-----------------------------------------------------------------------
-- FloatingPointPower, version 0.0
-----------------------------------------------------------------------

Library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity fpow_op is
Generic (
 INPUTS: integer := 2; 
 OUTPUTS: integer := 1; 
 DATA_SIZE_IN: integer := 32; --we default to single precision
 DATA_SIZE_OUT: integer := 32
);
port (
    -- inputs
    clk          : in std_logic;
    rst          : in std_logic;
     lhs          : in std_logic_vector(63 downto 0);
    lhs_valid    : in std_logic;
    rhs          : in std_logic_vector(63  downto 0);
    rhs_valid    : in std_logic;
    result_ready : in std_logic;
    -- outputs
     result       : out std_logic_vector(65  downto 0);
    result_valid : out std_logic;
    lhs_ready    : out std_logic;
    rhs_ready    : out std_logic
  );
end entity;

architecture arch of fpow_op is
    
    
    -- legacy comment : main_component went here in component based version

    signal join_valid : STD_LOGIC;

    signal buff_valid, oehb_valid, oehb_ready : STD_LOGIC;
    signal oehb_dataOut, oehb_datain : std_logic_vector(0 downto 0);

    --intermediate input signals for float conversion
    signal ip_lhs, ip_rhs : std_logic_vector(65 downto 0);

    --intermidiate output signal(s) for float conversion
    signal ip_result : std_logic_vector(65 downto 0);

    

    begin


          join_inputs : entity work.join(arch) generic map(2) 
    port map( 
      -- inputs 
      ins_valid(0) => lhs_valid,
      ins_valid(1) => rhs_valid,
      outs_ready   => oehb_ready,
      -- outputs 
      outs_valid   => join_valid, 
      ins_ready(0) => lhs_ready, 
      ins_ready(1) => rhs_ready
    );

        buff: entity work.delay_buffer(arch) generic map(526)
        port map(clk,
                rst,
                join_valid,
                oehb_ready,
                buff_valid);

        oehb: entity work.oehb_dataless(arch)
            port map(
            clk        => clk,
            rst        => rst,
            ins_valid  => buff_valid,
            outs_ready => result_ready,
            outs_valid => result_valid,
            ins_ready  => oehb_ready
            );

        ieee2nfloat_0: entity work.InputIEEE_64bit(arch)
                port map (
                    --input
                    X =>lhs,
                    --output
                    R => ip_lhs
                );

        ieee2nfloat_1: entity work.InputIEEE_64bit(arch)
                port map (
                    --input
                    X => rhs,
                    --output
                    R => ip_rhs
                );

        

        -- No output conversion: direct assignment
       result <= ip_result;

        operator : entity work.FloatingPointPower(arch)
        port map (
            clk   => clk,
            ce_1 => oehb_ready,
            ce_2 => oehb_ready,
            ce_3 => oehb_ready,
            ce_4 => oehb_ready,
            ce_5 => oehb_ready,
            ce_6 => oehb_ready,
            ce_7 => oehb_ready,
            ce_8 => oehb_ready,
            ce_9 => oehb_ready,
            ce_10 => oehb_ready,
            ce_11 => oehb_ready,
            ce_12 => oehb_ready,
            ce_13 => oehb_ready,
            ce_14 => oehb_ready,
            ce_15 => oehb_ready,
            ce_16 => oehb_ready,
            ce_17 => oehb_ready,
            ce_18 => oehb_ready,
            ce_19 => oehb_ready,
            ce_20 => oehb_ready,
            ce_21 => oehb_ready,
            ce_22 => oehb_ready,
            ce_23 => oehb_ready,
            ce_24 => oehb_ready,
            ce_25 => oehb_ready,
            ce_26 => oehb_ready,
            ce_27 => oehb_ready,
            ce_28 => oehb_ready,
            ce_29 => oehb_ready,
            ce_30 => oehb_ready,
            ce_31 => oehb_ready,
            ce_32 => oehb_ready,
            ce_33 => oehb_ready,
            ce_34 => oehb_ready,
            ce_35 => oehb_ready,
            ce_36 => oehb_ready,
            ce_37 => oehb_ready,
            ce_38 => oehb_ready,
            ce_39 => oehb_ready,
            ce_40 => oehb_ready,
            ce_41 => oehb_ready,
            ce_42 => oehb_ready,
            ce_43 => oehb_ready,
            ce_44 => oehb_ready,
            ce_45 => oehb_ready,
            ce_46 => oehb_ready,
            ce_47 => oehb_ready,
            ce_48 => oehb_ready,
            ce_49 => oehb_ready,
            ce_50 => oehb_ready,
            ce_51 => oehb_ready,
            ce_52 => oehb_ready,
            ce_53 => oehb_ready,
            ce_54 => oehb_ready,
            ce_55 => oehb_ready,
            ce_56 => oehb_ready,
            ce_57 => oehb_ready,
            ce_58 => oehb_ready,
            ce_59 => oehb_ready,
            ce_60 => oehb_ready,
            ce_61 => oehb_ready,
            ce_62 => oehb_ready,
            ce_63 => oehb_ready,
            ce_64 => oehb_ready,
            ce_65 => oehb_ready,
            ce_66 => oehb_ready,
            ce_67 => oehb_ready,
            ce_68 => oehb_ready,
            ce_69 => oehb_ready,
            ce_70 => oehb_ready,
            ce_71 => oehb_ready,
            ce_72 => oehb_ready,
            ce_73 => oehb_ready,
            ce_74 => oehb_ready,
            ce_75 => oehb_ready,
            ce_76 => oehb_ready,
            ce_77 => oehb_ready,
            ce_78 => oehb_ready,
            ce_79 => oehb_ready,
            ce_80 => oehb_ready,
            ce_81 => oehb_ready,
            ce_82 => oehb_ready,
            ce_83 => oehb_ready,
            ce_84 => oehb_ready,
            ce_85 => oehb_ready,
            ce_86 => oehb_ready,
            ce_87 => oehb_ready,
            ce_88 => oehb_ready,
            ce_89 => oehb_ready,
            ce_90 => oehb_ready,
            ce_91 => oehb_ready,
            ce_92 => oehb_ready,
            ce_93 => oehb_ready,
            ce_94 => oehb_ready,
            ce_95 => oehb_ready,
            ce_96 => oehb_ready,
            ce_97 => oehb_ready,
            ce_98 => oehb_ready,
            ce_99 => oehb_ready,
            ce_100 => oehb_ready,
            ce_101 => oehb_ready,
            ce_102 => oehb_ready,
            ce_103 => oehb_ready,
            ce_104 => oehb_ready,
            ce_105 => oehb_ready,
            ce_106 => oehb_ready,
            ce_107 => oehb_ready,
            ce_108 => oehb_ready,
            ce_109 => oehb_ready,
            ce_110 => oehb_ready,
            ce_111 => oehb_ready,
            ce_112 => oehb_ready,
            ce_113 => oehb_ready,
            ce_114 => oehb_ready,
            ce_115 => oehb_ready,
            ce_116 => oehb_ready,
            ce_117 => oehb_ready,
            ce_118 => oehb_ready,
            ce_119 => oehb_ready,
            ce_120 => oehb_ready,
            ce_121 => oehb_ready,
            ce_122 => oehb_ready,
            ce_123 => oehb_ready,
            ce_124 => oehb_ready,
            ce_125 => oehb_ready,
            ce_126 => oehb_ready,
            ce_127 => oehb_ready,
            ce_128 => oehb_ready,
            ce_129 => oehb_ready,
            ce_130 => oehb_ready,
            ce_131 => oehb_ready,
            ce_132 => oehb_ready,
            ce_133 => oehb_ready,
            ce_134 => oehb_ready,
            ce_135 => oehb_ready,
            ce_136 => oehb_ready,
            ce_137 => oehb_ready,
            ce_138 => oehb_ready,
            ce_139 => oehb_ready,
            ce_140 => oehb_ready,
            ce_141 => oehb_ready,
            ce_142 => oehb_ready,
            ce_143 => oehb_ready,
            ce_144 => oehb_ready,
            ce_145 => oehb_ready,
            ce_146 => oehb_ready,
            ce_147 => oehb_ready,
            ce_148 => oehb_ready,
            ce_149 => oehb_ready,
            ce_150 => oehb_ready,
            ce_151 => oehb_ready,
            ce_152 => oehb_ready,
            ce_153 => oehb_ready,
            ce_154 => oehb_ready,
            ce_155 => oehb_ready,
            ce_156 => oehb_ready,
            ce_157 => oehb_ready,
            ce_158 => oehb_ready,
            ce_159 => oehb_ready,
            ce_160 => oehb_ready,
            ce_161 => oehb_ready,
            ce_162 => oehb_ready,
            ce_163 => oehb_ready,
            ce_164 => oehb_ready,
            ce_165 => oehb_ready,
            ce_166 => oehb_ready,
            ce_167 => oehb_ready,
            ce_168 => oehb_ready,
            ce_169 => oehb_ready,
            ce_170 => oehb_ready,
            ce_171 => oehb_ready,
            ce_172 => oehb_ready,
            ce_173 => oehb_ready,
            ce_174 => oehb_ready,
            ce_175 => oehb_ready,
            ce_176 => oehb_ready,
            ce_177 => oehb_ready,
            ce_178 => oehb_ready,
            ce_179 => oehb_ready,
            ce_180 => oehb_ready,
            ce_181 => oehb_ready,
            ce_182 => oehb_ready,
            ce_183 => oehb_ready,
            ce_184 => oehb_ready,
            ce_185 => oehb_ready,
            ce_186 => oehb_ready,
            ce_187 => oehb_ready,
            ce_188 => oehb_ready,
            ce_189 => oehb_ready,
            ce_190 => oehb_ready,
            ce_191 => oehb_ready,
            ce_192 => oehb_ready,
            ce_193 => oehb_ready,
            ce_194 => oehb_ready,
            ce_195 => oehb_ready,
            ce_196 => oehb_ready,
            ce_197 => oehb_ready,
            ce_198 => oehb_ready,
            ce_199 => oehb_ready,
            ce_200 => oehb_ready,
            ce_201 => oehb_ready,
            ce_202 => oehb_ready,
            ce_203 => oehb_ready,
            ce_204 => oehb_ready,
            ce_205 => oehb_ready,
            ce_206 => oehb_ready,
            ce_207 => oehb_ready,
            ce_208 => oehb_ready,
            ce_209 => oehb_ready,
            ce_210 => oehb_ready,
            ce_211 => oehb_ready,
            ce_212 => oehb_ready,
            ce_213 => oehb_ready,
            ce_214 => oehb_ready,
            ce_215 => oehb_ready,
            ce_216 => oehb_ready,
            ce_217 => oehb_ready,
            ce_218 => oehb_ready,
            ce_219 => oehb_ready,
            ce_220 => oehb_ready,
            ce_221 => oehb_ready,
            ce_222 => oehb_ready,
            ce_223 => oehb_ready,
            ce_224 => oehb_ready,
            ce_225 => oehb_ready,
            ce_226 => oehb_ready,
            ce_227 => oehb_ready,
            ce_228 => oehb_ready,
            ce_229 => oehb_ready,
            ce_230 => oehb_ready,
            ce_231 => oehb_ready,
            ce_232 => oehb_ready,
            ce_233 => oehb_ready,
            ce_234 => oehb_ready,
            ce_235 => oehb_ready,
            ce_236 => oehb_ready,
            ce_237 => oehb_ready,
            ce_238 => oehb_ready,
            ce_239 => oehb_ready,
            ce_240 => oehb_ready,
            ce_241 => oehb_ready,
            ce_242 => oehb_ready,
            ce_243 => oehb_ready,
            ce_244 => oehb_ready,
            ce_245 => oehb_ready,
            ce_246 => oehb_ready,
            ce_247 => oehb_ready,
            ce_248 => oehb_ready,
            ce_249 => oehb_ready,
            ce_250 => oehb_ready,
            ce_251 => oehb_ready,
            ce_252 => oehb_ready,
            ce_253 => oehb_ready,
            ce_254 => oehb_ready,
            ce_255 => oehb_ready,
            ce_256 => oehb_ready,
            ce_257 => oehb_ready,
            ce_258 => oehb_ready,
            ce_259 => oehb_ready,
            ce_260 => oehb_ready,
            ce_261 => oehb_ready,
            ce_262 => oehb_ready,
            ce_263 => oehb_ready,
            ce_264 => oehb_ready,
            ce_265 => oehb_ready,
            ce_266 => oehb_ready,
            ce_267 => oehb_ready,
            ce_268 => oehb_ready,
            ce_269 => oehb_ready,
            ce_270 => oehb_ready,
            ce_271 => oehb_ready,
            ce_272 => oehb_ready,
            ce_273 => oehb_ready,
            ce_274 => oehb_ready,
            ce_275 => oehb_ready,
            ce_276 => oehb_ready,
            ce_277 => oehb_ready,
            ce_278 => oehb_ready,
            ce_279 => oehb_ready,
            ce_280 => oehb_ready,
            ce_281 => oehb_ready,
            ce_282 => oehb_ready,
            ce_283 => oehb_ready,
            ce_284 => oehb_ready,
            ce_285 => oehb_ready,
            ce_286 => oehb_ready,
            ce_287 => oehb_ready,
            ce_288 => oehb_ready,
            ce_289 => oehb_ready,
            ce_290 => oehb_ready,
            ce_291 => oehb_ready,
            ce_292 => oehb_ready,
            ce_293 => oehb_ready,
            ce_294 => oehb_ready,
            ce_295 => oehb_ready,
            ce_296 => oehb_ready,
            ce_297 => oehb_ready,
            ce_298 => oehb_ready,
            ce_299 => oehb_ready,
            ce_300 => oehb_ready,
            ce_301 => oehb_ready,
            ce_302 => oehb_ready,
            ce_303 => oehb_ready,
            ce_304 => oehb_ready,
            ce_305 => oehb_ready,
            ce_306 => oehb_ready,
            ce_307 => oehb_ready,
            ce_308 => oehb_ready,
            ce_309 => oehb_ready,
            ce_310 => oehb_ready,
            ce_311 => oehb_ready,
            ce_312 => oehb_ready,
            ce_313 => oehb_ready,
            ce_314 => oehb_ready,
            ce_315 => oehb_ready,
            ce_316 => oehb_ready,
            ce_317 => oehb_ready,
            ce_318 => oehb_ready,
            ce_319 => oehb_ready,
            ce_320 => oehb_ready,
            ce_321 => oehb_ready,
            ce_322 => oehb_ready,
            ce_323 => oehb_ready,
            ce_324 => oehb_ready,
            ce_325 => oehb_ready,
            ce_326 => oehb_ready,
            ce_327 => oehb_ready,
            ce_328 => oehb_ready,
            ce_329 => oehb_ready,
            ce_330 => oehb_ready,
            ce_331 => oehb_ready,
            ce_332 => oehb_ready,
            ce_333 => oehb_ready,
            ce_334 => oehb_ready,
            ce_335 => oehb_ready,
            ce_336 => oehb_ready,
            ce_337 => oehb_ready,
            ce_338 => oehb_ready,
            ce_339 => oehb_ready,
            ce_340 => oehb_ready,
            ce_341 => oehb_ready,
            ce_342 => oehb_ready,
            ce_343 => oehb_ready,
            ce_344 => oehb_ready,
            ce_345 => oehb_ready,
            ce_346 => oehb_ready,
            ce_347 => oehb_ready,
            ce_348 => oehb_ready,
            ce_349 => oehb_ready,
            ce_350 => oehb_ready,
            ce_351 => oehb_ready,
            ce_352 => oehb_ready,
            ce_353 => oehb_ready,
            ce_354 => oehb_ready,
            ce_355 => oehb_ready,
            ce_356 => oehb_ready,
            ce_357 => oehb_ready,
            ce_358 => oehb_ready,
            ce_359 => oehb_ready,
            ce_360 => oehb_ready,
            ce_361 => oehb_ready,
            ce_362 => oehb_ready,
            ce_363 => oehb_ready,
            ce_364 => oehb_ready,
            ce_365 => oehb_ready,
            ce_366 => oehb_ready,
            ce_367 => oehb_ready,
            ce_368 => oehb_ready,
            ce_369 => oehb_ready,
            ce_370 => oehb_ready,
            ce_371 => oehb_ready,
            ce_372 => oehb_ready,
            ce_373 => oehb_ready,
            ce_374 => oehb_ready,
            ce_375 => oehb_ready,
            ce_376 => oehb_ready,
            ce_377 => oehb_ready,
            ce_378 => oehb_ready,
            ce_379 => oehb_ready,
            ce_380 => oehb_ready,
            ce_381 => oehb_ready,
            ce_382 => oehb_ready,
            ce_383 => oehb_ready,
            ce_384 => oehb_ready,
            ce_385 => oehb_ready,
            ce_386 => oehb_ready,
            ce_387 => oehb_ready,
            ce_388 => oehb_ready,
            ce_389 => oehb_ready,
            ce_390 => oehb_ready,
            ce_391 => oehb_ready,
            ce_392 => oehb_ready,
            ce_393 => oehb_ready,
            ce_394 => oehb_ready,
            ce_395 => oehb_ready,
            ce_396 => oehb_ready,
            ce_397 => oehb_ready,
            ce_398 => oehb_ready,
            ce_399 => oehb_ready,
            ce_400 => oehb_ready,
            ce_401 => oehb_ready,
            ce_402 => oehb_ready,
            ce_403 => oehb_ready,
            ce_404 => oehb_ready,
            ce_405 => oehb_ready,
            ce_406 => oehb_ready,
            ce_407 => oehb_ready,
            ce_408 => oehb_ready,
            ce_409 => oehb_ready,
            ce_410 => oehb_ready,
            ce_411 => oehb_ready,
            ce_412 => oehb_ready,
            ce_413 => oehb_ready,
            ce_414 => oehb_ready,
            ce_415 => oehb_ready,
            ce_416 => oehb_ready,
            ce_417 => oehb_ready,
            ce_418 => oehb_ready,
            ce_419 => oehb_ready,
            ce_420 => oehb_ready,
            ce_421 => oehb_ready,
            ce_422 => oehb_ready,
            ce_423 => oehb_ready,
            ce_424 => oehb_ready,
            ce_425 => oehb_ready,
            ce_426 => oehb_ready,
            ce_427 => oehb_ready,
            ce_428 => oehb_ready,
            ce_429 => oehb_ready,
            ce_430 => oehb_ready,
            ce_431 => oehb_ready,
            ce_432 => oehb_ready,
            ce_433 => oehb_ready,
            ce_434 => oehb_ready,
            ce_435 => oehb_ready,
            ce_436 => oehb_ready,
            ce_437 => oehb_ready,
            ce_438 => oehb_ready,
            ce_439 => oehb_ready,
            ce_440 => oehb_ready,
            ce_441 => oehb_ready,
            ce_442 => oehb_ready,
            ce_443 => oehb_ready,
            ce_444 => oehb_ready,
            ce_445 => oehb_ready,
            ce_446 => oehb_ready,
            ce_447 => oehb_ready,
            ce_448 => oehb_ready,
            ce_449 => oehb_ready,
            ce_450 => oehb_ready,
            ce_451 => oehb_ready,
            ce_452 => oehb_ready,
            ce_453 => oehb_ready,
            ce_454 => oehb_ready,
            ce_455 => oehb_ready,
            ce_456 => oehb_ready,
            ce_457 => oehb_ready,
            ce_458 => oehb_ready,
            ce_459 => oehb_ready,
            ce_460 => oehb_ready,
            ce_461 => oehb_ready,
            ce_462 => oehb_ready,
            ce_463 => oehb_ready,
            ce_464 => oehb_ready,
            ce_465 => oehb_ready,
            ce_466 => oehb_ready,
            ce_467 => oehb_ready,
            ce_468 => oehb_ready,
            ce_469 => oehb_ready,
            ce_470 => oehb_ready,
            ce_471 => oehb_ready,
            ce_472 => oehb_ready,
            ce_473 => oehb_ready,
            ce_474 => oehb_ready,
            ce_475 => oehb_ready,
            ce_476 => oehb_ready,
            ce_477 => oehb_ready,
            ce_478 => oehb_ready,
            ce_479 => oehb_ready,
            ce_480 => oehb_ready,
            ce_481 => oehb_ready,
            ce_482 => oehb_ready,
            ce_483 => oehb_ready,
            ce_484 => oehb_ready,
            ce_485 => oehb_ready,
            ce_486 => oehb_ready,
            ce_487 => oehb_ready,
            ce_488 => oehb_ready,
            ce_489 => oehb_ready,
            ce_490 => oehb_ready,
            ce_491 => oehb_ready,
            ce_492 => oehb_ready,
            ce_493 => oehb_ready,
            ce_494 => oehb_ready,
            ce_495 => oehb_ready,
            ce_496 => oehb_ready,
            ce_497 => oehb_ready,
            ce_498 => oehb_ready,
            ce_499 => oehb_ready,
            ce_500 => oehb_ready,
            ce_501 => oehb_ready,
            ce_502 => oehb_ready,
            ce_503 => oehb_ready,
            ce_504 => oehb_ready,
            ce_505 => oehb_ready,
            ce_506 => oehb_ready,
            ce_507 => oehb_ready,
            ce_508 => oehb_ready,
            ce_509 => oehb_ready,
            ce_510 => oehb_ready,
            ce_511 => oehb_ready,
            ce_512 => oehb_ready,
            ce_513 => oehb_ready,
            ce_514 => oehb_ready,
            ce_515 => oehb_ready,
            ce_516 => oehb_ready,
            ce_517 => oehb_ready,
            ce_518 => oehb_ready,
            ce_519 => oehb_ready,
            ce_520 => oehb_ready,
            ce_521 => oehb_ready,
            ce_522 => oehb_ready,
            ce_523 => oehb_ready,
            ce_524 => oehb_ready,
            ce_525 => oehb_ready,
            ce_526 => oehb_ready,
            ce_527 => oehb_ready,
            X     => ip_lhs,
            Y     => ip_rhs,
            R     => ip_result
        );
end architecture;



