--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid17
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid17 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid17 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid22
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid22 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid22 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid27
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid27 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid27 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid32
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid32 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid32 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid37
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid37 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid37 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid42
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid42 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid42 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid47
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid47 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid47 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid52
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid52 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid52 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid63
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid63 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid63 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid68
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid68 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid68 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid73
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid73 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid73 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid78
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid78 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid78 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid83
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid83 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid83 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid88
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid88 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid88 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid93
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid93 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid93 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid98
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid98 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid98 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid113
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid113 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid113 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid118
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid118 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid118 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid123
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid128
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid128 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid128 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid133
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid133 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid133 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid138
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid138 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid138 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid143
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid143 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid143 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid148
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid148 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid148 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid153
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid153 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid153 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid158
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid158 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid158 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid163
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid163 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid163 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid168
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid168 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid168 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid183
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid183 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid183 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid188
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid188 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid188 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid193
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid193 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid193 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid198
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid198 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid198 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid203
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid203 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid203 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid208
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid208 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid208 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid213
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid213 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid213 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid218
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid218 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid218 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid223
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid223 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid223 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid228
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid228 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid228 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid233
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid233 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid233 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid238
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid238 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid238 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid253
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid253 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid253 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid258
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid258 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid258 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid263
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid263 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid263 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid268
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid268 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid268 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid273
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid273 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid273 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid278
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid278 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid278 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid283
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid283 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid283 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid288
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid288 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid288 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid293
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid293 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid293 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid298
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid298 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid298 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid303
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid303 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid303 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid308
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid308 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid308 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid313
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid313 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid313 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid318
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid318 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid318 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq300_uid322
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid322 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid322 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq300_uid326
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid326 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid326 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid334
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid334 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid334 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq300_uid400
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq300_uid400 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq300_uid400 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid432
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid432 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid432 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid9
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid9 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid9 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid11
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid11 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid11 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid13
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid13 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid13 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid15
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid15 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid15 is
   component MultTable_Freq300_uid17 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy18_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid17
      port map ( X => Xtable_c0,
                 Y => Y1_copy18_c0);
   Y1_c0 <= Y1_copy18_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid20
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid20 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid20 is
   component MultTable_Freq300_uid22 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy23_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid22
      port map ( X => Xtable_c0,
                 Y => Y1_copy23_c0);
   Y1_c0 <= Y1_copy23_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid25
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid25 is
   component MultTable_Freq300_uid27 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy28_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid27
      port map ( X => Xtable_c0,
                 Y => Y1_copy28_c0);
   Y1_c0 <= Y1_copy28_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid30
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid30 is
   component MultTable_Freq300_uid32 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy33_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid32
      port map ( X => Xtable_c0,
                 Y => Y1_copy33_c0);
   Y1_c0 <= Y1_copy33_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid35
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid35 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid35 is
   component MultTable_Freq300_uid37 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy38_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid37
      port map ( X => Xtable_c0,
                 Y => Y1_copy38_c0);
   Y1_c0 <= Y1_copy38_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid40
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid40 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid40 is
   component MultTable_Freq300_uid42 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy43_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid42
      port map ( X => Xtable_c0,
                 Y => Y1_copy43_c0);
   Y1_c0 <= Y1_copy43_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid45
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid45 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid45 is
   component MultTable_Freq300_uid47 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy48_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid47
      port map ( X => Xtable_c0,
                 Y => Y1_copy48_c0);
   Y1_c0 <= Y1_copy48_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid50
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid50 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid50 is
   component MultTable_Freq300_uid52 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy53_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid52
      port map ( X => Xtable_c0,
                 Y => Y1_copy53_c0);
   Y1_c0 <= Y1_copy53_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid55
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid55 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid55 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid57
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid57 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid57 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid59
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid59 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid59 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid61
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid61 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid61 is
   component MultTable_Freq300_uid63 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy64_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid63
      port map ( X => Xtable_c0,
                 Y => Y1_copy64_c0);
   Y1_c0 <= Y1_copy64_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid66
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid66 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid66 is
   component MultTable_Freq300_uid68 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy69_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid68
      port map ( X => Xtable_c0,
                 Y => Y1_copy69_c0);
   Y1_c0 <= Y1_copy69_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid71
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid71 is
   component MultTable_Freq300_uid73 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy74_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid73
      port map ( X => Xtable_c0,
                 Y => Y1_copy74_c0);
   Y1_c0 <= Y1_copy74_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid76
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid76 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid76 is
   component MultTable_Freq300_uid78 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy79_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid78
      port map ( X => Xtable_c0,
                 Y => Y1_copy79_c0);
   Y1_c0 <= Y1_copy79_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid81
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid81 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid81 is
   component MultTable_Freq300_uid83 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy84_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid83
      port map ( X => Xtable_c0,
                 Y => Y1_copy84_c0);
   Y1_c0 <= Y1_copy84_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid86
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid86 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid86 is
   component MultTable_Freq300_uid88 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy89_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid88
      port map ( X => Xtable_c0,
                 Y => Y1_copy89_c0);
   Y1_c0 <= Y1_copy89_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid91
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid91 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid91 is
   component MultTable_Freq300_uid93 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy94_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid93
      port map ( X => Xtable_c0,
                 Y => Y1_copy94_c0);
   Y1_c0 <= Y1_copy94_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid96
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid96 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid96 is
   component MultTable_Freq300_uid98 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy99_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid98
      port map ( X => Xtable_c0,
                 Y => Y1_copy99_c0);
   Y1_c0 <= Y1_copy99_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid101
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid101 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid101 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid103
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid103 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid103 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid105
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid105 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid105 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid107
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid107 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid107 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid109
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid109 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid109 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid111
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid111 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid111 is
   component MultTable_Freq300_uid113 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy114_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid113
      port map ( X => Xtable_c0,
                 Y => Y1_copy114_c0);
   Y1_c0 <= Y1_copy114_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid116
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid116 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid116 is
   component MultTable_Freq300_uid118 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy119_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid118
      port map ( X => Xtable_c0,
                 Y => Y1_copy119_c0);
   Y1_c0 <= Y1_copy119_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid121
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid121 is
   component MultTable_Freq300_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy124_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid123
      port map ( X => Xtable_c0,
                 Y => Y1_copy124_c0);
   Y1_c0 <= Y1_copy124_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid126
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid126 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid126 is
   component MultTable_Freq300_uid128 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy129_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid128
      port map ( X => Xtable_c0,
                 Y => Y1_copy129_c0);
   Y1_c0 <= Y1_copy129_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid131
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid131 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid131 is
   component MultTable_Freq300_uid133 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy134_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid133
      port map ( X => Xtable_c0,
                 Y => Y1_copy134_c0);
   Y1_c0 <= Y1_copy134_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid136
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid136 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid136 is
   component MultTable_Freq300_uid138 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy139_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid138
      port map ( X => Xtable_c0,
                 Y => Y1_copy139_c0);
   Y1_c0 <= Y1_copy139_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid141
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid141 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid141 is
   component MultTable_Freq300_uid143 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy144_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid143
      port map ( X => Xtable_c0,
                 Y => Y1_copy144_c0);
   Y1_c0 <= Y1_copy144_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid146
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid146 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid146 is
   component MultTable_Freq300_uid148 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy149_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid148
      port map ( X => Xtable_c0,
                 Y => Y1_copy149_c0);
   Y1_c0 <= Y1_copy149_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid151
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid151 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid151 is
   component MultTable_Freq300_uid153 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy154_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid153
      port map ( X => Xtable_c0,
                 Y => Y1_copy154_c0);
   Y1_c0 <= Y1_copy154_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid156
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid156 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid156 is
   component MultTable_Freq300_uid158 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy159_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid158
      port map ( X => Xtable_c0,
                 Y => Y1_copy159_c0);
   Y1_c0 <= Y1_copy159_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid161
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid161 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid161 is
   component MultTable_Freq300_uid163 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy164_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid163
      port map ( X => Xtable_c0,
                 Y => Y1_copy164_c0);
   Y1_c0 <= Y1_copy164_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid166
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid166 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid166 is
   component MultTable_Freq300_uid168 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy169_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid168
      port map ( X => Xtable_c0,
                 Y => Y1_copy169_c0);
   Y1_c0 <= Y1_copy169_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid171
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid171 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid171 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid173
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid173 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid173 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid175
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid175 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid175 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid177
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid177 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid177 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid179
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid179 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid179 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid181
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid181 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid181 is
   component MultTable_Freq300_uid183 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy184_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid183
      port map ( X => Xtable_c0,
                 Y => Y1_copy184_c0);
   Y1_c0 <= Y1_copy184_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid186
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid186 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid186 is
   component MultTable_Freq300_uid188 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy189_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid188
      port map ( X => Xtable_c0,
                 Y => Y1_copy189_c0);
   Y1_c0 <= Y1_copy189_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid191
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid191 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid191 is
   component MultTable_Freq300_uid193 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy194_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid193
      port map ( X => Xtable_c0,
                 Y => Y1_copy194_c0);
   Y1_c0 <= Y1_copy194_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid196
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid196 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid196 is
   component MultTable_Freq300_uid198 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy199_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid198
      port map ( X => Xtable_c0,
                 Y => Y1_copy199_c0);
   Y1_c0 <= Y1_copy199_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid201
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid201 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid201 is
   component MultTable_Freq300_uid203 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy204_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid203
      port map ( X => Xtable_c0,
                 Y => Y1_copy204_c0);
   Y1_c0 <= Y1_copy204_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid206
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid206 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid206 is
   component MultTable_Freq300_uid208 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy209_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid208
      port map ( X => Xtable_c0,
                 Y => Y1_copy209_c0);
   Y1_c0 <= Y1_copy209_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid211
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid211 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid211 is
   component MultTable_Freq300_uid213 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy214_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid213
      port map ( X => Xtable_c0,
                 Y => Y1_copy214_c0);
   Y1_c0 <= Y1_copy214_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid216
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid216 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid216 is
   component MultTable_Freq300_uid218 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy219_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid218
      port map ( X => Xtable_c0,
                 Y => Y1_copy219_c0);
   Y1_c0 <= Y1_copy219_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid221
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid221 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid221 is
   component MultTable_Freq300_uid223 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy224_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid223
      port map ( X => Xtable_c0,
                 Y => Y1_copy224_c0);
   Y1_c0 <= Y1_copy224_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid226
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid226 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid226 is
   component MultTable_Freq300_uid228 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy229_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid228
      port map ( X => Xtable_c0,
                 Y => Y1_copy229_c0);
   Y1_c0 <= Y1_copy229_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid231
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid231 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid231 is
   component MultTable_Freq300_uid233 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy234_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid233
      port map ( X => Xtable_c0,
                 Y => Y1_copy234_c0);
   Y1_c0 <= Y1_copy234_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid236
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid236 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid236 is
   component MultTable_Freq300_uid238 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy239_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid238
      port map ( X => Xtable_c0,
                 Y => Y1_copy239_c0);
   Y1_c0 <= Y1_copy239_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid241
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid241 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid241 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid243
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid243 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid243 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid245
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid245 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid245 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid247
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid247 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid247 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid249
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid249 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid249 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid251
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid251 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid251 is
   component MultTable_Freq300_uid253 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy254_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid253
      port map ( X => Xtable_c0,
                 Y => Y1_copy254_c0);
   Y1_c0 <= Y1_copy254_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid256
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid256 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid256 is
   component MultTable_Freq300_uid258 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy259_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid258
      port map ( X => Xtable_c0,
                 Y => Y1_copy259_c0);
   Y1_c0 <= Y1_copy259_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid261
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid261 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid261 is
   component MultTable_Freq300_uid263 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy264_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid263
      port map ( X => Xtable_c0,
                 Y => Y1_copy264_c0);
   Y1_c0 <= Y1_copy264_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid266
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid266 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid266 is
   component MultTable_Freq300_uid268 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy269_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid268
      port map ( X => Xtable_c0,
                 Y => Y1_copy269_c0);
   Y1_c0 <= Y1_copy269_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid271
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid271 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid271 is
   component MultTable_Freq300_uid273 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy274_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid273
      port map ( X => Xtable_c0,
                 Y => Y1_copy274_c0);
   Y1_c0 <= Y1_copy274_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid276
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid276 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid276 is
   component MultTable_Freq300_uid278 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy279_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid278
      port map ( X => Xtable_c0,
                 Y => Y1_copy279_c0);
   Y1_c0 <= Y1_copy279_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid281
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid281 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid281 is
   component MultTable_Freq300_uid283 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy284_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid283
      port map ( X => Xtable_c0,
                 Y => Y1_copy284_c0);
   Y1_c0 <= Y1_copy284_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid286
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid286 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid286 is
   component MultTable_Freq300_uid288 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy289_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid288
      port map ( X => Xtable_c0,
                 Y => Y1_copy289_c0);
   Y1_c0 <= Y1_copy289_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid291
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid291 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid291 is
   component MultTable_Freq300_uid293 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy294_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid293
      port map ( X => Xtable_c0,
                 Y => Y1_copy294_c0);
   Y1_c0 <= Y1_copy294_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid296
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid296 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid296 is
   component MultTable_Freq300_uid298 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy299_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid298
      port map ( X => Xtable_c0,
                 Y => Y1_copy299_c0);
   Y1_c0 <= Y1_copy299_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid301
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid301 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid301 is
   component MultTable_Freq300_uid303 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy304_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid303
      port map ( X => Xtable_c0,
                 Y => Y1_copy304_c0);
   Y1_c0 <= Y1_copy304_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid306
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid306 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid306 is
   component MultTable_Freq300_uid308 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy309_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid308
      port map ( X => Xtable_c0,
                 Y => Y1_copy309_c0);
   Y1_c0 <= Y1_copy309_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid311
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid311 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid311 is
   component MultTable_Freq300_uid313 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy314_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid313
      port map ( X => Xtable_c0,
                 Y => Y1_copy314_c0);
   Y1_c0 <= Y1_copy314_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x3_Freq300_uid316
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid316 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid316 is
   component MultTable_Freq300_uid318 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy319_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid318
      port map ( X => Xtable_c0,
                 Y => Y1_copy319_c0);
   Y1_c0 <= Y1_copy319_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_84_Freq300_uid972
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_84_Freq300_uid972 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(83 downto 0);
          Y : in  std_logic_vector(83 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(83 downto 0)   );
end entity;

architecture arch of IntAdder_84_Freq300_uid972 is
signal Rtmp_c2 :  std_logic_vector(83 downto 0);
signal X_c2 :  std_logic_vector(83 downto 0);
signal Y_c2 :  std_logic_vector(83 downto 0);
signal Cin_c1, Cin_c2 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               X_c2 <= X;
               Y_c2 <= Y;
               Cin_c2 <= Cin_c1;
            end if;
         end if;
      end process;
   Rtmp_c2 <= X_c2 + Y_c2 + Cin_c2;
   R <= Rtmp_c2;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_53x53_106_Freq300_uid5
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_53x53_106_Freq300_uid5 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          Y : in  std_logic_vector(52 downto 0);
          R : out  std_logic_vector(105 downto 0)   );
end entity;

architecture arch of IntMultiplier_53x53_106_Freq300_uid5 is
   component DSPBlock_17x24_Freq300_uid9 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid11 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid13 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid15 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid20 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid35 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid40 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid45 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid50 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid55 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid57 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid59 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid61 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid66 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid76 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid81 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid86 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid91 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid96 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid101 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid103 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid105 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid107 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid109 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid111 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid116 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid126 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid131 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid136 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid141 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid146 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid151 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid156 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid161 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid166 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid171 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid173 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid175 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid177 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid179 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid181 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid186 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid191 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid196 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid201 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid206 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid211 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid216 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid221 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid226 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid231 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid236 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid241 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid243 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid245 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid247 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid249 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid251 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid256 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid261 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid266 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid271 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid276 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid281 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid286 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid291 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid296 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid301 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid306 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid311 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid316 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid322 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid326 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid334 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq300_uid400 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid432 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntAdder_84_Freq300_uid972 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(83 downto 0);
             Y : in  std_logic_vector(83 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(83 downto 0)   );
   end component;

signal XX_m6_c0 :  std_logic_vector(52 downto 0);
signal YY_m6_c0 :  std_logic_vector(52 downto 0);
signal tile_0_X_c0 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_0_output_c0 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w0_0_c0, bh7_w0_0_c1 :  std_logic;
signal bh7_w1_0_c0, bh7_w1_0_c1 :  std_logic;
signal bh7_w2_0_c0, bh7_w2_0_c1 :  std_logic;
signal bh7_w3_0_c0, bh7_w3_0_c1 :  std_logic;
signal bh7_w4_0_c0, bh7_w4_0_c1 :  std_logic;
signal bh7_w5_0_c0, bh7_w5_0_c1 :  std_logic;
signal bh7_w6_0_c0, bh7_w6_0_c1 :  std_logic;
signal bh7_w7_0_c0, bh7_w7_0_c1 :  std_logic;
signal bh7_w8_0_c0, bh7_w8_0_c1 :  std_logic;
signal bh7_w9_0_c0, bh7_w9_0_c1 :  std_logic;
signal bh7_w10_0_c0, bh7_w10_0_c1 :  std_logic;
signal bh7_w11_0_c0, bh7_w11_0_c1 :  std_logic;
signal bh7_w12_0_c0, bh7_w12_0_c1 :  std_logic;
signal bh7_w13_0_c0, bh7_w13_0_c1 :  std_logic;
signal bh7_w14_0_c0, bh7_w14_0_c1 :  std_logic;
signal bh7_w15_0_c0, bh7_w15_0_c1 :  std_logic;
signal bh7_w16_0_c0, bh7_w16_0_c1 :  std_logic;
signal bh7_w17_0_c0 :  std_logic;
signal bh7_w18_0_c0 :  std_logic;
signal bh7_w19_0_c0 :  std_logic;
signal bh7_w20_0_c0 :  std_logic;
signal bh7_w21_0_c0 :  std_logic;
signal bh7_w22_0_c0 :  std_logic;
signal bh7_w23_0_c0 :  std_logic;
signal bh7_w24_0_c0 :  std_logic;
signal bh7_w25_0_c0 :  std_logic;
signal bh7_w26_0_c0 :  std_logic;
signal bh7_w27_0_c0 :  std_logic;
signal bh7_w28_0_c0 :  std_logic;
signal bh7_w29_0_c0 :  std_logic;
signal bh7_w30_0_c0 :  std_logic;
signal bh7_w31_0_c0 :  std_logic;
signal bh7_w32_0_c0 :  std_logic;
signal bh7_w33_0_c0 :  std_logic;
signal bh7_w34_0_c0 :  std_logic;
signal bh7_w35_0_c0 :  std_logic;
signal bh7_w36_0_c0 :  std_logic;
signal bh7_w37_0_c0 :  std_logic;
signal bh7_w38_0_c0 :  std_logic;
signal bh7_w39_0_c0 :  std_logic;
signal bh7_w40_0_c0 :  std_logic;
signal tile_1_X_c0 :  std_logic_vector(16 downto 0);
signal tile_1_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_1_output_c0 :  std_logic_vector(40 downto 0);
signal tile_1_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w17_1_c0 :  std_logic;
signal bh7_w18_1_c0 :  std_logic;
signal bh7_w19_1_c0 :  std_logic;
signal bh7_w20_1_c0 :  std_logic;
signal bh7_w21_1_c0 :  std_logic;
signal bh7_w22_1_c0 :  std_logic;
signal bh7_w23_1_c0 :  std_logic;
signal bh7_w24_1_c0 :  std_logic;
signal bh7_w25_1_c0 :  std_logic;
signal bh7_w26_1_c0 :  std_logic;
signal bh7_w27_1_c0 :  std_logic;
signal bh7_w28_1_c0 :  std_logic;
signal bh7_w29_1_c0 :  std_logic;
signal bh7_w30_1_c0 :  std_logic;
signal bh7_w31_1_c0 :  std_logic;
signal bh7_w32_1_c0 :  std_logic;
signal bh7_w33_1_c0 :  std_logic;
signal bh7_w34_1_c0 :  std_logic;
signal bh7_w35_1_c0 :  std_logic;
signal bh7_w36_1_c0 :  std_logic;
signal bh7_w37_1_c0 :  std_logic;
signal bh7_w38_1_c0 :  std_logic;
signal bh7_w39_1_c0 :  std_logic;
signal bh7_w40_1_c0 :  std_logic;
signal bh7_w41_0_c0 :  std_logic;
signal bh7_w42_0_c0 :  std_logic;
signal bh7_w43_0_c0 :  std_logic;
signal bh7_w44_0_c0 :  std_logic;
signal bh7_w45_0_c0 :  std_logic;
signal bh7_w46_0_c0 :  std_logic;
signal bh7_w47_0_c0 :  std_logic;
signal bh7_w48_0_c0 :  std_logic;
signal bh7_w49_0_c0 :  std_logic;
signal bh7_w50_0_c0 :  std_logic;
signal bh7_w51_0_c0 :  std_logic;
signal bh7_w52_0_c0 :  std_logic;
signal bh7_w53_0_c0 :  std_logic;
signal bh7_w54_0_c0 :  std_logic;
signal bh7_w55_0_c0 :  std_logic;
signal bh7_w56_0_c0 :  std_logic;
signal bh7_w57_0_c0 :  std_logic;
signal tile_2_X_c0 :  std_logic_vector(16 downto 0);
signal tile_2_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_2_output_c0 :  std_logic_vector(40 downto 0);
signal tile_2_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w34_2_c0 :  std_logic;
signal bh7_w35_2_c0 :  std_logic;
signal bh7_w36_2_c0 :  std_logic;
signal bh7_w37_2_c0 :  std_logic;
signal bh7_w38_2_c0 :  std_logic;
signal bh7_w39_2_c0 :  std_logic;
signal bh7_w40_2_c0 :  std_logic;
signal bh7_w41_1_c0 :  std_logic;
signal bh7_w42_1_c0 :  std_logic;
signal bh7_w43_1_c0 :  std_logic;
signal bh7_w44_1_c0 :  std_logic;
signal bh7_w45_1_c0 :  std_logic;
signal bh7_w46_1_c0 :  std_logic;
signal bh7_w47_1_c0 :  std_logic;
signal bh7_w48_1_c0 :  std_logic;
signal bh7_w49_1_c0 :  std_logic;
signal bh7_w50_1_c0 :  std_logic;
signal bh7_w51_1_c0 :  std_logic;
signal bh7_w52_1_c0 :  std_logic;
signal bh7_w53_1_c0 :  std_logic;
signal bh7_w54_1_c0 :  std_logic;
signal bh7_w55_1_c0 :  std_logic;
signal bh7_w56_1_c0 :  std_logic;
signal bh7_w57_1_c0 :  std_logic;
signal bh7_w58_0_c0 :  std_logic;
signal bh7_w59_0_c0, bh7_w59_0_c1 :  std_logic;
signal bh7_w60_0_c0, bh7_w60_0_c1 :  std_logic;
signal bh7_w61_0_c0, bh7_w61_0_c1 :  std_logic;
signal bh7_w62_0_c0, bh7_w62_0_c1 :  std_logic;
signal bh7_w63_0_c0 :  std_logic;
signal bh7_w64_0_c0, bh7_w64_0_c1 :  std_logic;
signal bh7_w65_0_c0, bh7_w65_0_c1 :  std_logic;
signal bh7_w66_0_c0 :  std_logic;
signal bh7_w67_0_c0, bh7_w67_0_c1 :  std_logic;
signal bh7_w68_0_c0 :  std_logic;
signal bh7_w69_0_c0, bh7_w69_0_c1 :  std_logic;
signal bh7_w70_0_c0, bh7_w70_0_c1 :  std_logic;
signal bh7_w71_0_c0 :  std_logic;
signal bh7_w72_0_c0, bh7_w72_0_c1 :  std_logic;
signal bh7_w73_0_c0 :  std_logic;
signal bh7_w74_0_c0, bh7_w74_0_c1 :  std_logic;
signal tile_3_X_c0 :  std_logic_vector(1 downto 0);
signal tile_3_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_3_output_c0 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w72_1_c0 :  std_logic;
signal bh7_w73_1_c0 :  std_logic;
signal bh7_w74_1_c0 :  std_logic;
signal bh7_w75_0_c0 :  std_logic;
signal bh7_w76_0_c0 :  std_logic;
signal tile_4_X_c0 :  std_logic_vector(1 downto 0);
signal tile_4_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_4_output_c0 :  std_logic_vector(4 downto 0);
signal tile_4_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w69_1_c0 :  std_logic;
signal bh7_w70_1_c0 :  std_logic;
signal bh7_w71_1_c0 :  std_logic;
signal bh7_w72_2_c0 :  std_logic;
signal bh7_w73_2_c0 :  std_logic;
signal tile_5_X_c0 :  std_logic_vector(1 downto 0);
signal tile_5_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_5_output_c0 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w66_1_c0 :  std_logic;
signal bh7_w67_1_c0 :  std_logic;
signal bh7_w68_1_c0 :  std_logic;
signal bh7_w69_2_c0 :  std_logic;
signal bh7_w70_2_c0 :  std_logic;
signal tile_6_X_c0 :  std_logic_vector(1 downto 0);
signal tile_6_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_6_output_c0 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w63_1_c0 :  std_logic;
signal bh7_w64_1_c0 :  std_logic;
signal bh7_w65_1_c0 :  std_logic;
signal bh7_w66_2_c0 :  std_logic;
signal bh7_w67_2_c0 :  std_logic;
signal tile_7_X_c0 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_7_output_c0 :  std_logic_vector(4 downto 0);
signal tile_7_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_1_c0 :  std_logic;
signal bh7_w61_1_c0 :  std_logic;
signal bh7_w62_1_c0 :  std_logic;
signal bh7_w63_2_c0 :  std_logic;
signal bh7_w64_2_c0 :  std_logic;
signal tile_8_X_c0 :  std_logic_vector(1 downto 0);
signal tile_8_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_8_output_c0 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_2_c0 :  std_logic;
signal bh7_w58_1_c0 :  std_logic;
signal bh7_w59_1_c0 :  std_logic;
signal bh7_w60_2_c0 :  std_logic;
signal bh7_w61_2_c0 :  std_logic;
signal tile_9_X_c0 :  std_logic_vector(1 downto 0);
signal tile_9_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_9_output_c0 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_2_c0 :  std_logic;
signal bh7_w55_2_c0 :  std_logic;
signal bh7_w56_2_c0 :  std_logic;
signal bh7_w57_3_c0 :  std_logic;
signal bh7_w58_2_c0 :  std_logic;
signal tile_10_X_c0 :  std_logic_vector(1 downto 0);
signal tile_10_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_10_output_c0 :  std_logic_vector(4 downto 0);
signal tile_10_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_2_c0 :  std_logic;
signal bh7_w52_2_c0 :  std_logic;
signal bh7_w53_2_c0 :  std_logic;
signal bh7_w54_3_c0 :  std_logic;
signal bh7_w55_3_c0 :  std_logic;
signal tile_11_X_c0 :  std_logic_vector(16 downto 0);
signal tile_11_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_11_output_c0 :  std_logic_vector(40 downto 0);
signal tile_11_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w24_2_c0 :  std_logic;
signal bh7_w25_2_c0, bh7_w25_2_c1 :  std_logic;
signal bh7_w26_2_c0 :  std_logic;
signal bh7_w27_2_c0, bh7_w27_2_c1 :  std_logic;
signal bh7_w28_2_c0 :  std_logic;
signal bh7_w29_2_c0, bh7_w29_2_c1 :  std_logic;
signal bh7_w30_2_c0 :  std_logic;
signal bh7_w31_2_c0, bh7_w31_2_c1 :  std_logic;
signal bh7_w32_2_c0 :  std_logic;
signal bh7_w33_2_c0, bh7_w33_2_c1 :  std_logic;
signal bh7_w34_3_c0 :  std_logic;
signal bh7_w35_3_c0 :  std_logic;
signal bh7_w36_3_c0 :  std_logic;
signal bh7_w37_3_c0 :  std_logic;
signal bh7_w38_3_c0 :  std_logic;
signal bh7_w39_3_c0 :  std_logic;
signal bh7_w40_3_c0 :  std_logic;
signal bh7_w41_2_c0 :  std_logic;
signal bh7_w42_2_c0 :  std_logic;
signal bh7_w43_2_c0 :  std_logic;
signal bh7_w44_2_c0 :  std_logic;
signal bh7_w45_2_c0 :  std_logic;
signal bh7_w46_2_c0 :  std_logic;
signal bh7_w47_2_c0 :  std_logic;
signal bh7_w48_2_c0 :  std_logic;
signal bh7_w49_2_c0 :  std_logic;
signal bh7_w50_2_c0 :  std_logic;
signal bh7_w51_3_c0 :  std_logic;
signal bh7_w52_3_c0 :  std_logic;
signal bh7_w53_3_c0 :  std_logic;
signal bh7_w54_4_c0 :  std_logic;
signal bh7_w55_4_c0 :  std_logic;
signal bh7_w56_3_c0 :  std_logic;
signal bh7_w57_4_c0 :  std_logic;
signal bh7_w58_3_c0 :  std_logic;
signal bh7_w59_2_c0, bh7_w59_2_c1 :  std_logic;
signal bh7_w60_3_c0, bh7_w60_3_c1 :  std_logic;
signal bh7_w61_3_c0, bh7_w61_3_c1 :  std_logic;
signal bh7_w62_2_c0, bh7_w62_2_c1 :  std_logic;
signal bh7_w63_3_c0 :  std_logic;
signal bh7_w64_3_c0, bh7_w64_3_c1 :  std_logic;
signal tile_12_X_c0 :  std_logic_vector(16 downto 0);
signal tile_12_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_12_output_c0 :  std_logic_vector(40 downto 0);
signal tile_12_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w41_3_c0 :  std_logic;
signal bh7_w42_3_c0 :  std_logic;
signal bh7_w43_3_c0 :  std_logic;
signal bh7_w44_3_c0 :  std_logic;
signal bh7_w45_3_c0 :  std_logic;
signal bh7_w46_3_c0 :  std_logic;
signal bh7_w47_3_c0 :  std_logic;
signal bh7_w48_3_c0, bh7_w48_3_c1 :  std_logic;
signal bh7_w49_3_c0 :  std_logic;
signal bh7_w50_3_c0 :  std_logic;
signal bh7_w51_4_c0 :  std_logic;
signal bh7_w52_4_c0 :  std_logic;
signal bh7_w53_4_c0 :  std_logic;
signal bh7_w54_5_c0 :  std_logic;
signal bh7_w55_5_c0 :  std_logic;
signal bh7_w56_4_c0 :  std_logic;
signal bh7_w57_5_c0 :  std_logic;
signal bh7_w58_4_c0 :  std_logic;
signal bh7_w59_3_c0, bh7_w59_3_c1 :  std_logic;
signal bh7_w60_4_c0, bh7_w60_4_c1 :  std_logic;
signal bh7_w61_4_c0, bh7_w61_4_c1 :  std_logic;
signal bh7_w62_3_c0, bh7_w62_3_c1 :  std_logic;
signal bh7_w63_4_c0 :  std_logic;
signal bh7_w64_4_c0, bh7_w64_4_c1 :  std_logic;
signal bh7_w65_2_c0, bh7_w65_2_c1 :  std_logic;
signal bh7_w66_3_c0 :  std_logic;
signal bh7_w67_3_c0, bh7_w67_3_c1 :  std_logic;
signal bh7_w68_2_c0 :  std_logic;
signal bh7_w69_3_c0, bh7_w69_3_c1 :  std_logic;
signal bh7_w70_3_c0, bh7_w70_3_c1 :  std_logic;
signal bh7_w71_2_c0 :  std_logic;
signal bh7_w72_3_c0, bh7_w72_3_c1 :  std_logic;
signal bh7_w73_3_c0 :  std_logic;
signal bh7_w74_2_c0, bh7_w74_2_c1 :  std_logic;
signal bh7_w75_1_c0 :  std_logic;
signal bh7_w76_1_c0, bh7_w76_1_c1 :  std_logic;
signal bh7_w77_0_c0, bh7_w77_0_c1 :  std_logic;
signal bh7_w78_0_c0, bh7_w78_0_c1 :  std_logic;
signal bh7_w79_0_c0, bh7_w79_0_c1 :  std_logic;
signal bh7_w80_0_c0, bh7_w80_0_c1 :  std_logic;
signal bh7_w81_0_c0, bh7_w81_0_c1 :  std_logic;
signal tile_13_X_c0 :  std_logic_vector(16 downto 0);
signal tile_13_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_13_output_c0 :  std_logic_vector(40 downto 0);
signal tile_13_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w58_5_c0, bh7_w58_5_c1 :  std_logic;
signal bh7_w59_4_c0, bh7_w59_4_c1 :  std_logic;
signal bh7_w60_5_c0, bh7_w60_5_c1 :  std_logic;
signal bh7_w61_5_c0, bh7_w61_5_c1 :  std_logic;
signal bh7_w62_4_c0, bh7_w62_4_c1 :  std_logic;
signal bh7_w63_5_c0, bh7_w63_5_c1 :  std_logic;
signal bh7_w64_5_c0, bh7_w64_5_c1 :  std_logic;
signal bh7_w65_3_c0, bh7_w65_3_c1 :  std_logic;
signal bh7_w66_4_c0 :  std_logic;
signal bh7_w67_4_c0, bh7_w67_4_c1 :  std_logic;
signal bh7_w68_3_c0 :  std_logic;
signal bh7_w69_4_c0, bh7_w69_4_c1 :  std_logic;
signal bh7_w70_4_c0, bh7_w70_4_c1 :  std_logic;
signal bh7_w71_3_c0 :  std_logic;
signal bh7_w72_4_c0, bh7_w72_4_c1 :  std_logic;
signal bh7_w73_4_c0 :  std_logic;
signal bh7_w74_3_c0, bh7_w74_3_c1 :  std_logic;
signal bh7_w75_2_c0, bh7_w75_2_c1 :  std_logic;
signal bh7_w76_2_c0, bh7_w76_2_c1 :  std_logic;
signal bh7_w77_1_c0, bh7_w77_1_c1 :  std_logic;
signal bh7_w78_1_c0, bh7_w78_1_c1 :  std_logic;
signal bh7_w79_1_c0, bh7_w79_1_c1 :  std_logic;
signal bh7_w80_1_c0, bh7_w80_1_c1 :  std_logic;
signal bh7_w81_1_c0, bh7_w81_1_c1 :  std_logic;
signal bh7_w82_0_c0, bh7_w82_0_c1 :  std_logic;
signal bh7_w83_0_c0, bh7_w83_0_c1 :  std_logic;
signal bh7_w84_0_c0, bh7_w84_0_c1 :  std_logic;
signal bh7_w85_0_c0, bh7_w85_0_c1 :  std_logic;
signal bh7_w86_0_c0, bh7_w86_0_c1 :  std_logic;
signal bh7_w87_0_c0, bh7_w87_0_c1 :  std_logic;
signal bh7_w88_0_c0, bh7_w88_0_c1 :  std_logic;
signal bh7_w89_0_c0, bh7_w89_0_c1 :  std_logic;
signal bh7_w90_0_c0, bh7_w90_0_c1 :  std_logic;
signal bh7_w91_0_c0, bh7_w91_0_c1 :  std_logic;
signal bh7_w92_0_c0, bh7_w92_0_c1 :  std_logic;
signal bh7_w93_0_c0, bh7_w93_0_c1 :  std_logic;
signal bh7_w94_0_c0, bh7_w94_0_c1 :  std_logic;
signal bh7_w95_0_c0, bh7_w95_0_c1 :  std_logic;
signal bh7_w96_0_c0, bh7_w96_0_c1 :  std_logic;
signal bh7_w97_0_c0, bh7_w97_0_c1 :  std_logic;
signal bh7_w98_0_c0, bh7_w98_0_c1 :  std_logic;
signal tile_14_X_c0 :  std_logic_vector(1 downto 0);
signal tile_14_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_14_output_c0 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_1_c0 :  std_logic;
signal bh7_w97_1_c0 :  std_logic;
signal bh7_w98_1_c0 :  std_logic;
signal bh7_w99_0_c0 :  std_logic;
signal bh7_w100_0_c0 :  std_logic;
signal tile_15_X_c0 :  std_logic_vector(1 downto 0);
signal tile_15_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_15_output_c0 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_1_c0 :  std_logic;
signal bh7_w94_1_c0 :  std_logic;
signal bh7_w95_1_c0 :  std_logic;
signal bh7_w96_2_c0 :  std_logic;
signal bh7_w97_2_c0 :  std_logic;
signal tile_16_X_c0 :  std_logic_vector(1 downto 0);
signal tile_16_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_16_output_c0 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_1_c0 :  std_logic;
signal bh7_w91_1_c0 :  std_logic;
signal bh7_w92_1_c0 :  std_logic;
signal bh7_w93_2_c0 :  std_logic;
signal bh7_w94_2_c0 :  std_logic;
signal tile_17_X_c0 :  std_logic_vector(1 downto 0);
signal tile_17_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_17_output_c0 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_1_c0 :  std_logic;
signal bh7_w88_1_c0 :  std_logic;
signal bh7_w89_1_c0 :  std_logic;
signal bh7_w90_2_c0 :  std_logic;
signal bh7_w91_2_c0 :  std_logic;
signal tile_18_X_c0 :  std_logic_vector(1 downto 0);
signal tile_18_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_18_output_c0 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_1_c0 :  std_logic;
signal bh7_w85_1_c0 :  std_logic;
signal bh7_w86_1_c0 :  std_logic;
signal bh7_w87_2_c0 :  std_logic;
signal bh7_w88_2_c0 :  std_logic;
signal tile_19_X_c0 :  std_logic_vector(1 downto 0);
signal tile_19_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_19_output_c0 :  std_logic_vector(4 downto 0);
signal tile_19_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w81_2_c0 :  std_logic;
signal bh7_w82_1_c0 :  std_logic;
signal bh7_w83_1_c0 :  std_logic;
signal bh7_w84_2_c0 :  std_logic;
signal bh7_w85_2_c0 :  std_logic;
signal tile_20_X_c0 :  std_logic_vector(1 downto 0);
signal tile_20_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_20_output_c0 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w78_2_c0 :  std_logic;
signal bh7_w79_2_c0 :  std_logic;
signal bh7_w80_2_c0 :  std_logic;
signal bh7_w81_3_c0 :  std_logic;
signal bh7_w82_2_c0 :  std_logic;
signal tile_21_X_c0 :  std_logic_vector(1 downto 0);
signal tile_21_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_21_output_c0 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w75_3_c0 :  std_logic;
signal bh7_w76_3_c0 :  std_logic;
signal bh7_w77_2_c0 :  std_logic;
signal bh7_w78_3_c0 :  std_logic;
signal bh7_w79_3_c0 :  std_logic;
signal tile_22_X_c0 :  std_logic_vector(0 downto 0);
signal tile_22_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_22_output_c0 :  std_logic_vector(0 downto 0);
signal tile_22_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w68_4_c0 :  std_logic;
signal tile_23_X_c0 :  std_logic_vector(3 downto 0);
signal tile_23_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_23_output_c0 :  std_logic_vector(3 downto 0);
signal tile_23_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w64_6_c0 :  std_logic;
signal bh7_w65_4_c0 :  std_logic;
signal bh7_w66_5_c0 :  std_logic;
signal bh7_w67_5_c0 :  std_logic;
signal tile_24_X_c0 :  std_logic_vector(3 downto 0);
signal tile_24_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_24_output_c0 :  std_logic_vector(3 downto 0);
signal tile_24_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w60_6_c0 :  std_logic;
signal bh7_w61_6_c0 :  std_logic;
signal bh7_w62_5_c0 :  std_logic;
signal bh7_w63_6_c0 :  std_logic;
signal tile_25_X_c0 :  std_logic_vector(3 downto 0);
signal tile_25_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_25_output_c0 :  std_logic_vector(3 downto 0);
signal tile_25_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w56_5_c0 :  std_logic;
signal bh7_w57_6_c0 :  std_logic;
signal bh7_w58_6_c0 :  std_logic;
signal bh7_w59_5_c0 :  std_logic;
signal tile_26_X_c0 :  std_logic_vector(3 downto 0);
signal tile_26_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_26_output_c0 :  std_logic_vector(3 downto 0);
signal tile_26_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w52_5_c0 :  std_logic;
signal bh7_w53_5_c0 :  std_logic;
signal bh7_w54_6_c0 :  std_logic;
signal bh7_w55_6_c0 :  std_logic;
signal tile_27_X_c0 :  std_logic_vector(1 downto 0);
signal tile_27_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_27_output_c0 :  std_logic_vector(3 downto 0);
signal tile_27_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w65_5_c0 :  std_logic;
signal bh7_w66_6_c0 :  std_logic;
signal bh7_w67_6_c0 :  std_logic;
signal bh7_w68_5_c0 :  std_logic;
signal tile_28_X_c0 :  std_logic_vector(2 downto 0);
signal tile_28_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_28_output_c0 :  std_logic_vector(4 downto 0);
signal tile_28_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w62_6_c0 :  std_logic;
signal bh7_w63_7_c0 :  std_logic;
signal bh7_w64_7_c0 :  std_logic;
signal bh7_w65_6_c0 :  std_logic;
signal bh7_w66_7_c0 :  std_logic;
signal tile_29_X_c0 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_29_output_c0 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w59_6_c0 :  std_logic;
signal bh7_w60_7_c0 :  std_logic;
signal bh7_w61_7_c0 :  std_logic;
signal bh7_w62_7_c0 :  std_logic;
signal bh7_w63_8_c0 :  std_logic;
signal tile_30_X_c0 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_30_output_c0 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w56_6_c0 :  std_logic;
signal bh7_w57_7_c0 :  std_logic;
signal bh7_w58_7_c0 :  std_logic;
signal bh7_w59_7_c0 :  std_logic;
signal bh7_w60_8_c0 :  std_logic;
signal tile_31_X_c0 :  std_logic_vector(2 downto 0);
signal tile_31_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_31_output_c0 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w53_6_c0 :  std_logic;
signal bh7_w54_7_c0 :  std_logic;
signal bh7_w55_7_c0 :  std_logic;
signal bh7_w56_7_c0 :  std_logic;
signal bh7_w57_8_c0 :  std_logic;
signal tile_32_X_c0 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_32_output_c0 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w50_4_c0 :  std_logic;
signal bh7_w51_5_c0 :  std_logic;
signal bh7_w52_6_c0 :  std_logic;
signal bh7_w53_7_c0 :  std_logic;
signal bh7_w54_8_c0 :  std_logic;
signal tile_33_X_c0 :  std_logic_vector(1 downto 0);
signal tile_33_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_33_output_c0 :  std_logic_vector(3 downto 0);
signal tile_33_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w63_9_c0 :  std_logic;
signal bh7_w64_8_c0 :  std_logic;
signal bh7_w65_7_c0 :  std_logic;
signal bh7_w66_8_c0 :  std_logic;
signal tile_34_X_c0 :  std_logic_vector(2 downto 0);
signal tile_34_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_34_output_c0 :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_9_c0 :  std_logic;
signal bh7_w61_8_c0 :  std_logic;
signal bh7_w62_8_c0 :  std_logic;
signal bh7_w63_10_c0 :  std_logic;
signal bh7_w64_9_c0 :  std_logic;
signal tile_35_X_c0 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_35_output_c0 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_9_c0 :  std_logic;
signal bh7_w58_8_c0 :  std_logic;
signal bh7_w59_8_c0 :  std_logic;
signal bh7_w60_10_c0 :  std_logic;
signal bh7_w61_9_c0 :  std_logic;
signal tile_36_X_c0 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_36_output_c0 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_9_c0 :  std_logic;
signal bh7_w55_8_c0 :  std_logic;
signal bh7_w56_8_c0 :  std_logic;
signal bh7_w57_10_c0 :  std_logic;
signal bh7_w58_9_c0 :  std_logic;
signal tile_37_X_c0 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_37_output_c0 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_6_c0 :  std_logic;
signal bh7_w52_7_c0 :  std_logic;
signal bh7_w53_8_c0 :  std_logic;
signal bh7_w54_10_c0 :  std_logic;
signal bh7_w55_9_c0 :  std_logic;
signal tile_38_X_c0 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_38_output_c0 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w48_4_c0 :  std_logic;
signal bh7_w49_4_c0 :  std_logic;
signal bh7_w50_5_c0 :  std_logic;
signal bh7_w51_7_c0 :  std_logic;
signal bh7_w52_8_c0 :  std_logic;
signal tile_39_X_c0 :  std_logic_vector(0 downto 0);
signal tile_39_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_39_output_c0 :  std_logic_vector(0 downto 0);
signal tile_39_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w85_3_c0 :  std_logic;
signal tile_40_X_c0 :  std_logic_vector(3 downto 0);
signal tile_40_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_40_output_c0 :  std_logic_vector(3 downto 0);
signal tile_40_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w81_4_c0 :  std_logic;
signal bh7_w82_3_c0 :  std_logic;
signal bh7_w83_2_c0 :  std_logic;
signal bh7_w84_3_c0 :  std_logic;
signal tile_41_X_c0 :  std_logic_vector(3 downto 0);
signal tile_41_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_41_output_c0 :  std_logic_vector(3 downto 0);
signal tile_41_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w77_3_c0 :  std_logic;
signal bh7_w78_4_c0 :  std_logic;
signal bh7_w79_4_c0 :  std_logic;
signal bh7_w80_3_c0 :  std_logic;
signal tile_42_X_c0 :  std_logic_vector(3 downto 0);
signal tile_42_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_42_output_c0 :  std_logic_vector(3 downto 0);
signal tile_42_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w73_5_c0 :  std_logic;
signal bh7_w74_4_c0 :  std_logic;
signal bh7_w75_4_c0 :  std_logic;
signal bh7_w76_4_c0 :  std_logic;
signal tile_43_X_c0 :  std_logic_vector(3 downto 0);
signal tile_43_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_43_output_c0 :  std_logic_vector(3 downto 0);
signal tile_43_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w69_5_c0 :  std_logic;
signal bh7_w70_5_c0 :  std_logic;
signal bh7_w71_4_c0 :  std_logic;
signal bh7_w72_5_c0 :  std_logic;
signal tile_44_X_c0 :  std_logic_vector(1 downto 0);
signal tile_44_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_44_output_c0 :  std_logic_vector(3 downto 0);
signal tile_44_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w82_4_c0 :  std_logic;
signal bh7_w83_3_c0 :  std_logic;
signal bh7_w84_4_c0 :  std_logic;
signal bh7_w85_4_c0 :  std_logic;
signal tile_45_X_c0 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_45_output_c0 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w79_5_c0 :  std_logic;
signal bh7_w80_4_c0 :  std_logic;
signal bh7_w81_5_c0 :  std_logic;
signal bh7_w82_5_c0 :  std_logic;
signal bh7_w83_4_c0 :  std_logic;
signal tile_46_X_c0 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_46_output_c0 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w76_5_c0 :  std_logic;
signal bh7_w77_4_c0 :  std_logic;
signal bh7_w78_5_c0 :  std_logic;
signal bh7_w79_6_c0 :  std_logic;
signal bh7_w80_5_c0 :  std_logic;
signal tile_47_X_c0 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_47_output_c0 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w73_6_c0 :  std_logic;
signal bh7_w74_5_c0 :  std_logic;
signal bh7_w75_5_c0 :  std_logic;
signal bh7_w76_6_c0 :  std_logic;
signal bh7_w77_5_c0 :  std_logic;
signal tile_48_X_c0 :  std_logic_vector(2 downto 0);
signal tile_48_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_48_output_c0 :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w70_6_c0 :  std_logic;
signal bh7_w71_5_c0 :  std_logic;
signal bh7_w72_6_c0 :  std_logic;
signal bh7_w73_7_c0 :  std_logic;
signal bh7_w74_6_c0 :  std_logic;
signal tile_49_X_c0 :  std_logic_vector(2 downto 0);
signal tile_49_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_49_output_c0 :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w67_7_c0 :  std_logic;
signal bh7_w68_6_c0 :  std_logic;
signal bh7_w69_6_c0 :  std_logic;
signal bh7_w70_7_c0 :  std_logic;
signal bh7_w71_6_c0 :  std_logic;
signal tile_50_X_c0 :  std_logic_vector(1 downto 0);
signal tile_50_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_50_output_c0 :  std_logic_vector(3 downto 0);
signal tile_50_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w80_6_c0 :  std_logic;
signal bh7_w81_6_c0 :  std_logic;
signal bh7_w82_6_c0 :  std_logic;
signal bh7_w83_5_c0 :  std_logic;
signal tile_51_X_c0 :  std_logic_vector(2 downto 0);
signal tile_51_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_51_output_c0 :  std_logic_vector(4 downto 0);
signal tile_51_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w77_6_c0 :  std_logic;
signal bh7_w78_6_c0 :  std_logic;
signal bh7_w79_7_c0 :  std_logic;
signal bh7_w80_7_c0 :  std_logic;
signal bh7_w81_7_c0 :  std_logic;
signal tile_52_X_c0 :  std_logic_vector(2 downto 0);
signal tile_52_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_52_output_c0 :  std_logic_vector(4 downto 0);
signal tile_52_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w74_7_c0 :  std_logic;
signal bh7_w75_6_c0 :  std_logic;
signal bh7_w76_7_c0 :  std_logic;
signal bh7_w77_7_c0 :  std_logic;
signal bh7_w78_7_c0 :  std_logic;
signal tile_53_X_c0 :  std_logic_vector(2 downto 0);
signal tile_53_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_53_output_c0 :  std_logic_vector(4 downto 0);
signal tile_53_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w71_7_c0 :  std_logic;
signal bh7_w72_7_c0 :  std_logic;
signal bh7_w73_8_c0 :  std_logic;
signal bh7_w74_8_c0 :  std_logic;
signal bh7_w75_7_c0 :  std_logic;
signal tile_54_X_c0 :  std_logic_vector(2 downto 0);
signal tile_54_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_54_output_c0 :  std_logic_vector(4 downto 0);
signal tile_54_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w68_7_c0 :  std_logic;
signal bh7_w69_7_c0 :  std_logic;
signal bh7_w70_8_c0 :  std_logic;
signal bh7_w71_8_c0 :  std_logic;
signal bh7_w72_8_c0 :  std_logic;
signal tile_55_X_c0 :  std_logic_vector(2 downto 0);
signal tile_55_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_55_output_c0 :  std_logic_vector(4 downto 0);
signal tile_55_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w65_8_c0 :  std_logic;
signal bh7_w66_9_c0 :  std_logic;
signal bh7_w67_8_c0 :  std_logic;
signal bh7_w68_8_c0 :  std_logic;
signal bh7_w69_8_c0 :  std_logic;
signal tile_56_X_c0 :  std_logic_vector(0 downto 0);
signal tile_56_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_56_output_c0 :  std_logic_vector(0 downto 0);
signal tile_56_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w102_0_c0 :  std_logic;
signal tile_57_X_c0 :  std_logic_vector(3 downto 0);
signal tile_57_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_57_output_c0 :  std_logic_vector(3 downto 0);
signal tile_57_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w98_2_c0 :  std_logic;
signal bh7_w99_1_c0 :  std_logic;
signal bh7_w100_1_c0 :  std_logic;
signal bh7_w101_0_c0 :  std_logic;
signal tile_58_X_c0 :  std_logic_vector(3 downto 0);
signal tile_58_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_58_output_c0 :  std_logic_vector(3 downto 0);
signal tile_58_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w94_3_c0 :  std_logic;
signal bh7_w95_2_c0 :  std_logic;
signal bh7_w96_3_c0 :  std_logic;
signal bh7_w97_3_c0 :  std_logic;
signal tile_59_X_c0 :  std_logic_vector(3 downto 0);
signal tile_59_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_59_output_c0 :  std_logic_vector(3 downto 0);
signal tile_59_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w90_3_c0 :  std_logic;
signal bh7_w91_3_c0 :  std_logic;
signal bh7_w92_2_c0 :  std_logic;
signal bh7_w93_3_c0 :  std_logic;
signal tile_60_X_c0 :  std_logic_vector(3 downto 0);
signal tile_60_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_60_output_c0 :  std_logic_vector(3 downto 0);
signal tile_60_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w86_2_c0 :  std_logic;
signal bh7_w87_3_c0 :  std_logic;
signal bh7_w88_3_c0 :  std_logic;
signal bh7_w89_2_c0 :  std_logic;
signal tile_61_X_c0 :  std_logic_vector(1 downto 0);
signal tile_61_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_61_output_c0 :  std_logic_vector(3 downto 0);
signal tile_61_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w99_2_c0 :  std_logic;
signal bh7_w100_2_c0 :  std_logic;
signal bh7_w101_1_c0 :  std_logic;
signal bh7_w102_1_c0 :  std_logic;
signal tile_62_X_c0 :  std_logic_vector(2 downto 0);
signal tile_62_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_62_output_c0 :  std_logic_vector(4 downto 0);
signal tile_62_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_4_c0 :  std_logic;
signal bh7_w97_4_c0 :  std_logic;
signal bh7_w98_3_c0 :  std_logic;
signal bh7_w99_3_c0 :  std_logic;
signal bh7_w100_3_c0 :  std_logic;
signal tile_63_X_c0 :  std_logic_vector(2 downto 0);
signal tile_63_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_63_output_c0 :  std_logic_vector(4 downto 0);
signal tile_63_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_4_c0 :  std_logic;
signal bh7_w94_4_c0 :  std_logic;
signal bh7_w95_3_c0 :  std_logic;
signal bh7_w96_5_c0 :  std_logic;
signal bh7_w97_5_c0 :  std_logic;
signal tile_64_X_c0 :  std_logic_vector(2 downto 0);
signal tile_64_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_64_output_c0 :  std_logic_vector(4 downto 0);
signal tile_64_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_4_c0 :  std_logic;
signal bh7_w91_4_c0 :  std_logic;
signal bh7_w92_3_c0 :  std_logic;
signal bh7_w93_5_c0 :  std_logic;
signal bh7_w94_5_c0 :  std_logic;
signal tile_65_X_c0 :  std_logic_vector(2 downto 0);
signal tile_65_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_65_output_c0 :  std_logic_vector(4 downto 0);
signal tile_65_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_4_c0 :  std_logic;
signal bh7_w88_4_c0 :  std_logic;
signal bh7_w89_3_c0 :  std_logic;
signal bh7_w90_5_c0 :  std_logic;
signal bh7_w91_5_c0 :  std_logic;
signal tile_66_X_c0 :  std_logic_vector(2 downto 0);
signal tile_66_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_66_output_c0 :  std_logic_vector(4 downto 0);
signal tile_66_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_5_c0 :  std_logic;
signal bh7_w85_5_c0 :  std_logic;
signal bh7_w86_3_c0 :  std_logic;
signal bh7_w87_5_c0 :  std_logic;
signal bh7_w88_5_c0 :  std_logic;
signal tile_67_X_c0 :  std_logic_vector(1 downto 0);
signal tile_67_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_67_output_c0 :  std_logic_vector(3 downto 0);
signal tile_67_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w97_6_c0 :  std_logic;
signal bh7_w98_4_c0 :  std_logic;
signal bh7_w99_4_c0 :  std_logic;
signal bh7_w100_4_c0 :  std_logic;
signal tile_68_X_c0 :  std_logic_vector(2 downto 0);
signal tile_68_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_68_output_c0 :  std_logic_vector(4 downto 0);
signal tile_68_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w94_6_c0 :  std_logic;
signal bh7_w95_4_c0 :  std_logic;
signal bh7_w96_6_c0 :  std_logic;
signal bh7_w97_7_c0 :  std_logic;
signal bh7_w98_5_c0 :  std_logic;
signal tile_69_X_c0 :  std_logic_vector(2 downto 0);
signal tile_69_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_69_output_c0 :  std_logic_vector(4 downto 0);
signal tile_69_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w91_6_c0 :  std_logic;
signal bh7_w92_4_c0 :  std_logic;
signal bh7_w93_6_c0 :  std_logic;
signal bh7_w94_7_c0 :  std_logic;
signal bh7_w95_5_c0 :  std_logic;
signal tile_70_X_c0 :  std_logic_vector(2 downto 0);
signal tile_70_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_70_output_c0 :  std_logic_vector(4 downto 0);
signal tile_70_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w88_6_c0 :  std_logic;
signal bh7_w89_4_c0 :  std_logic;
signal bh7_w90_6_c0 :  std_logic;
signal bh7_w91_7_c0 :  std_logic;
signal bh7_w92_5_c0 :  std_logic;
signal tile_71_X_c0 :  std_logic_vector(2 downto 0);
signal tile_71_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_71_output_c0 :  std_logic_vector(4 downto 0);
signal tile_71_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w85_6_c0 :  std_logic;
signal bh7_w86_4_c0 :  std_logic;
signal bh7_w87_6_c0 :  std_logic;
signal bh7_w88_7_c0 :  std_logic;
signal bh7_w89_5_c0 :  std_logic;
signal tile_72_X_c0 :  std_logic_vector(2 downto 0);
signal tile_72_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_72_output_c0 :  std_logic_vector(4 downto 0);
signal tile_72_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w82_7_c0 :  std_logic;
signal bh7_w83_6_c0 :  std_logic;
signal bh7_w84_6_c0 :  std_logic;
signal bh7_w85_7_c0 :  std_logic;
signal bh7_w86_5_c0 :  std_logic;
signal tile_73_X_c0 :  std_logic_vector(1 downto 0);
signal tile_73_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_73_output_c0 :  std_logic_vector(3 downto 0);
signal tile_73_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w102_2_c0 :  std_logic;
signal bh7_w103_0_c0 :  std_logic;
signal bh7_w104_0_c0 :  std_logic;
signal bh7_w105_0_c0 :  std_logic;
signal tile_74_X_c0 :  std_logic_vector(1 downto 0);
signal tile_74_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_74_output_c0 :  std_logic_vector(4 downto 0);
signal tile_74_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w99_5_c0 :  std_logic;
signal bh7_w100_5_c0 :  std_logic;
signal bh7_w101_2_c0 :  std_logic;
signal bh7_w102_3_c0 :  std_logic;
signal bh7_w103_1_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid323_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid323_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w49_5_c0 :  std_logic;
signal bh7_w50_6_c0 :  std_logic;
signal bh7_w51_8_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_copy324_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid327_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid327_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w51_9_c0 :  std_logic;
signal bh7_w52_9_c0 :  std_logic;
signal bh7_w53_9_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_copy328_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid329_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid329_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w52_10_c0 :  std_logic;
signal bh7_w53_10_c0 :  std_logic;
signal bh7_w54_11_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_copy330_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid331_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid331_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w53_11_c0 :  std_logic;
signal bh7_w54_12_c0 :  std_logic;
signal bh7_w55_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_copy332_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid335_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w54_13_c0 :  std_logic;
signal bh7_w55_11_c0 :  std_logic;
signal bh7_w56_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_copy336_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid337_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w55_12_c0 :  std_logic;
signal bh7_w56_10_c0 :  std_logic;
signal bh7_w57_11_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_copy338_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid339_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid339_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w56_11_c0 :  std_logic;
signal bh7_w57_12_c0 :  std_logic;
signal bh7_w58_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_copy340_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid341_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w57_13_c0 :  std_logic;
signal bh7_w58_11_c0 :  std_logic;
signal bh7_w59_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_copy342_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid343_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w58_12_c0 :  std_logic;
signal bh7_w59_10_c0 :  std_logic;
signal bh7_w60_11_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_copy344_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid345_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid345_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w59_11_c0 :  std_logic;
signal bh7_w60_12_c0 :  std_logic;
signal bh7_w61_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_copy346_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid347_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w60_13_c0 :  std_logic;
signal bh7_w61_11_c0 :  std_logic;
signal bh7_w62_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_copy348_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid349_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w61_12_c0 :  std_logic;
signal bh7_w62_10_c0 :  std_logic;
signal bh7_w63_11_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_copy350_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid351_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid351_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w62_11_c0 :  std_logic;
signal bh7_w63_12_c0 :  std_logic;
signal bh7_w64_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_copy352_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid353_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w63_13_c0 :  std_logic;
signal bh7_w64_11_c0 :  std_logic;
signal bh7_w65_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_copy354_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid355_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w64_12_c0 :  std_logic;
signal bh7_w65_10_c0 :  std_logic;
signal bh7_w66_10_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_copy356_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid357_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w65_11_c0 :  std_logic;
signal bh7_w66_11_c0 :  std_logic;
signal bh7_w67_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_copy358_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid359_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_12_c0 :  std_logic;
signal bh7_w67_10_c0 :  std_logic;
signal bh7_w68_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_copy360_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid361_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w67_11_c0 :  std_logic;
signal bh7_w68_10_c0 :  std_logic;
signal bh7_w69_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_copy362_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid363_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_11_c0 :  std_logic;
signal bh7_w69_10_c0 :  std_logic;
signal bh7_w70_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_copy364_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid365_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w69_11_c0 :  std_logic;
signal bh7_w70_10_c0 :  std_logic;
signal bh7_w71_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_copy366_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid367_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_11_c0 :  std_logic;
signal bh7_w71_10_c0 :  std_logic;
signal bh7_w72_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_copy368_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid369_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w71_11_c0 :  std_logic;
signal bh7_w72_10_c0 :  std_logic;
signal bh7_w73_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_copy370_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid371_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_11_c0 :  std_logic;
signal bh7_w73_10_c0 :  std_logic;
signal bh7_w74_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_copy372_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid373_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w73_11_c0 :  std_logic;
signal bh7_w74_10_c0 :  std_logic;
signal bh7_w75_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_copy374_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid375_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_11_c0 :  std_logic;
signal bh7_w75_9_c0 :  std_logic;
signal bh7_w76_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_copy376_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid377_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w75_10_c0 :  std_logic;
signal bh7_w76_9_c0 :  std_logic;
signal bh7_w77_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_copy378_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid379_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_10_c0 :  std_logic;
signal bh7_w77_9_c0 :  std_logic;
signal bh7_w78_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_copy380_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid381_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w77_10_c0 :  std_logic;
signal bh7_w78_9_c0 :  std_logic;
signal bh7_w79_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_copy382_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid383_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_10_c0 :  std_logic;
signal bh7_w79_9_c0 :  std_logic;
signal bh7_w80_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_copy384_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid385_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w79_10_c0 :  std_logic;
signal bh7_w80_9_c0 :  std_logic;
signal bh7_w81_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_copy386_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid387_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_10_c0 :  std_logic;
signal bh7_w81_9_c0 :  std_logic;
signal bh7_w82_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_copy388_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid389_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w81_10_c0 :  std_logic;
signal bh7_w82_9_c0 :  std_logic;
signal bh7_w83_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_copy390_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid391_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_10_c0 :  std_logic;
signal bh7_w83_8_c0 :  std_logic;
signal bh7_w84_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_copy392_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid393_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w83_9_c0 :  std_logic;
signal bh7_w84_8_c0 :  std_logic;
signal bh7_w85_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_copy394_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid395_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w84_9_c0 :  std_logic;
signal bh7_w85_9_c0 :  std_logic;
signal bh7_w86_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_copy396_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid397_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w85_10_c0 :  std_logic;
signal bh7_w86_7_c0 :  std_logic;
signal bh7_w87_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_copy398_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid401_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w86_8_c0 :  std_logic;
signal bh7_w87_8_c0 :  std_logic;
signal bh7_w88_8_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_copy402_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid403_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w87_9_c0 :  std_logic;
signal bh7_w88_9_c0 :  std_logic;
signal bh7_w89_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_copy404_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid405_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w88_10_c0 :  std_logic;
signal bh7_w89_7_c0 :  std_logic;
signal bh7_w90_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_copy406_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid407_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w89_8_c0 :  std_logic;
signal bh7_w90_8_c0 :  std_logic;
signal bh7_w91_8_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_copy408_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid409_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w90_9_c0 :  std_logic;
signal bh7_w91_9_c0 :  std_logic;
signal bh7_w92_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_copy410_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid411_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w91_10_c0 :  std_logic;
signal bh7_w92_7_c0 :  std_logic;
signal bh7_w93_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_copy412_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid413_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w92_8_c0 :  std_logic;
signal bh7_w93_8_c0 :  std_logic;
signal bh7_w94_8_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_copy414_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid415_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w93_9_c0 :  std_logic;
signal bh7_w94_9_c0 :  std_logic;
signal bh7_w95_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_copy416_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid417_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w94_10_c0 :  std_logic;
signal bh7_w95_7_c0 :  std_logic;
signal bh7_w96_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_copy418_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid419_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w95_8_c0 :  std_logic;
signal bh7_w96_8_c0 :  std_logic;
signal bh7_w97_8_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_copy420_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid421_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w96_9_c0 :  std_logic;
signal bh7_w97_9_c0 :  std_logic;
signal bh7_w98_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_copy422_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid423_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w97_10_c0 :  std_logic;
signal bh7_w98_7_c0 :  std_logic;
signal bh7_w99_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_copy424_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid425_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w98_8_c0 :  std_logic;
signal bh7_w99_7_c0 :  std_logic;
signal bh7_w100_6_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_copy426_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid427_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w99_8_c0 :  std_logic;
signal bh7_w100_7_c0 :  std_logic;
signal bh7_w101_3_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_copy428_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid429_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w100_8_c0 :  std_logic;
signal bh7_w101_4_c0 :  std_logic;
signal bh7_w102_4_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_copy430_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid433_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w101_5_c0 :  std_logic;
signal bh7_w102_5_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_copy434_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid435_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid435_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w102_6_c0 :  std_logic;
signal bh7_w103_2_c0 :  std_logic;
signal bh7_w104_1_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_copy436_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid437_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid437_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w51_10_c0 :  std_logic;
signal bh7_w52_11_c0 :  std_logic;
signal bh7_w53_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_copy438_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid439_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid439_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w53_13_c0 :  std_logic;
signal bh7_w54_14_c0 :  std_logic;
signal bh7_w55_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_copy440_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid441_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w55_14_c0 :  std_logic;
signal bh7_w56_12_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_copy442_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid443_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid443_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w56_13_c0 :  std_logic;
signal bh7_w57_14_c0 :  std_logic;
signal bh7_w58_13_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_copy444_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid445_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w57_15_c0 :  std_logic;
signal bh7_w58_14_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_copy446_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid447_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w58_15_c0 :  std_logic;
signal bh7_w59_12_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_copy448_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid449_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid449_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w59_13_c0 :  std_logic;
signal bh7_w60_14_c0 :  std_logic;
signal bh7_w61_13_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_copy450_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid451_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w60_15_c0 :  std_logic;
signal bh7_w61_14_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_copy452_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid453_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w61_15_c0 :  std_logic;
signal bh7_w62_12_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_copy454_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid455_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid455_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w62_13_c0 :  std_logic;
signal bh7_w63_14_c0 :  std_logic;
signal bh7_w64_13_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_copy456_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid457_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w63_15_c0 :  std_logic;
signal bh7_w64_14_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_copy458_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid459_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid459_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w64_15_c0 :  std_logic;
signal bh7_w65_12_c0 :  std_logic;
signal bh7_w66_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_copy460_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid461_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid461_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_14_c0 :  std_logic;
signal bh7_w67_12_c0 :  std_logic;
signal bh7_w68_12_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_copy462_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid463_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w67_13_c0 :  std_logic;
signal bh7_w68_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_copy464_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid465_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid465_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_14_c0 :  std_logic;
signal bh7_w69_12_c0 :  std_logic;
signal bh7_w70_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_copy466_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid467_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid467_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_13_c0 :  std_logic;
signal bh7_w71_12_c0 :  std_logic;
signal bh7_w72_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_copy468_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid469_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid469_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_13_c0 :  std_logic;
signal bh7_w73_12_c0 :  std_logic;
signal bh7_w74_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_copy470_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid471_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid471_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_13_c0 :  std_logic;
signal bh7_w75_11_c0 :  std_logic;
signal bh7_w76_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_copy472_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid473_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid473_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_12_c0 :  std_logic;
signal bh7_w77_11_c0 :  std_logic;
signal bh7_w78_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_copy474_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid475_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid475_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_12_c0 :  std_logic;
signal bh7_w79_11_c0 :  std_logic;
signal bh7_w80_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_copy476_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid477_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid477_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_12_c0 :  std_logic;
signal bh7_w81_11_c0 :  std_logic;
signal bh7_w82_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_copy478_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid479_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid479_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_12_c0 :  std_logic;
signal bh7_w83_10_c0 :  std_logic;
signal bh7_w84_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_copy480_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid481_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w83_11_c0 :  std_logic;
signal bh7_w84_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_copy482_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid483_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w84_12_c0 :  std_logic;
signal bh7_w85_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_copy484_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid485_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid485_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w85_12_c0 :  std_logic;
signal bh7_w86_9_c0 :  std_logic;
signal bh7_w87_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_copy486_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid487_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w86_10_c0 :  std_logic;
signal bh7_w87_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_copy488_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid489_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w87_12_c0 :  std_logic;
signal bh7_w88_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_copy490_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid491_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid491_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w88_12_c0 :  std_logic;
signal bh7_w89_9_c0 :  std_logic;
signal bh7_w90_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_copy492_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid493_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w89_10_c0 :  std_logic;
signal bh7_w90_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_copy494_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid495_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w90_12_c0 :  std_logic;
signal bh7_w91_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_copy496_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid497_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid497_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w91_12_c0 :  std_logic;
signal bh7_w92_9_c0 :  std_logic;
signal bh7_w93_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_copy498_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid499_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w92_10_c0 :  std_logic;
signal bh7_w93_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_copy500_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid501_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w93_12_c0 :  std_logic;
signal bh7_w94_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_copy502_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid503_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid503_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w94_12_c0 :  std_logic;
signal bh7_w95_9_c0 :  std_logic;
signal bh7_w96_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_copy504_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid505_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w95_10_c0 :  std_logic;
signal bh7_w96_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_copy506_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid507_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w96_12_c0 :  std_logic;
signal bh7_w97_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_copy508_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid509_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid509_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w97_12_c0 :  std_logic;
signal bh7_w98_9_c0 :  std_logic;
signal bh7_w99_9_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_copy510_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid511_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w98_10_c0 :  std_logic;
signal bh7_w99_10_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_copy512_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid513_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid513_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w99_11_c0 :  std_logic;
signal bh7_w100_9_c0 :  std_logic;
signal bh7_w101_6_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_copy514_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid515_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid515_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w101_7_c0 :  std_logic;
signal bh7_w102_7_c0 :  std_logic;
signal bh7_w103_3_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_copy516_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid517_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid517_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w103_4_c0 :  std_logic;
signal bh7_w104_2_c0 :  std_logic;
signal bh7_w105_1_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_copy518_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid519_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid519_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w53_14_c0 :  std_logic;
signal bh7_w54_15_c0 :  std_logic;
signal bh7_w55_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_copy520_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid521_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid521_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w55_16_c0 :  std_logic;
signal bh7_w56_14_c0 :  std_logic;
signal bh7_w57_16_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_copy522_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid523_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w57_17_c0 :  std_logic;
signal bh7_w58_16_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_copy524_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid525_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid525_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w58_17_c0 :  std_logic;
signal bh7_w59_14_c0 :  std_logic;
signal bh7_w60_16_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_copy526_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid527_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w60_17_c0 :  std_logic;
signal bh7_w61_16_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_copy528_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid529_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid529_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w61_17_c0 :  std_logic;
signal bh7_w62_14_c0 :  std_logic;
signal bh7_w63_16_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_copy530_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid531_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w63_17_c0 :  std_logic;
signal bh7_w64_16_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_copy532_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid533_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid533_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w64_17_c0 :  std_logic;
signal bh7_w65_13_c0 :  std_logic;
signal bh7_w66_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_copy534_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid535_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid535_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_16_c0 :  std_logic;
signal bh7_w67_14_c0 :  std_logic;
signal bh7_w68_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_copy536_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid537_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid537_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_16_c0 :  std_logic;
signal bh7_w69_13_c0 :  std_logic;
signal bh7_w70_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_copy538_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid539_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid539_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_15_c0 :  std_logic;
signal bh7_w71_13_c0 :  std_logic;
signal bh7_w72_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_copy540_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid541_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid541_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_15_c0 :  std_logic;
signal bh7_w73_13_c0 :  std_logic;
signal bh7_w74_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_copy542_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid543_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid543_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_15_c0 :  std_logic;
signal bh7_w75_12_c0 :  std_logic;
signal bh7_w76_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_copy544_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid545_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid545_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_14_c0 :  std_logic;
signal bh7_w77_12_c0 :  std_logic;
signal bh7_w78_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_copy546_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid547_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid547_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_14_c0 :  std_logic;
signal bh7_w79_12_c0 :  std_logic;
signal bh7_w80_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_copy548_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid549_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid549_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_14_c0 :  std_logic;
signal bh7_w81_12_c0 :  std_logic;
signal bh7_w82_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_copy550_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid551_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid551_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_14_c0 :  std_logic;
signal bh7_w83_12_c0 :  std_logic;
signal bh7_w84_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_copy552_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid553_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid553_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w84_14_c0 :  std_logic;
signal bh7_w85_13_c0 :  std_logic;
signal bh7_w86_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_copy554_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid555_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w86_12_c0 :  std_logic;
signal bh7_w87_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_copy556_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid557_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid557_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w87_14_c0 :  std_logic;
signal bh7_w88_13_c0 :  std_logic;
signal bh7_w89_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_copy558_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid559_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w89_12_c0 :  std_logic;
signal bh7_w90_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_copy560_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid561_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid561_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w90_14_c0 :  std_logic;
signal bh7_w91_13_c0 :  std_logic;
signal bh7_w92_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_copy562_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid563_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w92_12_c0 :  std_logic;
signal bh7_w93_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_copy564_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid565_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid565_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w93_14_c0 :  std_logic;
signal bh7_w94_13_c0 :  std_logic;
signal bh7_w95_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_copy566_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid567_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w95_12_c0 :  std_logic;
signal bh7_w96_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_copy568_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid569_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid569_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w96_14_c0 :  std_logic;
signal bh7_w97_13_c0 :  std_logic;
signal bh7_w98_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_copy570_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid571_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w98_12_c0 :  std_logic;
signal bh7_w99_12_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_copy572_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid573_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid573_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w99_13_c0 :  std_logic;
signal bh7_w100_10_c0 :  std_logic;
signal bh7_w101_8_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_copy574_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid575_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid575_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w101_9_c0 :  std_logic;
signal bh7_w102_8_c0 :  std_logic;
signal bh7_w103_5_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_copy576_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid577_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid577_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w103_6_c0 :  std_logic;
signal bh7_w104_3_c0 :  std_logic;
signal bh7_w105_2_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_copy578_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid579_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w105_3_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_copy580_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid581_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid581_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w55_17_c0 :  std_logic;
signal bh7_w56_15_c0 :  std_logic;
signal bh7_w57_18_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_copy582_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid583_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid583_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w57_19_c0 :  std_logic;
signal bh7_w58_18_c0 :  std_logic;
signal bh7_w59_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_copy584_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid585_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid585_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w60_18_c0 :  std_logic;
signal bh7_w61_18_c0, bh7_w61_18_c1 :  std_logic;
signal bh7_w62_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_copy586_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid587_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid587_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w63_18_c0 :  std_logic;
signal bh7_w64_18_c0, bh7_w64_18_c1 :  std_logic;
signal bh7_w65_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_copy588_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid589_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid589_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_17_c0 :  std_logic;
signal bh7_w67_15_c0, bh7_w67_15_c1 :  std_logic;
signal bh7_w68_17_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_copy590_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid591_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid591_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_18_c0 :  std_logic;
signal bh7_w69_14_c0 :  std_logic;
signal bh7_w70_16_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_copy592_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid593_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid593_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_17_c0 :  std_logic;
signal bh7_w71_14_c0 :  std_logic;
signal bh7_w72_16_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_copy594_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid595_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid595_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_17_c0 :  std_logic;
signal bh7_w73_14_c0 :  std_logic;
signal bh7_w74_16_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_copy596_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid597_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid597_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_17_c0 :  std_logic;
signal bh7_w75_13_c0 :  std_logic;
signal bh7_w76_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_copy598_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid599_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid599_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_16_c0 :  std_logic;
signal bh7_w77_13_c0 :  std_logic;
signal bh7_w78_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_copy600_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid601_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid601_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_16_c0 :  std_logic;
signal bh7_w79_13_c0 :  std_logic;
signal bh7_w80_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_copy602_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid603_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid603_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_16_c0 :  std_logic;
signal bh7_w81_13_c0 :  std_logic;
signal bh7_w82_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_copy604_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid605_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid605_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_16_c0 :  std_logic;
signal bh7_w83_13_c0 :  std_logic;
signal bh7_w84_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_copy606_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid607_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid607_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w84_16_c0 :  std_logic;
signal bh7_w85_14_c0 :  std_logic;
signal bh7_w86_13_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_copy608_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid609_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid609_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w86_14_c0 :  std_logic;
signal bh7_w87_15_c0 :  std_logic;
signal bh7_w88_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_copy610_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid611_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid611_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w89_13_c0 :  std_logic;
signal bh7_w90_15_c0, bh7_w90_15_c1 :  std_logic;
signal bh7_w91_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_copy612_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid613_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid613_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w92_13_c0 :  std_logic;
signal bh7_w93_15_c0, bh7_w93_15_c1 :  std_logic;
signal bh7_w94_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_copy614_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid615_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid615_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w95_13_c0 :  std_logic;
signal bh7_w96_15_c0, bh7_w96_15_c1 :  std_logic;
signal bh7_w97_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_copy616_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid617_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid617_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w98_13_c0 :  std_logic;
signal bh7_w99_14_c0, bh7_w99_14_c1 :  std_logic;
signal bh7_w100_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_copy618_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid619_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid619_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w101_10_c0 :  std_logic;
signal bh7_w102_9_c0, bh7_w102_9_c1 :  std_logic;
signal bh7_w103_7_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_copy620_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid621_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid621_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w103_8_c0 :  std_logic;
signal bh7_w104_4_c0 :  std_logic;
signal bh7_w105_4_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_copy622_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid623_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid623_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w105_5_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_copy624_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid625_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid625_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w57_20_c1 :  std_logic;
signal bh7_w58_19_c1 :  std_logic;
signal bh7_w59_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c0, Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid627_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid627_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_17_c1 :  std_logic;
signal bh7_w60_19_c1 :  std_logic;
signal bh7_w61_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c0, Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid629_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid629_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_16_c1 :  std_logic;
signal bh7_w63_19_c1 :  std_logic;
signal bh7_w64_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c0, Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid631_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid631_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w65_15_c1 :  std_logic;
signal bh7_w66_18_c1 :  std_logic;
signal bh7_w67_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c0, Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid633_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid633_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_19_c1 :  std_logic;
signal bh7_w69_15_c1 :  std_logic;
signal bh7_w70_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c0, Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid635_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid635_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_19_c1 :  std_logic;
signal bh7_w71_15_c1 :  std_logic;
signal bh7_w72_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c0, Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid637_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid637_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_19_c1 :  std_logic;
signal bh7_w73_15_c1 :  std_logic;
signal bh7_w74_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c0, Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid639_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid639_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_19_c1 :  std_logic;
signal bh7_w75_14_c1 :  std_logic;
signal bh7_w76_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c0, Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid641_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid641_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_18_c1 :  std_logic;
signal bh7_w77_14_c1 :  std_logic;
signal bh7_w78_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c0, Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid643_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid643_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_18_c1 :  std_logic;
signal bh7_w79_14_c1 :  std_logic;
signal bh7_w80_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c0, Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid645_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid645_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_18_c1 :  std_logic;
signal bh7_w81_14_c1 :  std_logic;
signal bh7_w82_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c0, Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid647_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid647_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_18_c1 :  std_logic;
signal bh7_w83_14_c1 :  std_logic;
signal bh7_w84_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c0, Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid649_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid649_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_18_c1 :  std_logic;
signal bh7_w85_15_c1 :  std_logic;
signal bh7_w86_15_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c0, Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid651_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid651_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_16_c1 :  std_logic;
signal bh7_w87_16_c1 :  std_logic;
signal bh7_w88_15_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c0, Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid653_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid653_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_16_c1 :  std_logic;
signal bh7_w89_14_c1 :  std_logic;
signal bh7_w90_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c0, Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid655_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid655_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w91_15_c1 :  std_logic;
signal bh7_w92_14_c1 :  std_logic;
signal bh7_w93_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c0, Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid657_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid657_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w94_15_c1 :  std_logic;
signal bh7_w95_14_c1 :  std_logic;
signal bh7_w96_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c0, Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid659_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid659_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w97_15_c1 :  std_logic;
signal bh7_w98_14_c1 :  std_logic;
signal bh7_w99_15_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c0, Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid661_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid661_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w100_12_c1 :  std_logic;
signal bh7_w101_11_c1 :  std_logic;
signal bh7_w102_10_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c0, Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid663_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid663_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w103_9_c1 :  std_logic;
signal bh7_w104_5_c1 :  std_logic;
signal bh7_w105_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c0, Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid665_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid665_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w105_7_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c0, Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid667_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid667_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w17_2_c1 :  std_logic;
signal bh7_w18_2_c1 :  std_logic;
signal bh7_w19_2_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c0, Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid669_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid669_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w19_3_c1 :  std_logic;
signal bh7_w20_2_c1 :  std_logic;
signal bh7_w21_2_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c0, Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid671_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid671_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_3_c1 :  std_logic;
signal bh7_w22_2_c1 :  std_logic;
signal bh7_w23_2_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c0, Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid673_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w23_3_c1 :  std_logic;
signal bh7_w24_3_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c0, Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid675_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid675_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w24_4_c1 :  std_logic;
signal bh7_w25_3_c1 :  std_logic;
signal bh7_w26_3_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c0, Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid677_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid677_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w26_4_c1 :  std_logic;
signal bh7_w27_3_c1 :  std_logic;
signal bh7_w28_3_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c0, Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid679_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid679_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w28_4_c1 :  std_logic;
signal bh7_w29_3_c1 :  std_logic;
signal bh7_w30_3_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c0, Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid681_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid681_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w30_4_c1 :  std_logic;
signal bh7_w31_3_c1 :  std_logic;
signal bh7_w32_3_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c0, Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid683_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid683_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w32_4_c1 :  std_logic;
signal bh7_w33_3_c1 :  std_logic;
signal bh7_w34_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c0, Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid685_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid685_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w34_5_c1 :  std_logic;
signal bh7_w35_4_c1 :  std_logic;
signal bh7_w36_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c0, Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid687_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w35_5_c1 :  std_logic;
signal bh7_w36_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c0, Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid689_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid689_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w36_6_c1 :  std_logic;
signal bh7_w37_4_c1 :  std_logic;
signal bh7_w38_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c0, Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid691_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w37_5_c1 :  std_logic;
signal bh7_w38_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c0, Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid693_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid693_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w38_6_c1 :  std_logic;
signal bh7_w39_4_c1 :  std_logic;
signal bh7_w40_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c0, Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid695_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w39_5_c1 :  std_logic;
signal bh7_w40_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c0, Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid697_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid697_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w40_6_c1 :  std_logic;
signal bh7_w41_4_c1 :  std_logic;
signal bh7_w42_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c0, Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid699_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w41_5_c1 :  std_logic;
signal bh7_w42_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c0, Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid701_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid701_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w42_6_c1 :  std_logic;
signal bh7_w43_4_c1 :  std_logic;
signal bh7_w44_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c0, Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid703_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w43_5_c1 :  std_logic;
signal bh7_w44_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c0, Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid705_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid705_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w44_6_c1 :  std_logic;
signal bh7_w45_4_c1 :  std_logic;
signal bh7_w46_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c0, Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid707_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w45_5_c1 :  std_logic;
signal bh7_w46_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c0, Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid709_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid709_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w46_6_c1 :  std_logic;
signal bh7_w47_4_c1 :  std_logic;
signal bh7_w48_5_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c0, Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid711_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w47_5_c1 :  std_logic;
signal bh7_w48_6_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c0, Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid713_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid713_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w48_7_c1 :  std_logic;
signal bh7_w49_6_c1 :  std_logic;
signal bh7_w50_7_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c0, Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid715_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid715_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w49_7_c1 :  std_logic;
signal bh7_w50_8_c1 :  std_logic;
signal bh7_w51_11_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c0, Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid717_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid717_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w50_9_c1 :  std_logic;
signal bh7_w51_12_c1 :  std_logic;
signal bh7_w52_12_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c0, Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid719_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid719_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w51_13_c1 :  std_logic;
signal bh7_w52_13_c1 :  std_logic;
signal bh7_w53_15_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c0, Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid721_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid721_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w52_14_c1 :  std_logic;
signal bh7_w53_16_c1 :  std_logic;
signal bh7_w54_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c0, Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid723_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid723_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w53_17_c1 :  std_logic;
signal bh7_w54_17_c1 :  std_logic;
signal bh7_w55_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c0, Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid725_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid725_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w54_18_c1 :  std_logic;
signal bh7_w55_19_c1 :  std_logic;
signal bh7_w56_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c0, Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid727_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid727_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w55_20_c1 :  std_logic;
signal bh7_w56_17_c1 :  std_logic;
signal bh7_w57_21_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c0, Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c0, Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid729_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_18_c1 :  std_logic;
signal bh7_w57_22_c1 :  std_logic;
signal bh7_w58_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_copy730_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c0, Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid731_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w57_23_c1 :  std_logic;
signal bh7_w58_21_c1 :  std_logic;
signal bh7_w59_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_copy732_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid733_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w58_22_c1 :  std_logic;
signal bh7_w59_19_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c0, Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c1 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid735_In0_c1 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_20_c1 :  std_logic;
signal bh7_w60_20_c1 :  std_logic;
signal bh7_w61_20_c1 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_copy736_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid737_In0_c1 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w60_21_c1 :  std_logic;
signal bh7_w61_21_c1 :  std_logic;
signal bh7_w62_17_c1 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_copy738_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid739_In0_c1 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w61_22_c1 :  std_logic;
signal bh7_w62_18_c1 :  std_logic;
signal bh7_w63_20_c1 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_copy740_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid741_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid741_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_19_c1 :  std_logic;
signal bh7_w63_21_c1 :  std_logic;
signal bh7_w64_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_copy742_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid743_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w63_22_c1 :  std_logic;
signal bh7_w64_21_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c0, Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c1 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid745_In0_c1 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_22_c1 :  std_logic;
signal bh7_w65_16_c1 :  std_logic;
signal bh7_w66_19_c1 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_copy746_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid747_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid747_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w65_17_c1 :  std_logic;
signal bh7_w66_20_c1 :  std_logic;
signal bh7_w67_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_copy748_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid749_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w66_21_c1 :  std_logic;
signal bh7_w67_18_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c0, Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid751_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid751_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w67_19_c1 :  std_logic;
signal bh7_w68_20_c1 :  std_logic;
signal bh7_w69_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_copy752_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid753_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w68_21_c1 :  std_logic;
signal bh7_w69_17_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c0, Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid755_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid755_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w69_18_c1 :  std_logic;
signal bh7_w70_20_c1 :  std_logic;
signal bh7_w71_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_copy756_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid757_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid757_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_21_c1 :  std_logic;
signal bh7_w71_17_c1 :  std_logic;
signal bh7_w72_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_copy758_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid759_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w71_18_c1 :  std_logic;
signal bh7_w72_21_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c0, Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid761_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid761_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_22_c1 :  std_logic;
signal bh7_w73_16_c1 :  std_logic;
signal bh7_w74_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_copy762_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid763_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w73_17_c1 :  std_logic;
signal bh7_w74_21_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c0, Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid765_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_22_c1 :  std_logic;
signal bh7_w75_15_c1 :  std_logic;
signal bh7_w76_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_copy766_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid767_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid767_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_23_c1 :  std_logic;
signal bh7_w75_16_c1 :  std_logic;
signal bh7_w76_20_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_copy768_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid769_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_21_c1 :  std_logic;
signal bh7_w77_15_c1 :  std_logic;
signal bh7_w78_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_copy770_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid771_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w77_16_c1 :  std_logic;
signal bh7_w78_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_copy772_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid773_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_21_c1 :  std_logic;
signal bh7_w79_15_c1 :  std_logic;
signal bh7_w80_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_copy774_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid775_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w79_16_c1 :  std_logic;
signal bh7_w80_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_copy776_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid777_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_21_c1 :  std_logic;
signal bh7_w81_15_c1 :  std_logic;
signal bh7_w82_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_copy778_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid779_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w81_16_c1 :  std_logic;
signal bh7_w82_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_copy780_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid781_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid781_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_21_c1 :  std_logic;
signal bh7_w83_15_c1 :  std_logic;
signal bh7_w84_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_copy782_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid783_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid783_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_20_c1 :  std_logic;
signal bh7_w85_16_c1 :  std_logic;
signal bh7_w86_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_copy784_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid785_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid785_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_18_c1 :  std_logic;
signal bh7_w87_17_c1 :  std_logic;
signal bh7_w88_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_copy786_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid787_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid787_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_18_c1 :  std_logic;
signal bh7_w89_15_c1 :  std_logic;
signal bh7_w90_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_copy788_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid789_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid789_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w90_18_c1 :  std_logic;
signal bh7_w91_16_c1 :  std_logic;
signal bh7_w92_15_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_copy790_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid791_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w92_16_c1 :  std_logic;
signal bh7_w93_17_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_copy792_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid793_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid793_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w93_18_c1 :  std_logic;
signal bh7_w94_16_c1 :  std_logic;
signal bh7_w95_15_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_copy794_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid795_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w95_16_c1 :  std_logic;
signal bh7_w96_17_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_copy796_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid797_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid797_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w96_18_c1 :  std_logic;
signal bh7_w97_16_c1 :  std_logic;
signal bh7_w98_15_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_copy798_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid799_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid799_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w98_16_c1 :  std_logic;
signal bh7_w99_16_c1 :  std_logic;
signal bh7_w100_13_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_copy800_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid801_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid801_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w102_11_c1 :  std_logic;
signal bh7_w103_10_c1 :  std_logic;
signal bh7_w104_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_copy802_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid803_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w105_8_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_copy804_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid805_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid805_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w19_4_c1 :  std_logic;
signal bh7_w20_3_c1 :  std_logic;
signal bh7_w21_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_copy806_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid807_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid807_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_5_c1 :  std_logic;
signal bh7_w22_3_c1 :  std_logic;
signal bh7_w23_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_copy808_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid809_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid809_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w23_5_c1 :  std_logic;
signal bh7_w24_5_c1 :  std_logic;
signal bh7_w25_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_copy810_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid811_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid811_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w25_5_c1 :  std_logic;
signal bh7_w26_5_c1 :  std_logic;
signal bh7_w27_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_copy812_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid813_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid813_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w27_5_c1 :  std_logic;
signal bh7_w28_5_c1 :  std_logic;
signal bh7_w29_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_copy814_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid815_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid815_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_5_c1 :  std_logic;
signal bh7_w30_5_c1 :  std_logic;
signal bh7_w31_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_copy816_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid817_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid817_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_5_c1 :  std_logic;
signal bh7_w32_5_c1 :  std_logic;
signal bh7_w33_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_copy818_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid819_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid819_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_5_c1 :  std_logic;
signal bh7_w34_6_c1 :  std_logic;
signal bh7_w35_6_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_copy820_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid821_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w35_7_c1 :  std_logic;
signal bh7_w36_7_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_copy822_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid823_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid823_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w36_8_c1 :  std_logic;
signal bh7_w37_6_c1 :  std_logic;
signal bh7_w38_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_copy824_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid825_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid825_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w38_8_c1 :  std_logic;
signal bh7_w39_6_c1 :  std_logic;
signal bh7_w40_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_copy826_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid827_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid827_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w40_8_c1 :  std_logic;
signal bh7_w41_6_c1 :  std_logic;
signal bh7_w42_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_copy828_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid829_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid829_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w42_8_c1 :  std_logic;
signal bh7_w43_6_c1 :  std_logic;
signal bh7_w44_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_copy830_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid831_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid831_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w44_8_c1 :  std_logic;
signal bh7_w45_6_c1 :  std_logic;
signal bh7_w46_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_copy832_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid833_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid833_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w46_8_c1 :  std_logic;
signal bh7_w47_6_c1 :  std_logic;
signal bh7_w48_8_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_copy834_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid835_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid835_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w48_9_c1 :  std_logic;
signal bh7_w49_8_c1 :  std_logic;
signal bh7_w50_10_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_copy836_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid837_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid837_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w50_11_c1 :  std_logic;
signal bh7_w51_14_c1 :  std_logic;
signal bh7_w52_15_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_copy838_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid839_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid839_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w52_16_c1 :  std_logic;
signal bh7_w53_18_c1 :  std_logic;
signal bh7_w54_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_copy840_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid841_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid841_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w54_20_c1 :  std_logic;
signal bh7_w55_21_c1 :  std_logic;
signal bh7_w56_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_copy842_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid843_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid843_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_20_c1 :  std_logic;
signal bh7_w57_24_c1 :  std_logic;
signal bh7_w58_23_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_copy844_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid845_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w58_24_c1 :  std_logic;
signal bh7_w59_21_c1 :  std_logic;
signal bh7_w60_22_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_copy846_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid847_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid847_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_22_c1 :  std_logic;
signal bh7_w60_23_c1 :  std_logic;
signal bh7_w61_23_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_copy848_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid849_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w61_24_c1 :  std_logic;
signal bh7_w62_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_copy850_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid851_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid851_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_21_c1 :  std_logic;
signal bh7_w63_23_c1 :  std_logic;
signal bh7_w64_23_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_copy852_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid853_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c0, Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w63_24_c1 :  std_logic;
signal bh7_w64_24_c1 :  std_logic;
signal bh7_w65_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_copy854_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid855_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid855_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_25_c1 :  std_logic;
signal bh7_w65_19_c1 :  std_logic;
signal bh7_w66_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_copy856_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid857_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w66_23_c1 :  std_logic;
signal bh7_w67_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_copy858_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid859_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid859_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w67_21_c1 :  std_logic;
signal bh7_w68_22_c1 :  std_logic;
signal bh7_w69_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_copy860_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid861_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid861_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w69_20_c1 :  std_logic;
signal bh7_w70_22_c1 :  std_logic;
signal bh7_w71_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_copy862_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid863_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w71_20_c1 :  std_logic;
signal bh7_w72_23_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_copy864_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid865_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid865_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_24_c1 :  std_logic;
signal bh7_w73_18_c1 :  std_logic;
signal bh7_w74_24_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_copy866_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid867_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid867_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_25_c1 :  std_logic;
signal bh7_w75_17_c1 :  std_logic;
signal bh7_w76_22_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_copy868_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid869_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid869_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_23_c1 :  std_logic;
signal bh7_w77_17_c1 :  std_logic;
signal bh7_w78_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_copy870_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid871_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid871_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_23_c1 :  std_logic;
signal bh7_w79_17_c1 :  std_logic;
signal bh7_w80_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_copy872_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid873_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid873_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_23_c1 :  std_logic;
signal bh7_w81_17_c1 :  std_logic;
signal bh7_w82_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_copy874_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid875_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w82_23_c1 :  std_logic;
signal bh7_w83_16_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_copy876_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid877_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid877_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_21_c1 :  std_logic;
signal bh7_w85_17_c1 :  std_logic;
signal bh7_w86_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_copy878_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid879_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid879_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_20_c1 :  std_logic;
signal bh7_w87_18_c1 :  std_logic;
signal bh7_w88_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_copy880_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid881_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid881_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_20_c1 :  std_logic;
signal bh7_w89_16_c1 :  std_logic;
signal bh7_w90_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_copy882_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid883_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid883_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w90_20_c1 :  std_logic;
signal bh7_w91_17_c1 :  std_logic;
signal bh7_w92_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_copy884_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid885_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid885_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w92_18_c1 :  std_logic;
signal bh7_w93_19_c1 :  std_logic;
signal bh7_w94_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_copy886_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid887_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid887_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w95_17_c1 :  std_logic;
signal bh7_w96_19_c1 :  std_logic;
signal bh7_w97_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_copy888_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid889_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid889_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w98_17_c1 :  std_logic;
signal bh7_w99_17_c1 :  std_logic;
signal bh7_w100_14_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_copy890_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid891_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid891_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w100_15_c1 :  std_logic;
signal bh7_w101_12_c1 :  std_logic;
signal bh7_w102_12_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_copy892_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid893_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid893_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w104_7_c1 :  std_logic;
signal bh7_w105_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_copy894_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid895_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid895_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_6_c1 :  std_logic;
signal bh7_w22_4_c1 :  std_logic;
signal bh7_w23_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_copy896_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid897_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid897_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w23_7_c1 :  std_logic;
signal bh7_w24_6_c1 :  std_logic;
signal bh7_w25_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_copy898_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid899_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid899_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w25_7_c1 :  std_logic;
signal bh7_w26_6_c1 :  std_logic;
signal bh7_w27_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_copy900_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid901_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid901_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w27_7_c1 :  std_logic;
signal bh7_w28_6_c1 :  std_logic;
signal bh7_w29_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_copy902_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid903_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid903_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_7_c1 :  std_logic;
signal bh7_w30_6_c1 :  std_logic;
signal bh7_w31_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_copy904_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid905_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid905_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_7_c1 :  std_logic;
signal bh7_w32_6_c1 :  std_logic;
signal bh7_w33_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_copy906_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid907_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid907_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_7_c1 :  std_logic;
signal bh7_w34_7_c1 :  std_logic;
signal bh7_w35_8_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_copy908_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid909_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid909_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w35_9_c1 :  std_logic;
signal bh7_w36_9_c1 :  std_logic;
signal bh7_w37_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_copy910_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid911_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid911_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w38_9_c1 :  std_logic;
signal bh7_w39_7_c1 :  std_logic;
signal bh7_w40_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_copy912_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid913_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid913_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w40_10_c1 :  std_logic;
signal bh7_w41_7_c1 :  std_logic;
signal bh7_w42_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_copy914_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid915_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid915_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w42_10_c1 :  std_logic;
signal bh7_w43_7_c1 :  std_logic;
signal bh7_w44_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_copy916_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid917_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid917_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w44_10_c1 :  std_logic;
signal bh7_w45_7_c1 :  std_logic;
signal bh7_w46_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_copy918_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid919_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid919_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w46_10_c1 :  std_logic;
signal bh7_w47_7_c1 :  std_logic;
signal bh7_w48_10_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_copy920_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid921_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid921_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w48_11_c1 :  std_logic;
signal bh7_w49_9_c1 :  std_logic;
signal bh7_w50_12_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_copy922_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid923_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid923_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w50_13_c1 :  std_logic;
signal bh7_w51_15_c1 :  std_logic;
signal bh7_w52_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_copy924_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid925_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid925_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w52_18_c1 :  std_logic;
signal bh7_w53_19_c1 :  std_logic;
signal bh7_w54_21_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_copy926_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid927_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid927_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w54_22_c1 :  std_logic;
signal bh7_w55_22_c1 :  std_logic;
signal bh7_w56_21_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_copy928_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid929_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid929_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_22_c1 :  std_logic;
signal bh7_w57_25_c1 :  std_logic;
signal bh7_w58_25_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_copy930_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid931_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid931_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w58_26_c1 :  std_logic;
signal bh7_w59_23_c1 :  std_logic;
signal bh7_w60_24_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_copy932_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid933_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid933_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w60_25_c1 :  std_logic;
signal bh7_w61_25_c1 :  std_logic;
signal bh7_w62_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_copy934_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid935_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid935_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_23_c1 :  std_logic;
signal bh7_w63_25_c1 :  std_logic;
signal bh7_w64_26_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_copy936_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid937_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid937_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_27_c1 :  std_logic;
signal bh7_w65_20_c1 :  std_logic;
signal bh7_w66_24_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_copy938_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid939_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid939_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w66_25_c1 :  std_logic;
signal bh7_w67_22_c1 :  std_logic;
signal bh7_w68_23_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_copy940_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid941_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid941_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_24_c1 :  std_logic;
signal bh7_w69_21_c1 :  std_logic;
signal bh7_w70_23_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_copy942_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid943_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid943_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w71_21_c1 :  std_logic;
signal bh7_w72_25_c1 :  std_logic;
signal bh7_w73_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_copy944_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid945_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid945_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w73_20_c1 :  std_logic;
signal bh7_w74_26_c1 :  std_logic;
signal bh7_w75_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_copy946_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid947_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid947_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w75_19_c1 :  std_logic;
signal bh7_w76_24_c1 :  std_logic;
signal bh7_w77_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_copy948_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid949_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid949_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_24_c1 :  std_logic;
signal bh7_w79_18_c1 :  std_logic;
signal bh7_w80_24_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_copy950_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid951_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid951_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_25_c1 :  std_logic;
signal bh7_w81_18_c1 :  std_logic;
signal bh7_w82_24_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_copy952_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid953_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid953_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_25_c1 :  std_logic;
signal bh7_w83_17_c1 :  std_logic;
signal bh7_w84_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_copy954_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid955_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid955_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_21_c1 :  std_logic;
signal bh7_w87_19_c1 :  std_logic;
signal bh7_w88_21_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_copy956_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid957_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid957_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_22_c1 :  std_logic;
signal bh7_w89_17_c1 :  std_logic;
signal bh7_w90_21_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_copy958_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid959_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid959_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w90_22_c1 :  std_logic;
signal bh7_w91_18_c1 :  std_logic;
signal bh7_w92_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_copy960_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid961_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid961_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w92_20_c1 :  std_logic;
signal bh7_w93_20_c1 :  std_logic;
signal bh7_w94_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_copy962_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid963_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid963_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w94_19_c1 :  std_logic;
signal bh7_w95_18_c1 :  std_logic;
signal bh7_w96_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_copy964_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid965_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid965_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w97_18_c1 :  std_logic;
signal bh7_w98_18_c1 :  std_logic;
signal bh7_w99_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_copy966_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid967_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid967_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w100_16_c1 :  std_logic;
signal bh7_w101_13_c1 :  std_logic;
signal bh7_w102_13_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_copy968_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid969_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid969_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w102_14_c1 :  std_logic;
signal bh7_w103_11_c1 :  std_logic;
signal bh7_w104_8_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_copy970_c1 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh7_22_c1, tmp_bitheapResult_bh7_22_c2 :  std_logic_vector(22 downto 0);
signal bitheapFinalAdd_bh7_In0_c1 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_In1_c1 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh7_Out_c2 :  std_logic_vector(83 downto 0);
signal bitheapResult_bh7_c2 :  std_logic_vector(105 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               bh7_w0_0_c1 <= bh7_w0_0_c0;
               bh7_w1_0_c1 <= bh7_w1_0_c0;
               bh7_w2_0_c1 <= bh7_w2_0_c0;
               bh7_w3_0_c1 <= bh7_w3_0_c0;
               bh7_w4_0_c1 <= bh7_w4_0_c0;
               bh7_w5_0_c1 <= bh7_w5_0_c0;
               bh7_w6_0_c1 <= bh7_w6_0_c0;
               bh7_w7_0_c1 <= bh7_w7_0_c0;
               bh7_w8_0_c1 <= bh7_w8_0_c0;
               bh7_w9_0_c1 <= bh7_w9_0_c0;
               bh7_w10_0_c1 <= bh7_w10_0_c0;
               bh7_w11_0_c1 <= bh7_w11_0_c0;
               bh7_w12_0_c1 <= bh7_w12_0_c0;
               bh7_w13_0_c1 <= bh7_w13_0_c0;
               bh7_w14_0_c1 <= bh7_w14_0_c0;
               bh7_w15_0_c1 <= bh7_w15_0_c0;
               bh7_w16_0_c1 <= bh7_w16_0_c0;
               bh7_w59_0_c1 <= bh7_w59_0_c0;
               bh7_w60_0_c1 <= bh7_w60_0_c0;
               bh7_w61_0_c1 <= bh7_w61_0_c0;
               bh7_w62_0_c1 <= bh7_w62_0_c0;
               bh7_w64_0_c1 <= bh7_w64_0_c0;
               bh7_w65_0_c1 <= bh7_w65_0_c0;
               bh7_w67_0_c1 <= bh7_w67_0_c0;
               bh7_w69_0_c1 <= bh7_w69_0_c0;
               bh7_w70_0_c1 <= bh7_w70_0_c0;
               bh7_w72_0_c1 <= bh7_w72_0_c0;
               bh7_w74_0_c1 <= bh7_w74_0_c0;
               bh7_w25_2_c1 <= bh7_w25_2_c0;
               bh7_w27_2_c1 <= bh7_w27_2_c0;
               bh7_w29_2_c1 <= bh7_w29_2_c0;
               bh7_w31_2_c1 <= bh7_w31_2_c0;
               bh7_w33_2_c1 <= bh7_w33_2_c0;
               bh7_w59_2_c1 <= bh7_w59_2_c0;
               bh7_w60_3_c1 <= bh7_w60_3_c0;
               bh7_w61_3_c1 <= bh7_w61_3_c0;
               bh7_w62_2_c1 <= bh7_w62_2_c0;
               bh7_w64_3_c1 <= bh7_w64_3_c0;
               bh7_w48_3_c1 <= bh7_w48_3_c0;
               bh7_w59_3_c1 <= bh7_w59_3_c0;
               bh7_w60_4_c1 <= bh7_w60_4_c0;
               bh7_w61_4_c1 <= bh7_w61_4_c0;
               bh7_w62_3_c1 <= bh7_w62_3_c0;
               bh7_w64_4_c1 <= bh7_w64_4_c0;
               bh7_w65_2_c1 <= bh7_w65_2_c0;
               bh7_w67_3_c1 <= bh7_w67_3_c0;
               bh7_w69_3_c1 <= bh7_w69_3_c0;
               bh7_w70_3_c1 <= bh7_w70_3_c0;
               bh7_w72_3_c1 <= bh7_w72_3_c0;
               bh7_w74_2_c1 <= bh7_w74_2_c0;
               bh7_w76_1_c1 <= bh7_w76_1_c0;
               bh7_w77_0_c1 <= bh7_w77_0_c0;
               bh7_w78_0_c1 <= bh7_w78_0_c0;
               bh7_w79_0_c1 <= bh7_w79_0_c0;
               bh7_w80_0_c1 <= bh7_w80_0_c0;
               bh7_w81_0_c1 <= bh7_w81_0_c0;
               bh7_w58_5_c1 <= bh7_w58_5_c0;
               bh7_w59_4_c1 <= bh7_w59_4_c0;
               bh7_w60_5_c1 <= bh7_w60_5_c0;
               bh7_w61_5_c1 <= bh7_w61_5_c0;
               bh7_w62_4_c1 <= bh7_w62_4_c0;
               bh7_w63_5_c1 <= bh7_w63_5_c0;
               bh7_w64_5_c1 <= bh7_w64_5_c0;
               bh7_w65_3_c1 <= bh7_w65_3_c0;
               bh7_w67_4_c1 <= bh7_w67_4_c0;
               bh7_w69_4_c1 <= bh7_w69_4_c0;
               bh7_w70_4_c1 <= bh7_w70_4_c0;
               bh7_w72_4_c1 <= bh7_w72_4_c0;
               bh7_w74_3_c1 <= bh7_w74_3_c0;
               bh7_w75_2_c1 <= bh7_w75_2_c0;
               bh7_w76_2_c1 <= bh7_w76_2_c0;
               bh7_w77_1_c1 <= bh7_w77_1_c0;
               bh7_w78_1_c1 <= bh7_w78_1_c0;
               bh7_w79_1_c1 <= bh7_w79_1_c0;
               bh7_w80_1_c1 <= bh7_w80_1_c0;
               bh7_w81_1_c1 <= bh7_w81_1_c0;
               bh7_w82_0_c1 <= bh7_w82_0_c0;
               bh7_w83_0_c1 <= bh7_w83_0_c0;
               bh7_w84_0_c1 <= bh7_w84_0_c0;
               bh7_w85_0_c1 <= bh7_w85_0_c0;
               bh7_w86_0_c1 <= bh7_w86_0_c0;
               bh7_w87_0_c1 <= bh7_w87_0_c0;
               bh7_w88_0_c1 <= bh7_w88_0_c0;
               bh7_w89_0_c1 <= bh7_w89_0_c0;
               bh7_w90_0_c1 <= bh7_w90_0_c0;
               bh7_w91_0_c1 <= bh7_w91_0_c0;
               bh7_w92_0_c1 <= bh7_w92_0_c0;
               bh7_w93_0_c1 <= bh7_w93_0_c0;
               bh7_w94_0_c1 <= bh7_w94_0_c0;
               bh7_w95_0_c1 <= bh7_w95_0_c0;
               bh7_w96_0_c1 <= bh7_w96_0_c0;
               bh7_w97_0_c1 <= bh7_w97_0_c0;
               bh7_w98_0_c1 <= bh7_w98_0_c0;
               bh7_w61_18_c1 <= bh7_w61_18_c0;
               bh7_w64_18_c1 <= bh7_w64_18_c0;
               bh7_w67_15_c1 <= bh7_w67_15_c0;
               bh7_w90_15_c1 <= bh7_w90_15_c0;
               bh7_w93_15_c1 <= bh7_w93_15_c0;
               bh7_w96_15_c1 <= bh7_w96_15_c0;
               bh7_w99_14_c1 <= bh7_w99_14_c0;
               bh7_w102_9_c1 <= bh7_w102_9_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c0;
            end if;
            if ce_2 = '1' then
               tmp_bitheapResult_bh7_22_c2 <= tmp_bitheapResult_bh7_22_c1;
            end if;
         end if;
      end process;
   XX_m6_c0 <= X ;
   YY_m6_c0 <= Y ;
   tile_0_X_c0 <= X(16 downto 0);
   tile_0_Y_c0 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid9
      port map ( clk  => clk,
                 X => tile_0_X_c0,
                 Y => tile_0_Y_c0,
                 R => tile_0_output_c0);

   tile_0_filtered_output_c0 <= unsigned(tile_0_output_c0(40 downto 0));
   bh7_w0_0_c0 <= tile_0_filtered_output_c0(0);
   bh7_w1_0_c0 <= tile_0_filtered_output_c0(1);
   bh7_w2_0_c0 <= tile_0_filtered_output_c0(2);
   bh7_w3_0_c0 <= tile_0_filtered_output_c0(3);
   bh7_w4_0_c0 <= tile_0_filtered_output_c0(4);
   bh7_w5_0_c0 <= tile_0_filtered_output_c0(5);
   bh7_w6_0_c0 <= tile_0_filtered_output_c0(6);
   bh7_w7_0_c0 <= tile_0_filtered_output_c0(7);
   bh7_w8_0_c0 <= tile_0_filtered_output_c0(8);
   bh7_w9_0_c0 <= tile_0_filtered_output_c0(9);
   bh7_w10_0_c0 <= tile_0_filtered_output_c0(10);
   bh7_w11_0_c0 <= tile_0_filtered_output_c0(11);
   bh7_w12_0_c0 <= tile_0_filtered_output_c0(12);
   bh7_w13_0_c0 <= tile_0_filtered_output_c0(13);
   bh7_w14_0_c0 <= tile_0_filtered_output_c0(14);
   bh7_w15_0_c0 <= tile_0_filtered_output_c0(15);
   bh7_w16_0_c0 <= tile_0_filtered_output_c0(16);
   bh7_w17_0_c0 <= tile_0_filtered_output_c0(17);
   bh7_w18_0_c0 <= tile_0_filtered_output_c0(18);
   bh7_w19_0_c0 <= tile_0_filtered_output_c0(19);
   bh7_w20_0_c0 <= tile_0_filtered_output_c0(20);
   bh7_w21_0_c0 <= tile_0_filtered_output_c0(21);
   bh7_w22_0_c0 <= tile_0_filtered_output_c0(22);
   bh7_w23_0_c0 <= tile_0_filtered_output_c0(23);
   bh7_w24_0_c0 <= tile_0_filtered_output_c0(24);
   bh7_w25_0_c0 <= tile_0_filtered_output_c0(25);
   bh7_w26_0_c0 <= tile_0_filtered_output_c0(26);
   bh7_w27_0_c0 <= tile_0_filtered_output_c0(27);
   bh7_w28_0_c0 <= tile_0_filtered_output_c0(28);
   bh7_w29_0_c0 <= tile_0_filtered_output_c0(29);
   bh7_w30_0_c0 <= tile_0_filtered_output_c0(30);
   bh7_w31_0_c0 <= tile_0_filtered_output_c0(31);
   bh7_w32_0_c0 <= tile_0_filtered_output_c0(32);
   bh7_w33_0_c0 <= tile_0_filtered_output_c0(33);
   bh7_w34_0_c0 <= tile_0_filtered_output_c0(34);
   bh7_w35_0_c0 <= tile_0_filtered_output_c0(35);
   bh7_w36_0_c0 <= tile_0_filtered_output_c0(36);
   bh7_w37_0_c0 <= tile_0_filtered_output_c0(37);
   bh7_w38_0_c0 <= tile_0_filtered_output_c0(38);
   bh7_w39_0_c0 <= tile_0_filtered_output_c0(39);
   bh7_w40_0_c0 <= tile_0_filtered_output_c0(40);
   tile_1_X_c0 <= X(33 downto 17);
   tile_1_Y_c0 <= Y(23 downto 0);
   tile_1_mult: DSPBlock_17x24_Freq300_uid11
      port map ( clk  => clk,
                 X => tile_1_X_c0,
                 Y => tile_1_Y_c0,
                 R => tile_1_output_c0);

   tile_1_filtered_output_c0 <= unsigned(tile_1_output_c0(40 downto 0));
   bh7_w17_1_c0 <= tile_1_filtered_output_c0(0);
   bh7_w18_1_c0 <= tile_1_filtered_output_c0(1);
   bh7_w19_1_c0 <= tile_1_filtered_output_c0(2);
   bh7_w20_1_c0 <= tile_1_filtered_output_c0(3);
   bh7_w21_1_c0 <= tile_1_filtered_output_c0(4);
   bh7_w22_1_c0 <= tile_1_filtered_output_c0(5);
   bh7_w23_1_c0 <= tile_1_filtered_output_c0(6);
   bh7_w24_1_c0 <= tile_1_filtered_output_c0(7);
   bh7_w25_1_c0 <= tile_1_filtered_output_c0(8);
   bh7_w26_1_c0 <= tile_1_filtered_output_c0(9);
   bh7_w27_1_c0 <= tile_1_filtered_output_c0(10);
   bh7_w28_1_c0 <= tile_1_filtered_output_c0(11);
   bh7_w29_1_c0 <= tile_1_filtered_output_c0(12);
   bh7_w30_1_c0 <= tile_1_filtered_output_c0(13);
   bh7_w31_1_c0 <= tile_1_filtered_output_c0(14);
   bh7_w32_1_c0 <= tile_1_filtered_output_c0(15);
   bh7_w33_1_c0 <= tile_1_filtered_output_c0(16);
   bh7_w34_1_c0 <= tile_1_filtered_output_c0(17);
   bh7_w35_1_c0 <= tile_1_filtered_output_c0(18);
   bh7_w36_1_c0 <= tile_1_filtered_output_c0(19);
   bh7_w37_1_c0 <= tile_1_filtered_output_c0(20);
   bh7_w38_1_c0 <= tile_1_filtered_output_c0(21);
   bh7_w39_1_c0 <= tile_1_filtered_output_c0(22);
   bh7_w40_1_c0 <= tile_1_filtered_output_c0(23);
   bh7_w41_0_c0 <= tile_1_filtered_output_c0(24);
   bh7_w42_0_c0 <= tile_1_filtered_output_c0(25);
   bh7_w43_0_c0 <= tile_1_filtered_output_c0(26);
   bh7_w44_0_c0 <= tile_1_filtered_output_c0(27);
   bh7_w45_0_c0 <= tile_1_filtered_output_c0(28);
   bh7_w46_0_c0 <= tile_1_filtered_output_c0(29);
   bh7_w47_0_c0 <= tile_1_filtered_output_c0(30);
   bh7_w48_0_c0 <= tile_1_filtered_output_c0(31);
   bh7_w49_0_c0 <= tile_1_filtered_output_c0(32);
   bh7_w50_0_c0 <= tile_1_filtered_output_c0(33);
   bh7_w51_0_c0 <= tile_1_filtered_output_c0(34);
   bh7_w52_0_c0 <= tile_1_filtered_output_c0(35);
   bh7_w53_0_c0 <= tile_1_filtered_output_c0(36);
   bh7_w54_0_c0 <= tile_1_filtered_output_c0(37);
   bh7_w55_0_c0 <= tile_1_filtered_output_c0(38);
   bh7_w56_0_c0 <= tile_1_filtered_output_c0(39);
   bh7_w57_0_c0 <= tile_1_filtered_output_c0(40);
   tile_2_X_c0 <= X(50 downto 34);
   tile_2_Y_c0 <= Y(23 downto 0);
   tile_2_mult: DSPBlock_17x24_Freq300_uid13
      port map ( clk  => clk,
                 X => tile_2_X_c0,
                 Y => tile_2_Y_c0,
                 R => tile_2_output_c0);

   tile_2_filtered_output_c0 <= unsigned(tile_2_output_c0(40 downto 0));
   bh7_w34_2_c0 <= tile_2_filtered_output_c0(0);
   bh7_w35_2_c0 <= tile_2_filtered_output_c0(1);
   bh7_w36_2_c0 <= tile_2_filtered_output_c0(2);
   bh7_w37_2_c0 <= tile_2_filtered_output_c0(3);
   bh7_w38_2_c0 <= tile_2_filtered_output_c0(4);
   bh7_w39_2_c0 <= tile_2_filtered_output_c0(5);
   bh7_w40_2_c0 <= tile_2_filtered_output_c0(6);
   bh7_w41_1_c0 <= tile_2_filtered_output_c0(7);
   bh7_w42_1_c0 <= tile_2_filtered_output_c0(8);
   bh7_w43_1_c0 <= tile_2_filtered_output_c0(9);
   bh7_w44_1_c0 <= tile_2_filtered_output_c0(10);
   bh7_w45_1_c0 <= tile_2_filtered_output_c0(11);
   bh7_w46_1_c0 <= tile_2_filtered_output_c0(12);
   bh7_w47_1_c0 <= tile_2_filtered_output_c0(13);
   bh7_w48_1_c0 <= tile_2_filtered_output_c0(14);
   bh7_w49_1_c0 <= tile_2_filtered_output_c0(15);
   bh7_w50_1_c0 <= tile_2_filtered_output_c0(16);
   bh7_w51_1_c0 <= tile_2_filtered_output_c0(17);
   bh7_w52_1_c0 <= tile_2_filtered_output_c0(18);
   bh7_w53_1_c0 <= tile_2_filtered_output_c0(19);
   bh7_w54_1_c0 <= tile_2_filtered_output_c0(20);
   bh7_w55_1_c0 <= tile_2_filtered_output_c0(21);
   bh7_w56_1_c0 <= tile_2_filtered_output_c0(22);
   bh7_w57_1_c0 <= tile_2_filtered_output_c0(23);
   bh7_w58_0_c0 <= tile_2_filtered_output_c0(24);
   bh7_w59_0_c0 <= tile_2_filtered_output_c0(25);
   bh7_w60_0_c0 <= tile_2_filtered_output_c0(26);
   bh7_w61_0_c0 <= tile_2_filtered_output_c0(27);
   bh7_w62_0_c0 <= tile_2_filtered_output_c0(28);
   bh7_w63_0_c0 <= tile_2_filtered_output_c0(29);
   bh7_w64_0_c0 <= tile_2_filtered_output_c0(30);
   bh7_w65_0_c0 <= tile_2_filtered_output_c0(31);
   bh7_w66_0_c0 <= tile_2_filtered_output_c0(32);
   bh7_w67_0_c0 <= tile_2_filtered_output_c0(33);
   bh7_w68_0_c0 <= tile_2_filtered_output_c0(34);
   bh7_w69_0_c0 <= tile_2_filtered_output_c0(35);
   bh7_w70_0_c0 <= tile_2_filtered_output_c0(36);
   bh7_w71_0_c0 <= tile_2_filtered_output_c0(37);
   bh7_w72_0_c0 <= tile_2_filtered_output_c0(38);
   bh7_w73_0_c0 <= tile_2_filtered_output_c0(39);
   bh7_w74_0_c0 <= tile_2_filtered_output_c0(40);
   tile_3_X_c0 <= X(52 downto 51);
   tile_3_Y_c0 <= Y(23 downto 21);
   tile_3_mult: IntMultiplierLUT_2x3_Freq300_uid15
      port map ( clk  => clk,
                 X => tile_3_X_c0,
                 Y => tile_3_Y_c0,
                 R => tile_3_output_c0);

   tile_3_filtered_output_c0 <= unsigned(tile_3_output_c0(4 downto 0));
   bh7_w72_1_c0 <= tile_3_filtered_output_c0(0);
   bh7_w73_1_c0 <= tile_3_filtered_output_c0(1);
   bh7_w74_1_c0 <= tile_3_filtered_output_c0(2);
   bh7_w75_0_c0 <= tile_3_filtered_output_c0(3);
   bh7_w76_0_c0 <= tile_3_filtered_output_c0(4);
   tile_4_X_c0 <= X(52 downto 51);
   tile_4_Y_c0 <= Y(20 downto 18);
   tile_4_mult: IntMultiplierLUT_2x3_Freq300_uid20
      port map ( clk  => clk,
                 X => tile_4_X_c0,
                 Y => tile_4_Y_c0,
                 R => tile_4_output_c0);

   tile_4_filtered_output_c0 <= unsigned(tile_4_output_c0(4 downto 0));
   bh7_w69_1_c0 <= tile_4_filtered_output_c0(0);
   bh7_w70_1_c0 <= tile_4_filtered_output_c0(1);
   bh7_w71_1_c0 <= tile_4_filtered_output_c0(2);
   bh7_w72_2_c0 <= tile_4_filtered_output_c0(3);
   bh7_w73_2_c0 <= tile_4_filtered_output_c0(4);
   tile_5_X_c0 <= X(52 downto 51);
   tile_5_Y_c0 <= Y(17 downto 15);
   tile_5_mult: IntMultiplierLUT_2x3_Freq300_uid25
      port map ( clk  => clk,
                 X => tile_5_X_c0,
                 Y => tile_5_Y_c0,
                 R => tile_5_output_c0);

   tile_5_filtered_output_c0 <= unsigned(tile_5_output_c0(4 downto 0));
   bh7_w66_1_c0 <= tile_5_filtered_output_c0(0);
   bh7_w67_1_c0 <= tile_5_filtered_output_c0(1);
   bh7_w68_1_c0 <= tile_5_filtered_output_c0(2);
   bh7_w69_2_c0 <= tile_5_filtered_output_c0(3);
   bh7_w70_2_c0 <= tile_5_filtered_output_c0(4);
   tile_6_X_c0 <= X(52 downto 51);
   tile_6_Y_c0 <= Y(14 downto 12);
   tile_6_mult: IntMultiplierLUT_2x3_Freq300_uid30
      port map ( clk  => clk,
                 X => tile_6_X_c0,
                 Y => tile_6_Y_c0,
                 R => tile_6_output_c0);

   tile_6_filtered_output_c0 <= unsigned(tile_6_output_c0(4 downto 0));
   bh7_w63_1_c0 <= tile_6_filtered_output_c0(0);
   bh7_w64_1_c0 <= tile_6_filtered_output_c0(1);
   bh7_w65_1_c0 <= tile_6_filtered_output_c0(2);
   bh7_w66_2_c0 <= tile_6_filtered_output_c0(3);
   bh7_w67_2_c0 <= tile_6_filtered_output_c0(4);
   tile_7_X_c0 <= X(52 downto 51);
   tile_7_Y_c0 <= Y(11 downto 9);
   tile_7_mult: IntMultiplierLUT_2x3_Freq300_uid35
      port map ( clk  => clk,
                 X => tile_7_X_c0,
                 Y => tile_7_Y_c0,
                 R => tile_7_output_c0);

   tile_7_filtered_output_c0 <= unsigned(tile_7_output_c0(4 downto 0));
   bh7_w60_1_c0 <= tile_7_filtered_output_c0(0);
   bh7_w61_1_c0 <= tile_7_filtered_output_c0(1);
   bh7_w62_1_c0 <= tile_7_filtered_output_c0(2);
   bh7_w63_2_c0 <= tile_7_filtered_output_c0(3);
   bh7_w64_2_c0 <= tile_7_filtered_output_c0(4);
   tile_8_X_c0 <= X(52 downto 51);
   tile_8_Y_c0 <= Y(8 downto 6);
   tile_8_mult: IntMultiplierLUT_2x3_Freq300_uid40
      port map ( clk  => clk,
                 X => tile_8_X_c0,
                 Y => tile_8_Y_c0,
                 R => tile_8_output_c0);

   tile_8_filtered_output_c0 <= unsigned(tile_8_output_c0(4 downto 0));
   bh7_w57_2_c0 <= tile_8_filtered_output_c0(0);
   bh7_w58_1_c0 <= tile_8_filtered_output_c0(1);
   bh7_w59_1_c0 <= tile_8_filtered_output_c0(2);
   bh7_w60_2_c0 <= tile_8_filtered_output_c0(3);
   bh7_w61_2_c0 <= tile_8_filtered_output_c0(4);
   tile_9_X_c0 <= X(52 downto 51);
   tile_9_Y_c0 <= Y(5 downto 3);
   tile_9_mult: IntMultiplierLUT_2x3_Freq300_uid45
      port map ( clk  => clk,
                 X => tile_9_X_c0,
                 Y => tile_9_Y_c0,
                 R => tile_9_output_c0);

   tile_9_filtered_output_c0 <= unsigned(tile_9_output_c0(4 downto 0));
   bh7_w54_2_c0 <= tile_9_filtered_output_c0(0);
   bh7_w55_2_c0 <= tile_9_filtered_output_c0(1);
   bh7_w56_2_c0 <= tile_9_filtered_output_c0(2);
   bh7_w57_3_c0 <= tile_9_filtered_output_c0(3);
   bh7_w58_2_c0 <= tile_9_filtered_output_c0(4);
   tile_10_X_c0 <= X(52 downto 51);
   tile_10_Y_c0 <= Y(2 downto 0);
   tile_10_mult: IntMultiplierLUT_2x3_Freq300_uid50
      port map ( clk  => clk,
                 X => tile_10_X_c0,
                 Y => tile_10_Y_c0,
                 R => tile_10_output_c0);

   tile_10_filtered_output_c0 <= unsigned(tile_10_output_c0(4 downto 0));
   bh7_w51_2_c0 <= tile_10_filtered_output_c0(0);
   bh7_w52_2_c0 <= tile_10_filtered_output_c0(1);
   bh7_w53_2_c0 <= tile_10_filtered_output_c0(2);
   bh7_w54_3_c0 <= tile_10_filtered_output_c0(3);
   bh7_w55_3_c0 <= tile_10_filtered_output_c0(4);
   tile_11_X_c0 <= X(16 downto 0);
   tile_11_Y_c0 <= Y(47 downto 24);
   tile_11_mult: DSPBlock_17x24_Freq300_uid55
      port map ( clk  => clk,
                 X => tile_11_X_c0,
                 Y => tile_11_Y_c0,
                 R => tile_11_output_c0);

   tile_11_filtered_output_c0 <= unsigned(tile_11_output_c0(40 downto 0));
   bh7_w24_2_c0 <= tile_11_filtered_output_c0(0);
   bh7_w25_2_c0 <= tile_11_filtered_output_c0(1);
   bh7_w26_2_c0 <= tile_11_filtered_output_c0(2);
   bh7_w27_2_c0 <= tile_11_filtered_output_c0(3);
   bh7_w28_2_c0 <= tile_11_filtered_output_c0(4);
   bh7_w29_2_c0 <= tile_11_filtered_output_c0(5);
   bh7_w30_2_c0 <= tile_11_filtered_output_c0(6);
   bh7_w31_2_c0 <= tile_11_filtered_output_c0(7);
   bh7_w32_2_c0 <= tile_11_filtered_output_c0(8);
   bh7_w33_2_c0 <= tile_11_filtered_output_c0(9);
   bh7_w34_3_c0 <= tile_11_filtered_output_c0(10);
   bh7_w35_3_c0 <= tile_11_filtered_output_c0(11);
   bh7_w36_3_c0 <= tile_11_filtered_output_c0(12);
   bh7_w37_3_c0 <= tile_11_filtered_output_c0(13);
   bh7_w38_3_c0 <= tile_11_filtered_output_c0(14);
   bh7_w39_3_c0 <= tile_11_filtered_output_c0(15);
   bh7_w40_3_c0 <= tile_11_filtered_output_c0(16);
   bh7_w41_2_c0 <= tile_11_filtered_output_c0(17);
   bh7_w42_2_c0 <= tile_11_filtered_output_c0(18);
   bh7_w43_2_c0 <= tile_11_filtered_output_c0(19);
   bh7_w44_2_c0 <= tile_11_filtered_output_c0(20);
   bh7_w45_2_c0 <= tile_11_filtered_output_c0(21);
   bh7_w46_2_c0 <= tile_11_filtered_output_c0(22);
   bh7_w47_2_c0 <= tile_11_filtered_output_c0(23);
   bh7_w48_2_c0 <= tile_11_filtered_output_c0(24);
   bh7_w49_2_c0 <= tile_11_filtered_output_c0(25);
   bh7_w50_2_c0 <= tile_11_filtered_output_c0(26);
   bh7_w51_3_c0 <= tile_11_filtered_output_c0(27);
   bh7_w52_3_c0 <= tile_11_filtered_output_c0(28);
   bh7_w53_3_c0 <= tile_11_filtered_output_c0(29);
   bh7_w54_4_c0 <= tile_11_filtered_output_c0(30);
   bh7_w55_4_c0 <= tile_11_filtered_output_c0(31);
   bh7_w56_3_c0 <= tile_11_filtered_output_c0(32);
   bh7_w57_4_c0 <= tile_11_filtered_output_c0(33);
   bh7_w58_3_c0 <= tile_11_filtered_output_c0(34);
   bh7_w59_2_c0 <= tile_11_filtered_output_c0(35);
   bh7_w60_3_c0 <= tile_11_filtered_output_c0(36);
   bh7_w61_3_c0 <= tile_11_filtered_output_c0(37);
   bh7_w62_2_c0 <= tile_11_filtered_output_c0(38);
   bh7_w63_3_c0 <= tile_11_filtered_output_c0(39);
   bh7_w64_3_c0 <= tile_11_filtered_output_c0(40);
   tile_12_X_c0 <= X(33 downto 17);
   tile_12_Y_c0 <= Y(47 downto 24);
   tile_12_mult: DSPBlock_17x24_Freq300_uid57
      port map ( clk  => clk,
                 X => tile_12_X_c0,
                 Y => tile_12_Y_c0,
                 R => tile_12_output_c0);

   tile_12_filtered_output_c0 <= unsigned(tile_12_output_c0(40 downto 0));
   bh7_w41_3_c0 <= tile_12_filtered_output_c0(0);
   bh7_w42_3_c0 <= tile_12_filtered_output_c0(1);
   bh7_w43_3_c0 <= tile_12_filtered_output_c0(2);
   bh7_w44_3_c0 <= tile_12_filtered_output_c0(3);
   bh7_w45_3_c0 <= tile_12_filtered_output_c0(4);
   bh7_w46_3_c0 <= tile_12_filtered_output_c0(5);
   bh7_w47_3_c0 <= tile_12_filtered_output_c0(6);
   bh7_w48_3_c0 <= tile_12_filtered_output_c0(7);
   bh7_w49_3_c0 <= tile_12_filtered_output_c0(8);
   bh7_w50_3_c0 <= tile_12_filtered_output_c0(9);
   bh7_w51_4_c0 <= tile_12_filtered_output_c0(10);
   bh7_w52_4_c0 <= tile_12_filtered_output_c0(11);
   bh7_w53_4_c0 <= tile_12_filtered_output_c0(12);
   bh7_w54_5_c0 <= tile_12_filtered_output_c0(13);
   bh7_w55_5_c0 <= tile_12_filtered_output_c0(14);
   bh7_w56_4_c0 <= tile_12_filtered_output_c0(15);
   bh7_w57_5_c0 <= tile_12_filtered_output_c0(16);
   bh7_w58_4_c0 <= tile_12_filtered_output_c0(17);
   bh7_w59_3_c0 <= tile_12_filtered_output_c0(18);
   bh7_w60_4_c0 <= tile_12_filtered_output_c0(19);
   bh7_w61_4_c0 <= tile_12_filtered_output_c0(20);
   bh7_w62_3_c0 <= tile_12_filtered_output_c0(21);
   bh7_w63_4_c0 <= tile_12_filtered_output_c0(22);
   bh7_w64_4_c0 <= tile_12_filtered_output_c0(23);
   bh7_w65_2_c0 <= tile_12_filtered_output_c0(24);
   bh7_w66_3_c0 <= tile_12_filtered_output_c0(25);
   bh7_w67_3_c0 <= tile_12_filtered_output_c0(26);
   bh7_w68_2_c0 <= tile_12_filtered_output_c0(27);
   bh7_w69_3_c0 <= tile_12_filtered_output_c0(28);
   bh7_w70_3_c0 <= tile_12_filtered_output_c0(29);
   bh7_w71_2_c0 <= tile_12_filtered_output_c0(30);
   bh7_w72_3_c0 <= tile_12_filtered_output_c0(31);
   bh7_w73_3_c0 <= tile_12_filtered_output_c0(32);
   bh7_w74_2_c0 <= tile_12_filtered_output_c0(33);
   bh7_w75_1_c0 <= tile_12_filtered_output_c0(34);
   bh7_w76_1_c0 <= tile_12_filtered_output_c0(35);
   bh7_w77_0_c0 <= tile_12_filtered_output_c0(36);
   bh7_w78_0_c0 <= tile_12_filtered_output_c0(37);
   bh7_w79_0_c0 <= tile_12_filtered_output_c0(38);
   bh7_w80_0_c0 <= tile_12_filtered_output_c0(39);
   bh7_w81_0_c0 <= tile_12_filtered_output_c0(40);
   tile_13_X_c0 <= X(50 downto 34);
   tile_13_Y_c0 <= Y(47 downto 24);
   tile_13_mult: DSPBlock_17x24_Freq300_uid59
      port map ( clk  => clk,
                 X => tile_13_X_c0,
                 Y => tile_13_Y_c0,
                 R => tile_13_output_c0);

   tile_13_filtered_output_c0 <= unsigned(tile_13_output_c0(40 downto 0));
   bh7_w58_5_c0 <= tile_13_filtered_output_c0(0);
   bh7_w59_4_c0 <= tile_13_filtered_output_c0(1);
   bh7_w60_5_c0 <= tile_13_filtered_output_c0(2);
   bh7_w61_5_c0 <= tile_13_filtered_output_c0(3);
   bh7_w62_4_c0 <= tile_13_filtered_output_c0(4);
   bh7_w63_5_c0 <= tile_13_filtered_output_c0(5);
   bh7_w64_5_c0 <= tile_13_filtered_output_c0(6);
   bh7_w65_3_c0 <= tile_13_filtered_output_c0(7);
   bh7_w66_4_c0 <= tile_13_filtered_output_c0(8);
   bh7_w67_4_c0 <= tile_13_filtered_output_c0(9);
   bh7_w68_3_c0 <= tile_13_filtered_output_c0(10);
   bh7_w69_4_c0 <= tile_13_filtered_output_c0(11);
   bh7_w70_4_c0 <= tile_13_filtered_output_c0(12);
   bh7_w71_3_c0 <= tile_13_filtered_output_c0(13);
   bh7_w72_4_c0 <= tile_13_filtered_output_c0(14);
   bh7_w73_4_c0 <= tile_13_filtered_output_c0(15);
   bh7_w74_3_c0 <= tile_13_filtered_output_c0(16);
   bh7_w75_2_c0 <= tile_13_filtered_output_c0(17);
   bh7_w76_2_c0 <= tile_13_filtered_output_c0(18);
   bh7_w77_1_c0 <= tile_13_filtered_output_c0(19);
   bh7_w78_1_c0 <= tile_13_filtered_output_c0(20);
   bh7_w79_1_c0 <= tile_13_filtered_output_c0(21);
   bh7_w80_1_c0 <= tile_13_filtered_output_c0(22);
   bh7_w81_1_c0 <= tile_13_filtered_output_c0(23);
   bh7_w82_0_c0 <= tile_13_filtered_output_c0(24);
   bh7_w83_0_c0 <= tile_13_filtered_output_c0(25);
   bh7_w84_0_c0 <= tile_13_filtered_output_c0(26);
   bh7_w85_0_c0 <= tile_13_filtered_output_c0(27);
   bh7_w86_0_c0 <= tile_13_filtered_output_c0(28);
   bh7_w87_0_c0 <= tile_13_filtered_output_c0(29);
   bh7_w88_0_c0 <= tile_13_filtered_output_c0(30);
   bh7_w89_0_c0 <= tile_13_filtered_output_c0(31);
   bh7_w90_0_c0 <= tile_13_filtered_output_c0(32);
   bh7_w91_0_c0 <= tile_13_filtered_output_c0(33);
   bh7_w92_0_c0 <= tile_13_filtered_output_c0(34);
   bh7_w93_0_c0 <= tile_13_filtered_output_c0(35);
   bh7_w94_0_c0 <= tile_13_filtered_output_c0(36);
   bh7_w95_0_c0 <= tile_13_filtered_output_c0(37);
   bh7_w96_0_c0 <= tile_13_filtered_output_c0(38);
   bh7_w97_0_c0 <= tile_13_filtered_output_c0(39);
   bh7_w98_0_c0 <= tile_13_filtered_output_c0(40);
   tile_14_X_c0 <= X(52 downto 51);
   tile_14_Y_c0 <= Y(47 downto 45);
   tile_14_mult: IntMultiplierLUT_2x3_Freq300_uid61
      port map ( clk  => clk,
                 X => tile_14_X_c0,
                 Y => tile_14_Y_c0,
                 R => tile_14_output_c0);

   tile_14_filtered_output_c0 <= unsigned(tile_14_output_c0(4 downto 0));
   bh7_w96_1_c0 <= tile_14_filtered_output_c0(0);
   bh7_w97_1_c0 <= tile_14_filtered_output_c0(1);
   bh7_w98_1_c0 <= tile_14_filtered_output_c0(2);
   bh7_w99_0_c0 <= tile_14_filtered_output_c0(3);
   bh7_w100_0_c0 <= tile_14_filtered_output_c0(4);
   tile_15_X_c0 <= X(52 downto 51);
   tile_15_Y_c0 <= Y(44 downto 42);
   tile_15_mult: IntMultiplierLUT_2x3_Freq300_uid66
      port map ( clk  => clk,
                 X => tile_15_X_c0,
                 Y => tile_15_Y_c0,
                 R => tile_15_output_c0);

   tile_15_filtered_output_c0 <= unsigned(tile_15_output_c0(4 downto 0));
   bh7_w93_1_c0 <= tile_15_filtered_output_c0(0);
   bh7_w94_1_c0 <= tile_15_filtered_output_c0(1);
   bh7_w95_1_c0 <= tile_15_filtered_output_c0(2);
   bh7_w96_2_c0 <= tile_15_filtered_output_c0(3);
   bh7_w97_2_c0 <= tile_15_filtered_output_c0(4);
   tile_16_X_c0 <= X(52 downto 51);
   tile_16_Y_c0 <= Y(41 downto 39);
   tile_16_mult: IntMultiplierLUT_2x3_Freq300_uid71
      port map ( clk  => clk,
                 X => tile_16_X_c0,
                 Y => tile_16_Y_c0,
                 R => tile_16_output_c0);

   tile_16_filtered_output_c0 <= unsigned(tile_16_output_c0(4 downto 0));
   bh7_w90_1_c0 <= tile_16_filtered_output_c0(0);
   bh7_w91_1_c0 <= tile_16_filtered_output_c0(1);
   bh7_w92_1_c0 <= tile_16_filtered_output_c0(2);
   bh7_w93_2_c0 <= tile_16_filtered_output_c0(3);
   bh7_w94_2_c0 <= tile_16_filtered_output_c0(4);
   tile_17_X_c0 <= X(52 downto 51);
   tile_17_Y_c0 <= Y(38 downto 36);
   tile_17_mult: IntMultiplierLUT_2x3_Freq300_uid76
      port map ( clk  => clk,
                 X => tile_17_X_c0,
                 Y => tile_17_Y_c0,
                 R => tile_17_output_c0);

   tile_17_filtered_output_c0 <= unsigned(tile_17_output_c0(4 downto 0));
   bh7_w87_1_c0 <= tile_17_filtered_output_c0(0);
   bh7_w88_1_c0 <= tile_17_filtered_output_c0(1);
   bh7_w89_1_c0 <= tile_17_filtered_output_c0(2);
   bh7_w90_2_c0 <= tile_17_filtered_output_c0(3);
   bh7_w91_2_c0 <= tile_17_filtered_output_c0(4);
   tile_18_X_c0 <= X(52 downto 51);
   tile_18_Y_c0 <= Y(35 downto 33);
   tile_18_mult: IntMultiplierLUT_2x3_Freq300_uid81
      port map ( clk  => clk,
                 X => tile_18_X_c0,
                 Y => tile_18_Y_c0,
                 R => tile_18_output_c0);

   tile_18_filtered_output_c0 <= unsigned(tile_18_output_c0(4 downto 0));
   bh7_w84_1_c0 <= tile_18_filtered_output_c0(0);
   bh7_w85_1_c0 <= tile_18_filtered_output_c0(1);
   bh7_w86_1_c0 <= tile_18_filtered_output_c0(2);
   bh7_w87_2_c0 <= tile_18_filtered_output_c0(3);
   bh7_w88_2_c0 <= tile_18_filtered_output_c0(4);
   tile_19_X_c0 <= X(52 downto 51);
   tile_19_Y_c0 <= Y(32 downto 30);
   tile_19_mult: IntMultiplierLUT_2x3_Freq300_uid86
      port map ( clk  => clk,
                 X => tile_19_X_c0,
                 Y => tile_19_Y_c0,
                 R => tile_19_output_c0);

   tile_19_filtered_output_c0 <= unsigned(tile_19_output_c0(4 downto 0));
   bh7_w81_2_c0 <= tile_19_filtered_output_c0(0);
   bh7_w82_1_c0 <= tile_19_filtered_output_c0(1);
   bh7_w83_1_c0 <= tile_19_filtered_output_c0(2);
   bh7_w84_2_c0 <= tile_19_filtered_output_c0(3);
   bh7_w85_2_c0 <= tile_19_filtered_output_c0(4);
   tile_20_X_c0 <= X(52 downto 51);
   tile_20_Y_c0 <= Y(29 downto 27);
   tile_20_mult: IntMultiplierLUT_2x3_Freq300_uid91
      port map ( clk  => clk,
                 X => tile_20_X_c0,
                 Y => tile_20_Y_c0,
                 R => tile_20_output_c0);

   tile_20_filtered_output_c0 <= unsigned(tile_20_output_c0(4 downto 0));
   bh7_w78_2_c0 <= tile_20_filtered_output_c0(0);
   bh7_w79_2_c0 <= tile_20_filtered_output_c0(1);
   bh7_w80_2_c0 <= tile_20_filtered_output_c0(2);
   bh7_w81_3_c0 <= tile_20_filtered_output_c0(3);
   bh7_w82_2_c0 <= tile_20_filtered_output_c0(4);
   tile_21_X_c0 <= X(52 downto 51);
   tile_21_Y_c0 <= Y(26 downto 24);
   tile_21_mult: IntMultiplierLUT_2x3_Freq300_uid96
      port map ( clk  => clk,
                 X => tile_21_X_c0,
                 Y => tile_21_Y_c0,
                 R => tile_21_output_c0);

   tile_21_filtered_output_c0 <= unsigned(tile_21_output_c0(4 downto 0));
   bh7_w75_3_c0 <= tile_21_filtered_output_c0(0);
   bh7_w76_3_c0 <= tile_21_filtered_output_c0(1);
   bh7_w77_2_c0 <= tile_21_filtered_output_c0(2);
   bh7_w78_3_c0 <= tile_21_filtered_output_c0(3);
   bh7_w79_3_c0 <= tile_21_filtered_output_c0(4);
   tile_22_X_c0 <= X(16 downto 16);
   tile_22_Y_c0 <= Y(52 downto 52);
   tile_22_mult: IntMultiplierLUT_1x1_Freq300_uid101
      port map ( clk  => clk,
                 X => tile_22_X_c0,
                 Y => tile_22_Y_c0,
                 R => tile_22_output_c0);

   tile_22_filtered_output_c0 <= unsigned(tile_22_output_c0(0 downto 0));
   bh7_w68_4_c0 <= tile_22_filtered_output_c0(0);
   tile_23_X_c0 <= X(15 downto 12);
   tile_23_Y_c0 <= Y(52 downto 52);
   tile_23_mult: IntMultiplierLUT_4x1_Freq300_uid103
      port map ( clk  => clk,
                 X => tile_23_X_c0,
                 Y => tile_23_Y_c0,
                 R => tile_23_output_c0);

   tile_23_filtered_output_c0 <= unsigned(tile_23_output_c0(3 downto 0));
   bh7_w64_6_c0 <= tile_23_filtered_output_c0(0);
   bh7_w65_4_c0 <= tile_23_filtered_output_c0(1);
   bh7_w66_5_c0 <= tile_23_filtered_output_c0(2);
   bh7_w67_5_c0 <= tile_23_filtered_output_c0(3);
   tile_24_X_c0 <= X(11 downto 8);
   tile_24_Y_c0 <= Y(52 downto 52);
   tile_24_mult: IntMultiplierLUT_4x1_Freq300_uid105
      port map ( clk  => clk,
                 X => tile_24_X_c0,
                 Y => tile_24_Y_c0,
                 R => tile_24_output_c0);

   tile_24_filtered_output_c0 <= unsigned(tile_24_output_c0(3 downto 0));
   bh7_w60_6_c0 <= tile_24_filtered_output_c0(0);
   bh7_w61_6_c0 <= tile_24_filtered_output_c0(1);
   bh7_w62_5_c0 <= tile_24_filtered_output_c0(2);
   bh7_w63_6_c0 <= tile_24_filtered_output_c0(3);
   tile_25_X_c0 <= X(7 downto 4);
   tile_25_Y_c0 <= Y(52 downto 52);
   tile_25_mult: IntMultiplierLUT_4x1_Freq300_uid107
      port map ( clk  => clk,
                 X => tile_25_X_c0,
                 Y => tile_25_Y_c0,
                 R => tile_25_output_c0);

   tile_25_filtered_output_c0 <= unsigned(tile_25_output_c0(3 downto 0));
   bh7_w56_5_c0 <= tile_25_filtered_output_c0(0);
   bh7_w57_6_c0 <= tile_25_filtered_output_c0(1);
   bh7_w58_6_c0 <= tile_25_filtered_output_c0(2);
   bh7_w59_5_c0 <= tile_25_filtered_output_c0(3);
   tile_26_X_c0 <= X(3 downto 0);
   tile_26_Y_c0 <= Y(52 downto 52);
   tile_26_mult: IntMultiplierLUT_4x1_Freq300_uid109
      port map ( clk  => clk,
                 X => tile_26_X_c0,
                 Y => tile_26_Y_c0,
                 R => tile_26_output_c0);

   tile_26_filtered_output_c0 <= unsigned(tile_26_output_c0(3 downto 0));
   bh7_w52_5_c0 <= tile_26_filtered_output_c0(0);
   bh7_w53_5_c0 <= tile_26_filtered_output_c0(1);
   bh7_w54_6_c0 <= tile_26_filtered_output_c0(2);
   bh7_w55_6_c0 <= tile_26_filtered_output_c0(3);
   tile_27_X_c0 <= X(16 downto 15);
   tile_27_Y_c0 <= Y(51 downto 50);
   tile_27_mult: IntMultiplierLUT_2x2_Freq300_uid111
      port map ( clk  => clk,
                 X => tile_27_X_c0,
                 Y => tile_27_Y_c0,
                 R => tile_27_output_c0);

   tile_27_filtered_output_c0 <= unsigned(tile_27_output_c0(3 downto 0));
   bh7_w65_5_c0 <= tile_27_filtered_output_c0(0);
   bh7_w66_6_c0 <= tile_27_filtered_output_c0(1);
   bh7_w67_6_c0 <= tile_27_filtered_output_c0(2);
   bh7_w68_5_c0 <= tile_27_filtered_output_c0(3);
   tile_28_X_c0 <= X(14 downto 12);
   tile_28_Y_c0 <= Y(51 downto 50);
   tile_28_mult: IntMultiplierLUT_3x2_Freq300_uid116
      port map ( clk  => clk,
                 X => tile_28_X_c0,
                 Y => tile_28_Y_c0,
                 R => tile_28_output_c0);

   tile_28_filtered_output_c0 <= unsigned(tile_28_output_c0(4 downto 0));
   bh7_w62_6_c0 <= tile_28_filtered_output_c0(0);
   bh7_w63_7_c0 <= tile_28_filtered_output_c0(1);
   bh7_w64_7_c0 <= tile_28_filtered_output_c0(2);
   bh7_w65_6_c0 <= tile_28_filtered_output_c0(3);
   bh7_w66_7_c0 <= tile_28_filtered_output_c0(4);
   tile_29_X_c0 <= X(11 downto 9);
   tile_29_Y_c0 <= Y(51 downto 50);
   tile_29_mult: IntMultiplierLUT_3x2_Freq300_uid121
      port map ( clk  => clk,
                 X => tile_29_X_c0,
                 Y => tile_29_Y_c0,
                 R => tile_29_output_c0);

   tile_29_filtered_output_c0 <= unsigned(tile_29_output_c0(4 downto 0));
   bh7_w59_6_c0 <= tile_29_filtered_output_c0(0);
   bh7_w60_7_c0 <= tile_29_filtered_output_c0(1);
   bh7_w61_7_c0 <= tile_29_filtered_output_c0(2);
   bh7_w62_7_c0 <= tile_29_filtered_output_c0(3);
   bh7_w63_8_c0 <= tile_29_filtered_output_c0(4);
   tile_30_X_c0 <= X(8 downto 6);
   tile_30_Y_c0 <= Y(51 downto 50);
   tile_30_mult: IntMultiplierLUT_3x2_Freq300_uid126
      port map ( clk  => clk,
                 X => tile_30_X_c0,
                 Y => tile_30_Y_c0,
                 R => tile_30_output_c0);

   tile_30_filtered_output_c0 <= unsigned(tile_30_output_c0(4 downto 0));
   bh7_w56_6_c0 <= tile_30_filtered_output_c0(0);
   bh7_w57_7_c0 <= tile_30_filtered_output_c0(1);
   bh7_w58_7_c0 <= tile_30_filtered_output_c0(2);
   bh7_w59_7_c0 <= tile_30_filtered_output_c0(3);
   bh7_w60_8_c0 <= tile_30_filtered_output_c0(4);
   tile_31_X_c0 <= X(5 downto 3);
   tile_31_Y_c0 <= Y(51 downto 50);
   tile_31_mult: IntMultiplierLUT_3x2_Freq300_uid131
      port map ( clk  => clk,
                 X => tile_31_X_c0,
                 Y => tile_31_Y_c0,
                 R => tile_31_output_c0);

   tile_31_filtered_output_c0 <= unsigned(tile_31_output_c0(4 downto 0));
   bh7_w53_6_c0 <= tile_31_filtered_output_c0(0);
   bh7_w54_7_c0 <= tile_31_filtered_output_c0(1);
   bh7_w55_7_c0 <= tile_31_filtered_output_c0(2);
   bh7_w56_7_c0 <= tile_31_filtered_output_c0(3);
   bh7_w57_8_c0 <= tile_31_filtered_output_c0(4);
   tile_32_X_c0 <= X(2 downto 0);
   tile_32_Y_c0 <= Y(51 downto 50);
   tile_32_mult: IntMultiplierLUT_3x2_Freq300_uid136
      port map ( clk  => clk,
                 X => tile_32_X_c0,
                 Y => tile_32_Y_c0,
                 R => tile_32_output_c0);

   tile_32_filtered_output_c0 <= unsigned(tile_32_output_c0(4 downto 0));
   bh7_w50_4_c0 <= tile_32_filtered_output_c0(0);
   bh7_w51_5_c0 <= tile_32_filtered_output_c0(1);
   bh7_w52_6_c0 <= tile_32_filtered_output_c0(2);
   bh7_w53_7_c0 <= tile_32_filtered_output_c0(3);
   bh7_w54_8_c0 <= tile_32_filtered_output_c0(4);
   tile_33_X_c0 <= X(16 downto 15);
   tile_33_Y_c0 <= Y(49 downto 48);
   tile_33_mult: IntMultiplierLUT_2x2_Freq300_uid141
      port map ( clk  => clk,
                 X => tile_33_X_c0,
                 Y => tile_33_Y_c0,
                 R => tile_33_output_c0);

   tile_33_filtered_output_c0 <= unsigned(tile_33_output_c0(3 downto 0));
   bh7_w63_9_c0 <= tile_33_filtered_output_c0(0);
   bh7_w64_8_c0 <= tile_33_filtered_output_c0(1);
   bh7_w65_7_c0 <= tile_33_filtered_output_c0(2);
   bh7_w66_8_c0 <= tile_33_filtered_output_c0(3);
   tile_34_X_c0 <= X(14 downto 12);
   tile_34_Y_c0 <= Y(49 downto 48);
   tile_34_mult: IntMultiplierLUT_3x2_Freq300_uid146
      port map ( clk  => clk,
                 X => tile_34_X_c0,
                 Y => tile_34_Y_c0,
                 R => tile_34_output_c0);

   tile_34_filtered_output_c0 <= unsigned(tile_34_output_c0(4 downto 0));
   bh7_w60_9_c0 <= tile_34_filtered_output_c0(0);
   bh7_w61_8_c0 <= tile_34_filtered_output_c0(1);
   bh7_w62_8_c0 <= tile_34_filtered_output_c0(2);
   bh7_w63_10_c0 <= tile_34_filtered_output_c0(3);
   bh7_w64_9_c0 <= tile_34_filtered_output_c0(4);
   tile_35_X_c0 <= X(11 downto 9);
   tile_35_Y_c0 <= Y(49 downto 48);
   tile_35_mult: IntMultiplierLUT_3x2_Freq300_uid151
      port map ( clk  => clk,
                 X => tile_35_X_c0,
                 Y => tile_35_Y_c0,
                 R => tile_35_output_c0);

   tile_35_filtered_output_c0 <= unsigned(tile_35_output_c0(4 downto 0));
   bh7_w57_9_c0 <= tile_35_filtered_output_c0(0);
   bh7_w58_8_c0 <= tile_35_filtered_output_c0(1);
   bh7_w59_8_c0 <= tile_35_filtered_output_c0(2);
   bh7_w60_10_c0 <= tile_35_filtered_output_c0(3);
   bh7_w61_9_c0 <= tile_35_filtered_output_c0(4);
   tile_36_X_c0 <= X(8 downto 6);
   tile_36_Y_c0 <= Y(49 downto 48);
   tile_36_mult: IntMultiplierLUT_3x2_Freq300_uid156
      port map ( clk  => clk,
                 X => tile_36_X_c0,
                 Y => tile_36_Y_c0,
                 R => tile_36_output_c0);

   tile_36_filtered_output_c0 <= unsigned(tile_36_output_c0(4 downto 0));
   bh7_w54_9_c0 <= tile_36_filtered_output_c0(0);
   bh7_w55_8_c0 <= tile_36_filtered_output_c0(1);
   bh7_w56_8_c0 <= tile_36_filtered_output_c0(2);
   bh7_w57_10_c0 <= tile_36_filtered_output_c0(3);
   bh7_w58_9_c0 <= tile_36_filtered_output_c0(4);
   tile_37_X_c0 <= X(5 downto 3);
   tile_37_Y_c0 <= Y(49 downto 48);
   tile_37_mult: IntMultiplierLUT_3x2_Freq300_uid161
      port map ( clk  => clk,
                 X => tile_37_X_c0,
                 Y => tile_37_Y_c0,
                 R => tile_37_output_c0);

   tile_37_filtered_output_c0 <= unsigned(tile_37_output_c0(4 downto 0));
   bh7_w51_6_c0 <= tile_37_filtered_output_c0(0);
   bh7_w52_7_c0 <= tile_37_filtered_output_c0(1);
   bh7_w53_8_c0 <= tile_37_filtered_output_c0(2);
   bh7_w54_10_c0 <= tile_37_filtered_output_c0(3);
   bh7_w55_9_c0 <= tile_37_filtered_output_c0(4);
   tile_38_X_c0 <= X(2 downto 0);
   tile_38_Y_c0 <= Y(49 downto 48);
   tile_38_mult: IntMultiplierLUT_3x2_Freq300_uid166
      port map ( clk  => clk,
                 X => tile_38_X_c0,
                 Y => tile_38_Y_c0,
                 R => tile_38_output_c0);

   tile_38_filtered_output_c0 <= unsigned(tile_38_output_c0(4 downto 0));
   bh7_w48_4_c0 <= tile_38_filtered_output_c0(0);
   bh7_w49_4_c0 <= tile_38_filtered_output_c0(1);
   bh7_w50_5_c0 <= tile_38_filtered_output_c0(2);
   bh7_w51_7_c0 <= tile_38_filtered_output_c0(3);
   bh7_w52_8_c0 <= tile_38_filtered_output_c0(4);
   tile_39_X_c0 <= X(33 downto 33);
   tile_39_Y_c0 <= Y(52 downto 52);
   tile_39_mult: IntMultiplierLUT_1x1_Freq300_uid171
      port map ( clk  => clk,
                 X => tile_39_X_c0,
                 Y => tile_39_Y_c0,
                 R => tile_39_output_c0);

   tile_39_filtered_output_c0 <= unsigned(tile_39_output_c0(0 downto 0));
   bh7_w85_3_c0 <= tile_39_filtered_output_c0(0);
   tile_40_X_c0 <= X(32 downto 29);
   tile_40_Y_c0 <= Y(52 downto 52);
   tile_40_mult: IntMultiplierLUT_4x1_Freq300_uid173
      port map ( clk  => clk,
                 X => tile_40_X_c0,
                 Y => tile_40_Y_c0,
                 R => tile_40_output_c0);

   tile_40_filtered_output_c0 <= unsigned(tile_40_output_c0(3 downto 0));
   bh7_w81_4_c0 <= tile_40_filtered_output_c0(0);
   bh7_w82_3_c0 <= tile_40_filtered_output_c0(1);
   bh7_w83_2_c0 <= tile_40_filtered_output_c0(2);
   bh7_w84_3_c0 <= tile_40_filtered_output_c0(3);
   tile_41_X_c0 <= X(28 downto 25);
   tile_41_Y_c0 <= Y(52 downto 52);
   tile_41_mult: IntMultiplierLUT_4x1_Freq300_uid175
      port map ( clk  => clk,
                 X => tile_41_X_c0,
                 Y => tile_41_Y_c0,
                 R => tile_41_output_c0);

   tile_41_filtered_output_c0 <= unsigned(tile_41_output_c0(3 downto 0));
   bh7_w77_3_c0 <= tile_41_filtered_output_c0(0);
   bh7_w78_4_c0 <= tile_41_filtered_output_c0(1);
   bh7_w79_4_c0 <= tile_41_filtered_output_c0(2);
   bh7_w80_3_c0 <= tile_41_filtered_output_c0(3);
   tile_42_X_c0 <= X(24 downto 21);
   tile_42_Y_c0 <= Y(52 downto 52);
   tile_42_mult: IntMultiplierLUT_4x1_Freq300_uid177
      port map ( clk  => clk,
                 X => tile_42_X_c0,
                 Y => tile_42_Y_c0,
                 R => tile_42_output_c0);

   tile_42_filtered_output_c0 <= unsigned(tile_42_output_c0(3 downto 0));
   bh7_w73_5_c0 <= tile_42_filtered_output_c0(0);
   bh7_w74_4_c0 <= tile_42_filtered_output_c0(1);
   bh7_w75_4_c0 <= tile_42_filtered_output_c0(2);
   bh7_w76_4_c0 <= tile_42_filtered_output_c0(3);
   tile_43_X_c0 <= X(20 downto 17);
   tile_43_Y_c0 <= Y(52 downto 52);
   tile_43_mult: IntMultiplierLUT_4x1_Freq300_uid179
      port map ( clk  => clk,
                 X => tile_43_X_c0,
                 Y => tile_43_Y_c0,
                 R => tile_43_output_c0);

   tile_43_filtered_output_c0 <= unsigned(tile_43_output_c0(3 downto 0));
   bh7_w69_5_c0 <= tile_43_filtered_output_c0(0);
   bh7_w70_5_c0 <= tile_43_filtered_output_c0(1);
   bh7_w71_4_c0 <= tile_43_filtered_output_c0(2);
   bh7_w72_5_c0 <= tile_43_filtered_output_c0(3);
   tile_44_X_c0 <= X(33 downto 32);
   tile_44_Y_c0 <= Y(51 downto 50);
   tile_44_mult: IntMultiplierLUT_2x2_Freq300_uid181
      port map ( clk  => clk,
                 X => tile_44_X_c0,
                 Y => tile_44_Y_c0,
                 R => tile_44_output_c0);

   tile_44_filtered_output_c0 <= unsigned(tile_44_output_c0(3 downto 0));
   bh7_w82_4_c0 <= tile_44_filtered_output_c0(0);
   bh7_w83_3_c0 <= tile_44_filtered_output_c0(1);
   bh7_w84_4_c0 <= tile_44_filtered_output_c0(2);
   bh7_w85_4_c0 <= tile_44_filtered_output_c0(3);
   tile_45_X_c0 <= X(31 downto 29);
   tile_45_Y_c0 <= Y(51 downto 50);
   tile_45_mult: IntMultiplierLUT_3x2_Freq300_uid186
      port map ( clk  => clk,
                 X => tile_45_X_c0,
                 Y => tile_45_Y_c0,
                 R => tile_45_output_c0);

   tile_45_filtered_output_c0 <= unsigned(tile_45_output_c0(4 downto 0));
   bh7_w79_5_c0 <= tile_45_filtered_output_c0(0);
   bh7_w80_4_c0 <= tile_45_filtered_output_c0(1);
   bh7_w81_5_c0 <= tile_45_filtered_output_c0(2);
   bh7_w82_5_c0 <= tile_45_filtered_output_c0(3);
   bh7_w83_4_c0 <= tile_45_filtered_output_c0(4);
   tile_46_X_c0 <= X(28 downto 26);
   tile_46_Y_c0 <= Y(51 downto 50);
   tile_46_mult: IntMultiplierLUT_3x2_Freq300_uid191
      port map ( clk  => clk,
                 X => tile_46_X_c0,
                 Y => tile_46_Y_c0,
                 R => tile_46_output_c0);

   tile_46_filtered_output_c0 <= unsigned(tile_46_output_c0(4 downto 0));
   bh7_w76_5_c0 <= tile_46_filtered_output_c0(0);
   bh7_w77_4_c0 <= tile_46_filtered_output_c0(1);
   bh7_w78_5_c0 <= tile_46_filtered_output_c0(2);
   bh7_w79_6_c0 <= tile_46_filtered_output_c0(3);
   bh7_w80_5_c0 <= tile_46_filtered_output_c0(4);
   tile_47_X_c0 <= X(25 downto 23);
   tile_47_Y_c0 <= Y(51 downto 50);
   tile_47_mult: IntMultiplierLUT_3x2_Freq300_uid196
      port map ( clk  => clk,
                 X => tile_47_X_c0,
                 Y => tile_47_Y_c0,
                 R => tile_47_output_c0);

   tile_47_filtered_output_c0 <= unsigned(tile_47_output_c0(4 downto 0));
   bh7_w73_6_c0 <= tile_47_filtered_output_c0(0);
   bh7_w74_5_c0 <= tile_47_filtered_output_c0(1);
   bh7_w75_5_c0 <= tile_47_filtered_output_c0(2);
   bh7_w76_6_c0 <= tile_47_filtered_output_c0(3);
   bh7_w77_5_c0 <= tile_47_filtered_output_c0(4);
   tile_48_X_c0 <= X(22 downto 20);
   tile_48_Y_c0 <= Y(51 downto 50);
   tile_48_mult: IntMultiplierLUT_3x2_Freq300_uid201
      port map ( clk  => clk,
                 X => tile_48_X_c0,
                 Y => tile_48_Y_c0,
                 R => tile_48_output_c0);

   tile_48_filtered_output_c0 <= unsigned(tile_48_output_c0(4 downto 0));
   bh7_w70_6_c0 <= tile_48_filtered_output_c0(0);
   bh7_w71_5_c0 <= tile_48_filtered_output_c0(1);
   bh7_w72_6_c0 <= tile_48_filtered_output_c0(2);
   bh7_w73_7_c0 <= tile_48_filtered_output_c0(3);
   bh7_w74_6_c0 <= tile_48_filtered_output_c0(4);
   tile_49_X_c0 <= X(19 downto 17);
   tile_49_Y_c0 <= Y(51 downto 50);
   tile_49_mult: IntMultiplierLUT_3x2_Freq300_uid206
      port map ( clk  => clk,
                 X => tile_49_X_c0,
                 Y => tile_49_Y_c0,
                 R => tile_49_output_c0);

   tile_49_filtered_output_c0 <= unsigned(tile_49_output_c0(4 downto 0));
   bh7_w67_7_c0 <= tile_49_filtered_output_c0(0);
   bh7_w68_6_c0 <= tile_49_filtered_output_c0(1);
   bh7_w69_6_c0 <= tile_49_filtered_output_c0(2);
   bh7_w70_7_c0 <= tile_49_filtered_output_c0(3);
   bh7_w71_6_c0 <= tile_49_filtered_output_c0(4);
   tile_50_X_c0 <= X(33 downto 32);
   tile_50_Y_c0 <= Y(49 downto 48);
   tile_50_mult: IntMultiplierLUT_2x2_Freq300_uid211
      port map ( clk  => clk,
                 X => tile_50_X_c0,
                 Y => tile_50_Y_c0,
                 R => tile_50_output_c0);

   tile_50_filtered_output_c0 <= unsigned(tile_50_output_c0(3 downto 0));
   bh7_w80_6_c0 <= tile_50_filtered_output_c0(0);
   bh7_w81_6_c0 <= tile_50_filtered_output_c0(1);
   bh7_w82_6_c0 <= tile_50_filtered_output_c0(2);
   bh7_w83_5_c0 <= tile_50_filtered_output_c0(3);
   tile_51_X_c0 <= X(31 downto 29);
   tile_51_Y_c0 <= Y(49 downto 48);
   tile_51_mult: IntMultiplierLUT_3x2_Freq300_uid216
      port map ( clk  => clk,
                 X => tile_51_X_c0,
                 Y => tile_51_Y_c0,
                 R => tile_51_output_c0);

   tile_51_filtered_output_c0 <= unsigned(tile_51_output_c0(4 downto 0));
   bh7_w77_6_c0 <= tile_51_filtered_output_c0(0);
   bh7_w78_6_c0 <= tile_51_filtered_output_c0(1);
   bh7_w79_7_c0 <= tile_51_filtered_output_c0(2);
   bh7_w80_7_c0 <= tile_51_filtered_output_c0(3);
   bh7_w81_7_c0 <= tile_51_filtered_output_c0(4);
   tile_52_X_c0 <= X(28 downto 26);
   tile_52_Y_c0 <= Y(49 downto 48);
   tile_52_mult: IntMultiplierLUT_3x2_Freq300_uid221
      port map ( clk  => clk,
                 X => tile_52_X_c0,
                 Y => tile_52_Y_c0,
                 R => tile_52_output_c0);

   tile_52_filtered_output_c0 <= unsigned(tile_52_output_c0(4 downto 0));
   bh7_w74_7_c0 <= tile_52_filtered_output_c0(0);
   bh7_w75_6_c0 <= tile_52_filtered_output_c0(1);
   bh7_w76_7_c0 <= tile_52_filtered_output_c0(2);
   bh7_w77_7_c0 <= tile_52_filtered_output_c0(3);
   bh7_w78_7_c0 <= tile_52_filtered_output_c0(4);
   tile_53_X_c0 <= X(25 downto 23);
   tile_53_Y_c0 <= Y(49 downto 48);
   tile_53_mult: IntMultiplierLUT_3x2_Freq300_uid226
      port map ( clk  => clk,
                 X => tile_53_X_c0,
                 Y => tile_53_Y_c0,
                 R => tile_53_output_c0);

   tile_53_filtered_output_c0 <= unsigned(tile_53_output_c0(4 downto 0));
   bh7_w71_7_c0 <= tile_53_filtered_output_c0(0);
   bh7_w72_7_c0 <= tile_53_filtered_output_c0(1);
   bh7_w73_8_c0 <= tile_53_filtered_output_c0(2);
   bh7_w74_8_c0 <= tile_53_filtered_output_c0(3);
   bh7_w75_7_c0 <= tile_53_filtered_output_c0(4);
   tile_54_X_c0 <= X(22 downto 20);
   tile_54_Y_c0 <= Y(49 downto 48);
   tile_54_mult: IntMultiplierLUT_3x2_Freq300_uid231
      port map ( clk  => clk,
                 X => tile_54_X_c0,
                 Y => tile_54_Y_c0,
                 R => tile_54_output_c0);

   tile_54_filtered_output_c0 <= unsigned(tile_54_output_c0(4 downto 0));
   bh7_w68_7_c0 <= tile_54_filtered_output_c0(0);
   bh7_w69_7_c0 <= tile_54_filtered_output_c0(1);
   bh7_w70_8_c0 <= tile_54_filtered_output_c0(2);
   bh7_w71_8_c0 <= tile_54_filtered_output_c0(3);
   bh7_w72_8_c0 <= tile_54_filtered_output_c0(4);
   tile_55_X_c0 <= X(19 downto 17);
   tile_55_Y_c0 <= Y(49 downto 48);
   tile_55_mult: IntMultiplierLUT_3x2_Freq300_uid236
      port map ( clk  => clk,
                 X => tile_55_X_c0,
                 Y => tile_55_Y_c0,
                 R => tile_55_output_c0);

   tile_55_filtered_output_c0 <= unsigned(tile_55_output_c0(4 downto 0));
   bh7_w65_8_c0 <= tile_55_filtered_output_c0(0);
   bh7_w66_9_c0 <= tile_55_filtered_output_c0(1);
   bh7_w67_8_c0 <= tile_55_filtered_output_c0(2);
   bh7_w68_8_c0 <= tile_55_filtered_output_c0(3);
   bh7_w69_8_c0 <= tile_55_filtered_output_c0(4);
   tile_56_X_c0 <= X(50 downto 50);
   tile_56_Y_c0 <= Y(52 downto 52);
   tile_56_mult: IntMultiplierLUT_1x1_Freq300_uid241
      port map ( clk  => clk,
                 X => tile_56_X_c0,
                 Y => tile_56_Y_c0,
                 R => tile_56_output_c0);

   tile_56_filtered_output_c0 <= unsigned(tile_56_output_c0(0 downto 0));
   bh7_w102_0_c0 <= tile_56_filtered_output_c0(0);
   tile_57_X_c0 <= X(49 downto 46);
   tile_57_Y_c0 <= Y(52 downto 52);
   tile_57_mult: IntMultiplierLUT_4x1_Freq300_uid243
      port map ( clk  => clk,
                 X => tile_57_X_c0,
                 Y => tile_57_Y_c0,
                 R => tile_57_output_c0);

   tile_57_filtered_output_c0 <= unsigned(tile_57_output_c0(3 downto 0));
   bh7_w98_2_c0 <= tile_57_filtered_output_c0(0);
   bh7_w99_1_c0 <= tile_57_filtered_output_c0(1);
   bh7_w100_1_c0 <= tile_57_filtered_output_c0(2);
   bh7_w101_0_c0 <= tile_57_filtered_output_c0(3);
   tile_58_X_c0 <= X(45 downto 42);
   tile_58_Y_c0 <= Y(52 downto 52);
   tile_58_mult: IntMultiplierLUT_4x1_Freq300_uid245
      port map ( clk  => clk,
                 X => tile_58_X_c0,
                 Y => tile_58_Y_c0,
                 R => tile_58_output_c0);

   tile_58_filtered_output_c0 <= unsigned(tile_58_output_c0(3 downto 0));
   bh7_w94_3_c0 <= tile_58_filtered_output_c0(0);
   bh7_w95_2_c0 <= tile_58_filtered_output_c0(1);
   bh7_w96_3_c0 <= tile_58_filtered_output_c0(2);
   bh7_w97_3_c0 <= tile_58_filtered_output_c0(3);
   tile_59_X_c0 <= X(41 downto 38);
   tile_59_Y_c0 <= Y(52 downto 52);
   tile_59_mult: IntMultiplierLUT_4x1_Freq300_uid247
      port map ( clk  => clk,
                 X => tile_59_X_c0,
                 Y => tile_59_Y_c0,
                 R => tile_59_output_c0);

   tile_59_filtered_output_c0 <= unsigned(tile_59_output_c0(3 downto 0));
   bh7_w90_3_c0 <= tile_59_filtered_output_c0(0);
   bh7_w91_3_c0 <= tile_59_filtered_output_c0(1);
   bh7_w92_2_c0 <= tile_59_filtered_output_c0(2);
   bh7_w93_3_c0 <= tile_59_filtered_output_c0(3);
   tile_60_X_c0 <= X(37 downto 34);
   tile_60_Y_c0 <= Y(52 downto 52);
   tile_60_mult: IntMultiplierLUT_4x1_Freq300_uid249
      port map ( clk  => clk,
                 X => tile_60_X_c0,
                 Y => tile_60_Y_c0,
                 R => tile_60_output_c0);

   tile_60_filtered_output_c0 <= unsigned(tile_60_output_c0(3 downto 0));
   bh7_w86_2_c0 <= tile_60_filtered_output_c0(0);
   bh7_w87_3_c0 <= tile_60_filtered_output_c0(1);
   bh7_w88_3_c0 <= tile_60_filtered_output_c0(2);
   bh7_w89_2_c0 <= tile_60_filtered_output_c0(3);
   tile_61_X_c0 <= X(50 downto 49);
   tile_61_Y_c0 <= Y(51 downto 50);
   tile_61_mult: IntMultiplierLUT_2x2_Freq300_uid251
      port map ( clk  => clk,
                 X => tile_61_X_c0,
                 Y => tile_61_Y_c0,
                 R => tile_61_output_c0);

   tile_61_filtered_output_c0 <= unsigned(tile_61_output_c0(3 downto 0));
   bh7_w99_2_c0 <= tile_61_filtered_output_c0(0);
   bh7_w100_2_c0 <= tile_61_filtered_output_c0(1);
   bh7_w101_1_c0 <= tile_61_filtered_output_c0(2);
   bh7_w102_1_c0 <= tile_61_filtered_output_c0(3);
   tile_62_X_c0 <= X(48 downto 46);
   tile_62_Y_c0 <= Y(51 downto 50);
   tile_62_mult: IntMultiplierLUT_3x2_Freq300_uid256
      port map ( clk  => clk,
                 X => tile_62_X_c0,
                 Y => tile_62_Y_c0,
                 R => tile_62_output_c0);

   tile_62_filtered_output_c0 <= unsigned(tile_62_output_c0(4 downto 0));
   bh7_w96_4_c0 <= tile_62_filtered_output_c0(0);
   bh7_w97_4_c0 <= tile_62_filtered_output_c0(1);
   bh7_w98_3_c0 <= tile_62_filtered_output_c0(2);
   bh7_w99_3_c0 <= tile_62_filtered_output_c0(3);
   bh7_w100_3_c0 <= tile_62_filtered_output_c0(4);
   tile_63_X_c0 <= X(45 downto 43);
   tile_63_Y_c0 <= Y(51 downto 50);
   tile_63_mult: IntMultiplierLUT_3x2_Freq300_uid261
      port map ( clk  => clk,
                 X => tile_63_X_c0,
                 Y => tile_63_Y_c0,
                 R => tile_63_output_c0);

   tile_63_filtered_output_c0 <= unsigned(tile_63_output_c0(4 downto 0));
   bh7_w93_4_c0 <= tile_63_filtered_output_c0(0);
   bh7_w94_4_c0 <= tile_63_filtered_output_c0(1);
   bh7_w95_3_c0 <= tile_63_filtered_output_c0(2);
   bh7_w96_5_c0 <= tile_63_filtered_output_c0(3);
   bh7_w97_5_c0 <= tile_63_filtered_output_c0(4);
   tile_64_X_c0 <= X(42 downto 40);
   tile_64_Y_c0 <= Y(51 downto 50);
   tile_64_mult: IntMultiplierLUT_3x2_Freq300_uid266
      port map ( clk  => clk,
                 X => tile_64_X_c0,
                 Y => tile_64_Y_c0,
                 R => tile_64_output_c0);

   tile_64_filtered_output_c0 <= unsigned(tile_64_output_c0(4 downto 0));
   bh7_w90_4_c0 <= tile_64_filtered_output_c0(0);
   bh7_w91_4_c0 <= tile_64_filtered_output_c0(1);
   bh7_w92_3_c0 <= tile_64_filtered_output_c0(2);
   bh7_w93_5_c0 <= tile_64_filtered_output_c0(3);
   bh7_w94_5_c0 <= tile_64_filtered_output_c0(4);
   tile_65_X_c0 <= X(39 downto 37);
   tile_65_Y_c0 <= Y(51 downto 50);
   tile_65_mult: IntMultiplierLUT_3x2_Freq300_uid271
      port map ( clk  => clk,
                 X => tile_65_X_c0,
                 Y => tile_65_Y_c0,
                 R => tile_65_output_c0);

   tile_65_filtered_output_c0 <= unsigned(tile_65_output_c0(4 downto 0));
   bh7_w87_4_c0 <= tile_65_filtered_output_c0(0);
   bh7_w88_4_c0 <= tile_65_filtered_output_c0(1);
   bh7_w89_3_c0 <= tile_65_filtered_output_c0(2);
   bh7_w90_5_c0 <= tile_65_filtered_output_c0(3);
   bh7_w91_5_c0 <= tile_65_filtered_output_c0(4);
   tile_66_X_c0 <= X(36 downto 34);
   tile_66_Y_c0 <= Y(51 downto 50);
   tile_66_mult: IntMultiplierLUT_3x2_Freq300_uid276
      port map ( clk  => clk,
                 X => tile_66_X_c0,
                 Y => tile_66_Y_c0,
                 R => tile_66_output_c0);

   tile_66_filtered_output_c0 <= unsigned(tile_66_output_c0(4 downto 0));
   bh7_w84_5_c0 <= tile_66_filtered_output_c0(0);
   bh7_w85_5_c0 <= tile_66_filtered_output_c0(1);
   bh7_w86_3_c0 <= tile_66_filtered_output_c0(2);
   bh7_w87_5_c0 <= tile_66_filtered_output_c0(3);
   bh7_w88_5_c0 <= tile_66_filtered_output_c0(4);
   tile_67_X_c0 <= X(50 downto 49);
   tile_67_Y_c0 <= Y(49 downto 48);
   tile_67_mult: IntMultiplierLUT_2x2_Freq300_uid281
      port map ( clk  => clk,
                 X => tile_67_X_c0,
                 Y => tile_67_Y_c0,
                 R => tile_67_output_c0);

   tile_67_filtered_output_c0 <= unsigned(tile_67_output_c0(3 downto 0));
   bh7_w97_6_c0 <= tile_67_filtered_output_c0(0);
   bh7_w98_4_c0 <= tile_67_filtered_output_c0(1);
   bh7_w99_4_c0 <= tile_67_filtered_output_c0(2);
   bh7_w100_4_c0 <= tile_67_filtered_output_c0(3);
   tile_68_X_c0 <= X(48 downto 46);
   tile_68_Y_c0 <= Y(49 downto 48);
   tile_68_mult: IntMultiplierLUT_3x2_Freq300_uid286
      port map ( clk  => clk,
                 X => tile_68_X_c0,
                 Y => tile_68_Y_c0,
                 R => tile_68_output_c0);

   tile_68_filtered_output_c0 <= unsigned(tile_68_output_c0(4 downto 0));
   bh7_w94_6_c0 <= tile_68_filtered_output_c0(0);
   bh7_w95_4_c0 <= tile_68_filtered_output_c0(1);
   bh7_w96_6_c0 <= tile_68_filtered_output_c0(2);
   bh7_w97_7_c0 <= tile_68_filtered_output_c0(3);
   bh7_w98_5_c0 <= tile_68_filtered_output_c0(4);
   tile_69_X_c0 <= X(45 downto 43);
   tile_69_Y_c0 <= Y(49 downto 48);
   tile_69_mult: IntMultiplierLUT_3x2_Freq300_uid291
      port map ( clk  => clk,
                 X => tile_69_X_c0,
                 Y => tile_69_Y_c0,
                 R => tile_69_output_c0);

   tile_69_filtered_output_c0 <= unsigned(tile_69_output_c0(4 downto 0));
   bh7_w91_6_c0 <= tile_69_filtered_output_c0(0);
   bh7_w92_4_c0 <= tile_69_filtered_output_c0(1);
   bh7_w93_6_c0 <= tile_69_filtered_output_c0(2);
   bh7_w94_7_c0 <= tile_69_filtered_output_c0(3);
   bh7_w95_5_c0 <= tile_69_filtered_output_c0(4);
   tile_70_X_c0 <= X(42 downto 40);
   tile_70_Y_c0 <= Y(49 downto 48);
   tile_70_mult: IntMultiplierLUT_3x2_Freq300_uid296
      port map ( clk  => clk,
                 X => tile_70_X_c0,
                 Y => tile_70_Y_c0,
                 R => tile_70_output_c0);

   tile_70_filtered_output_c0 <= unsigned(tile_70_output_c0(4 downto 0));
   bh7_w88_6_c0 <= tile_70_filtered_output_c0(0);
   bh7_w89_4_c0 <= tile_70_filtered_output_c0(1);
   bh7_w90_6_c0 <= tile_70_filtered_output_c0(2);
   bh7_w91_7_c0 <= tile_70_filtered_output_c0(3);
   bh7_w92_5_c0 <= tile_70_filtered_output_c0(4);
   tile_71_X_c0 <= X(39 downto 37);
   tile_71_Y_c0 <= Y(49 downto 48);
   tile_71_mult: IntMultiplierLUT_3x2_Freq300_uid301
      port map ( clk  => clk,
                 X => tile_71_X_c0,
                 Y => tile_71_Y_c0,
                 R => tile_71_output_c0);

   tile_71_filtered_output_c0 <= unsigned(tile_71_output_c0(4 downto 0));
   bh7_w85_6_c0 <= tile_71_filtered_output_c0(0);
   bh7_w86_4_c0 <= tile_71_filtered_output_c0(1);
   bh7_w87_6_c0 <= tile_71_filtered_output_c0(2);
   bh7_w88_7_c0 <= tile_71_filtered_output_c0(3);
   bh7_w89_5_c0 <= tile_71_filtered_output_c0(4);
   tile_72_X_c0 <= X(36 downto 34);
   tile_72_Y_c0 <= Y(49 downto 48);
   tile_72_mult: IntMultiplierLUT_3x2_Freq300_uid306
      port map ( clk  => clk,
                 X => tile_72_X_c0,
                 Y => tile_72_Y_c0,
                 R => tile_72_output_c0);

   tile_72_filtered_output_c0 <= unsigned(tile_72_output_c0(4 downto 0));
   bh7_w82_7_c0 <= tile_72_filtered_output_c0(0);
   bh7_w83_6_c0 <= tile_72_filtered_output_c0(1);
   bh7_w84_6_c0 <= tile_72_filtered_output_c0(2);
   bh7_w85_7_c0 <= tile_72_filtered_output_c0(3);
   bh7_w86_5_c0 <= tile_72_filtered_output_c0(4);
   tile_73_X_c0 <= X(52 downto 51);
   tile_73_Y_c0 <= Y(52 downto 51);
   tile_73_mult: IntMultiplierLUT_2x2_Freq300_uid311
      port map ( clk  => clk,
                 X => tile_73_X_c0,
                 Y => tile_73_Y_c0,
                 R => tile_73_output_c0);

   tile_73_filtered_output_c0 <= unsigned(tile_73_output_c0(3 downto 0));
   bh7_w102_2_c0 <= tile_73_filtered_output_c0(0);
   bh7_w103_0_c0 <= tile_73_filtered_output_c0(1);
   bh7_w104_0_c0 <= tile_73_filtered_output_c0(2);
   bh7_w105_0_c0 <= tile_73_filtered_output_c0(3);
   tile_74_X_c0 <= X(52 downto 51);
   tile_74_Y_c0 <= Y(50 downto 48);
   tile_74_mult: IntMultiplierLUT_2x3_Freq300_uid316
      port map ( clk  => clk,
                 X => tile_74_X_c0,
                 Y => tile_74_Y_c0,
                 R => tile_74_output_c0);

   tile_74_filtered_output_c0 <= unsigned(tile_74_output_c0(4 downto 0));
   bh7_w99_5_c0 <= tile_74_filtered_output_c0(0);
   bh7_w100_5_c0 <= tile_74_filtered_output_c0(1);
   bh7_w101_2_c0 <= tile_74_filtered_output_c0(2);
   bh7_w102_3_c0 <= tile_74_filtered_output_c0(3);
   bh7_w103_1_c0 <= tile_74_filtered_output_c0(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq300_uid322_bh7_uid323_In0_c0 <= "" & bh7_w49_4_c0 & "0" & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid323_In1_c0 <= "" & bh7_w50_4_c0 & bh7_w50_5_c0;
   bh7_w49_5_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0(0);
   bh7_w50_6_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0(1);
   bh7_w51_8_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid323: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid323_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid323_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_copy324_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_copy324_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid327_In0_c0 <= "" & bh7_w51_2_c0 & bh7_w51_5_c0 & bh7_w51_6_c0 & bh7_w51_7_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid327_In1_c0 <= "" & bh7_w52_2_c0;
   bh7_w51_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0(0);
   bh7_w52_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0(1);
   bh7_w53_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid327: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid327_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid327_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_copy328_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_copy328_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid329_In0_c0 <= "" & bh7_w52_5_c0 & bh7_w52_6_c0 & bh7_w52_7_c0 & bh7_w52_8_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid329_In1_c0 <= "" & bh7_w53_2_c0;
   bh7_w52_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0(0);
   bh7_w53_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0(1);
   bh7_w54_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid329: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid329_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid329_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_copy330_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_copy330_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid331_In0_c0 <= "" & bh7_w53_5_c0 & bh7_w53_6_c0 & bh7_w53_7_c0 & bh7_w53_8_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid331_In1_c0 <= "" & bh7_w54_2_c0;
   bh7_w53_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0(0);
   bh7_w54_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0(1);
   bh7_w55_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid331: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid331_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid331_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_copy332_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_copy332_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid335_In0_c0 <= "" & bh7_w54_3_c0 & bh7_w54_6_c0 & bh7_w54_7_c0 & bh7_w54_8_c0 & bh7_w54_9_c0 & bh7_w54_10_c0;
   bh7_w54_13_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0(0);
   bh7_w55_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0(1);
   bh7_w56_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid335: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid335_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_copy336_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_copy336_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid337_In0_c0 <= "" & bh7_w55_2_c0 & bh7_w55_3_c0 & bh7_w55_6_c0 & bh7_w55_7_c0 & bh7_w55_8_c0 & bh7_w55_9_c0;
   bh7_w55_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0(0);
   bh7_w56_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0(1);
   bh7_w57_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid337: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid337_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_copy338_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_copy338_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid339_In0_c0 <= "" & bh7_w56_2_c0 & bh7_w56_5_c0 & bh7_w56_6_c0 & bh7_w56_7_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid339_In1_c0 <= "" & bh7_w57_2_c0;
   bh7_w56_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0(0);
   bh7_w57_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0(1);
   bh7_w58_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid339: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid339_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid339_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_copy340_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_copy340_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid341_In0_c0 <= "" & bh7_w57_3_c0 & bh7_w57_6_c0 & bh7_w57_7_c0 & bh7_w57_8_c0 & bh7_w57_9_c0 & bh7_w57_10_c0;
   bh7_w57_13_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0(0);
   bh7_w58_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0(1);
   bh7_w59_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid341: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid341_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_copy342_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_copy342_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid343_In0_c0 <= "" & bh7_w58_1_c0 & bh7_w58_2_c0 & bh7_w58_6_c0 & bh7_w58_7_c0 & bh7_w58_8_c0 & bh7_w58_9_c0;
   bh7_w58_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0(0);
   bh7_w59_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0(1);
   bh7_w60_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid343: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid343_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_copy344_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_copy344_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid345_In0_c0 <= "" & bh7_w59_1_c0 & bh7_w59_5_c0 & bh7_w59_6_c0 & bh7_w59_7_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid345_In1_c0 <= "" & bh7_w60_1_c0;
   bh7_w59_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0(0);
   bh7_w60_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0(1);
   bh7_w61_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid345: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid345_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid345_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_copy346_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_copy346_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid347_In0_c0 <= "" & bh7_w60_2_c0 & bh7_w60_6_c0 & bh7_w60_7_c0 & bh7_w60_8_c0 & bh7_w60_9_c0 & bh7_w60_10_c0;
   bh7_w60_13_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0(0);
   bh7_w61_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0(1);
   bh7_w62_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid347: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid347_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_copy348_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_copy348_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid349_In0_c0 <= "" & bh7_w61_1_c0 & bh7_w61_2_c0 & bh7_w61_6_c0 & bh7_w61_7_c0 & bh7_w61_8_c0 & bh7_w61_9_c0;
   bh7_w61_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0(0);
   bh7_w62_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0(1);
   bh7_w63_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid349: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid349_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_copy350_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_copy350_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid351_In0_c0 <= "" & bh7_w62_1_c0 & bh7_w62_5_c0 & bh7_w62_6_c0 & bh7_w62_7_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid351_In1_c0 <= "" & bh7_w63_1_c0;
   bh7_w62_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0(0);
   bh7_w63_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0(1);
   bh7_w64_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid351: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid351_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid351_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_copy352_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_copy352_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid353_In0_c0 <= "" & bh7_w63_2_c0 & bh7_w63_6_c0 & bh7_w63_7_c0 & bh7_w63_8_c0 & bh7_w63_9_c0 & bh7_w63_10_c0;
   bh7_w63_13_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0(0);
   bh7_w64_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0(1);
   bh7_w65_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid353: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid353_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_copy354_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_copy354_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid355_In0_c0 <= "" & bh7_w64_1_c0 & bh7_w64_2_c0 & bh7_w64_6_c0 & bh7_w64_7_c0 & bh7_w64_8_c0 & bh7_w64_9_c0;
   bh7_w64_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0(0);
   bh7_w65_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0(1);
   bh7_w66_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid355: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid355_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_copy356_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_copy356_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid357_In0_c0 <= "" & bh7_w65_1_c0 & bh7_w65_4_c0 & bh7_w65_5_c0 & bh7_w65_6_c0 & bh7_w65_7_c0 & bh7_w65_8_c0;
   bh7_w65_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0(0);
   bh7_w66_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0(1);
   bh7_w67_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid357: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid357_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_copy358_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_copy358_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid359_In0_c0 <= "" & bh7_w66_1_c0 & bh7_w66_2_c0 & bh7_w66_5_c0 & bh7_w66_6_c0 & bh7_w66_7_c0 & bh7_w66_8_c0;
   bh7_w66_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0(0);
   bh7_w67_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0(1);
   bh7_w68_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid359: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid359_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_copy360_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_copy360_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid361_In0_c0 <= "" & bh7_w67_1_c0 & bh7_w67_2_c0 & bh7_w67_5_c0 & bh7_w67_6_c0 & bh7_w67_7_c0 & bh7_w67_8_c0;
   bh7_w67_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0(0);
   bh7_w68_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0(1);
   bh7_w69_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid361: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid361_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_copy362_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_copy362_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid363_In0_c0 <= "" & bh7_w68_1_c0 & bh7_w68_4_c0 & bh7_w68_5_c0 & bh7_w68_6_c0 & bh7_w68_7_c0 & bh7_w68_8_c0;
   bh7_w68_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0(0);
   bh7_w69_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0(1);
   bh7_w70_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid363: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid363_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_copy364_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_copy364_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid365_In0_c0 <= "" & bh7_w69_1_c0 & bh7_w69_2_c0 & bh7_w69_5_c0 & bh7_w69_6_c0 & bh7_w69_7_c0 & bh7_w69_8_c0;
   bh7_w69_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0(0);
   bh7_w70_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0(1);
   bh7_w71_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid365: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid365_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_copy366_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_copy366_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid367_In0_c0 <= "" & bh7_w70_1_c0 & bh7_w70_2_c0 & bh7_w70_5_c0 & bh7_w70_6_c0 & bh7_w70_7_c0 & bh7_w70_8_c0;
   bh7_w70_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0(0);
   bh7_w71_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0(1);
   bh7_w72_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid367: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid367_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_copy368_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_copy368_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid369_In0_c0 <= "" & bh7_w71_1_c0 & bh7_w71_4_c0 & bh7_w71_5_c0 & bh7_w71_6_c0 & bh7_w71_7_c0 & bh7_w71_8_c0;
   bh7_w71_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0(0);
   bh7_w72_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0(1);
   bh7_w73_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid369: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid369_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_copy370_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_copy370_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid371_In0_c0 <= "" & bh7_w72_1_c0 & bh7_w72_2_c0 & bh7_w72_5_c0 & bh7_w72_6_c0 & bh7_w72_7_c0 & bh7_w72_8_c0;
   bh7_w72_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0(0);
   bh7_w73_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0(1);
   bh7_w74_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid371: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid371_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_copy372_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_copy372_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid373_In0_c0 <= "" & bh7_w73_1_c0 & bh7_w73_2_c0 & bh7_w73_5_c0 & bh7_w73_6_c0 & bh7_w73_7_c0 & bh7_w73_8_c0;
   bh7_w73_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0(0);
   bh7_w74_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0(1);
   bh7_w75_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid373: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid373_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_copy374_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_copy374_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid375_In0_c0 <= "" & bh7_w74_1_c0 & bh7_w74_4_c0 & bh7_w74_5_c0 & bh7_w74_6_c0 & bh7_w74_7_c0 & bh7_w74_8_c0;
   bh7_w74_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0(0);
   bh7_w75_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0(1);
   bh7_w76_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid375: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid375_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_copy376_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_copy376_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid377_In0_c0 <= "" & bh7_w75_0_c0 & bh7_w75_3_c0 & bh7_w75_4_c0 & bh7_w75_5_c0 & bh7_w75_6_c0 & bh7_w75_7_c0;
   bh7_w75_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0(0);
   bh7_w76_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0(1);
   bh7_w77_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid377: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid377_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_copy378_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_copy378_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid379_In0_c0 <= "" & bh7_w76_0_c0 & bh7_w76_3_c0 & bh7_w76_4_c0 & bh7_w76_5_c0 & bh7_w76_6_c0 & bh7_w76_7_c0;
   bh7_w76_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0(0);
   bh7_w77_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0(1);
   bh7_w78_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid379: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid379_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_copy380_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_copy380_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid381_In0_c0 <= "" & bh7_w77_2_c0 & bh7_w77_3_c0 & bh7_w77_4_c0 & bh7_w77_5_c0 & bh7_w77_6_c0 & bh7_w77_7_c0;
   bh7_w77_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0(0);
   bh7_w78_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0(1);
   bh7_w79_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid381: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid381_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_copy382_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_copy382_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid383_In0_c0 <= "" & bh7_w78_2_c0 & bh7_w78_3_c0 & bh7_w78_4_c0 & bh7_w78_5_c0 & bh7_w78_6_c0 & bh7_w78_7_c0;
   bh7_w78_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0(0);
   bh7_w79_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0(1);
   bh7_w80_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid383: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid383_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_copy384_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_copy384_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid385_In0_c0 <= "" & bh7_w79_2_c0 & bh7_w79_3_c0 & bh7_w79_4_c0 & bh7_w79_5_c0 & bh7_w79_6_c0 & bh7_w79_7_c0;
   bh7_w79_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0(0);
   bh7_w80_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0(1);
   bh7_w81_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid385: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid385_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_copy386_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_copy386_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid387_In0_c0 <= "" & bh7_w80_2_c0 & bh7_w80_3_c0 & bh7_w80_4_c0 & bh7_w80_5_c0 & bh7_w80_6_c0 & bh7_w80_7_c0;
   bh7_w80_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0(0);
   bh7_w81_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0(1);
   bh7_w82_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid387: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid387_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_copy388_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_copy388_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid389_In0_c0 <= "" & bh7_w81_2_c0 & bh7_w81_3_c0 & bh7_w81_4_c0 & bh7_w81_5_c0 & bh7_w81_6_c0 & bh7_w81_7_c0;
   bh7_w81_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0(0);
   bh7_w82_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0(1);
   bh7_w83_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid389: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid389_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_copy390_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_copy390_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid391_In0_c0 <= "" & bh7_w82_1_c0 & bh7_w82_2_c0 & bh7_w82_3_c0 & bh7_w82_4_c0 & bh7_w82_5_c0 & bh7_w82_6_c0;
   bh7_w82_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0(0);
   bh7_w83_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0(1);
   bh7_w84_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid391: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid391_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_copy392_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_copy392_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid393_In0_c0 <= "" & bh7_w83_1_c0 & bh7_w83_2_c0 & bh7_w83_3_c0 & bh7_w83_4_c0 & bh7_w83_5_c0 & bh7_w83_6_c0;
   bh7_w83_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0(0);
   bh7_w84_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0(1);
   bh7_w85_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid393: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid393_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_copy394_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_copy394_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid395_In0_c0 <= "" & bh7_w84_1_c0 & bh7_w84_2_c0 & bh7_w84_3_c0 & bh7_w84_4_c0 & bh7_w84_5_c0 & bh7_w84_6_c0;
   bh7_w84_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0(0);
   bh7_w85_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0(1);
   bh7_w86_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid395: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid395_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_copy396_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_copy396_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid397_In0_c0 <= "" & bh7_w85_1_c0 & bh7_w85_2_c0 & bh7_w85_3_c0 & bh7_w85_4_c0 & bh7_w85_5_c0 & bh7_w85_6_c0;
   bh7_w85_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0(0);
   bh7_w86_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0(1);
   bh7_w87_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid397: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid397_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_copy398_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_copy398_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid401_In0_c0 <= "" & bh7_w86_1_c0 & bh7_w86_2_c0 & bh7_w86_3_c0 & bh7_w86_4_c0 & bh7_w86_5_c0;
   bh7_w86_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0(0);
   bh7_w87_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0(1);
   bh7_w88_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid401: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid401_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_copy402_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_copy402_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid403_In0_c0 <= "" & bh7_w87_1_c0 & bh7_w87_2_c0 & bh7_w87_3_c0 & bh7_w87_4_c0 & bh7_w87_5_c0 & bh7_w87_6_c0;
   bh7_w87_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0(0);
   bh7_w88_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0(1);
   bh7_w89_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid403: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid403_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_copy404_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_copy404_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid405_In0_c0 <= "" & bh7_w88_1_c0 & bh7_w88_2_c0 & bh7_w88_3_c0 & bh7_w88_4_c0 & bh7_w88_5_c0 & bh7_w88_6_c0;
   bh7_w88_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0(0);
   bh7_w89_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0(1);
   bh7_w90_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid405: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid405_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_copy406_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_copy406_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid407_In0_c0 <= "" & bh7_w89_1_c0 & bh7_w89_2_c0 & bh7_w89_3_c0 & bh7_w89_4_c0 & bh7_w89_5_c0;
   bh7_w89_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0(0);
   bh7_w90_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0(1);
   bh7_w91_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid407: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid407_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_copy408_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_copy408_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid409_In0_c0 <= "" & bh7_w90_1_c0 & bh7_w90_2_c0 & bh7_w90_3_c0 & bh7_w90_4_c0 & bh7_w90_5_c0 & bh7_w90_6_c0;
   bh7_w90_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0(0);
   bh7_w91_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0(1);
   bh7_w92_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid409: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid409_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_copy410_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_copy410_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid411_In0_c0 <= "" & bh7_w91_1_c0 & bh7_w91_2_c0 & bh7_w91_3_c0 & bh7_w91_4_c0 & bh7_w91_5_c0 & bh7_w91_6_c0;
   bh7_w91_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0(0);
   bh7_w92_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0(1);
   bh7_w93_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid411: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid411_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_copy412_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_copy412_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid413_In0_c0 <= "" & bh7_w92_1_c0 & bh7_w92_2_c0 & bh7_w92_3_c0 & bh7_w92_4_c0 & bh7_w92_5_c0;
   bh7_w92_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0(0);
   bh7_w93_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0(1);
   bh7_w94_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid413: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid413_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_copy414_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_copy414_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid415_In0_c0 <= "" & bh7_w93_1_c0 & bh7_w93_2_c0 & bh7_w93_3_c0 & bh7_w93_4_c0 & bh7_w93_5_c0 & bh7_w93_6_c0;
   bh7_w93_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0(0);
   bh7_w94_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0(1);
   bh7_w95_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid415: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid415_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_copy416_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_copy416_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid417_In0_c0 <= "" & bh7_w94_1_c0 & bh7_w94_2_c0 & bh7_w94_3_c0 & bh7_w94_4_c0 & bh7_w94_5_c0 & bh7_w94_6_c0;
   bh7_w94_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0(0);
   bh7_w95_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0(1);
   bh7_w96_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid417: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid417_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_copy418_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_copy418_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid419_In0_c0 <= "" & bh7_w95_1_c0 & bh7_w95_2_c0 & bh7_w95_3_c0 & bh7_w95_4_c0 & bh7_w95_5_c0;
   bh7_w95_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0(0);
   bh7_w96_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0(1);
   bh7_w97_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid419: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid419_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_copy420_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_copy420_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid421_In0_c0 <= "" & bh7_w96_1_c0 & bh7_w96_2_c0 & bh7_w96_3_c0 & bh7_w96_4_c0 & bh7_w96_5_c0 & bh7_w96_6_c0;
   bh7_w96_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0(0);
   bh7_w97_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0(1);
   bh7_w98_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid421: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid421_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_copy422_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_copy422_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid423_In0_c0 <= "" & bh7_w97_1_c0 & bh7_w97_2_c0 & bh7_w97_3_c0 & bh7_w97_4_c0 & bh7_w97_5_c0 & bh7_w97_6_c0;
   bh7_w97_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0(0);
   bh7_w98_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0(1);
   bh7_w99_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid423: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid423_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_copy424_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_copy424_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid425_In0_c0 <= "" & bh7_w98_1_c0 & bh7_w98_2_c0 & bh7_w98_3_c0 & bh7_w98_4_c0 & bh7_w98_5_c0;
   bh7_w98_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0(0);
   bh7_w99_7_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0(1);
   bh7_w100_6_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid425: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid425_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_copy426_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_copy426_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid427_In0_c0 <= "" & bh7_w99_0_c0 & bh7_w99_1_c0 & bh7_w99_2_c0 & bh7_w99_3_c0 & bh7_w99_4_c0 & bh7_w99_5_c0;
   bh7_w99_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0(0);
   bh7_w100_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0(1);
   bh7_w101_3_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid427: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid427_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_copy428_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_copy428_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid429_In0_c0 <= "" & bh7_w100_0_c0 & bh7_w100_1_c0 & bh7_w100_2_c0 & bh7_w100_3_c0 & bh7_w100_4_c0 & bh7_w100_5_c0;
   bh7_w100_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0(0);
   bh7_w101_4_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0(1);
   bh7_w102_4_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid429: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid429_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_copy430_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_copy430_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid433_In0_c0 <= "" & bh7_w101_0_c0 & bh7_w101_1_c0 & bh7_w101_2_c0;
   bh7_w101_5_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_c0(0);
   bh7_w102_5_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid433: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid433_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_copy434_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_copy434_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid435_In0_c0 <= "" & bh7_w102_0_c0 & bh7_w102_1_c0 & bh7_w102_2_c0 & bh7_w102_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid435_In1_c0 <= "" & bh7_w103_0_c0;
   bh7_w102_6_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0(0);
   bh7_w103_2_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0(1);
   bh7_w104_1_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid435: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid435_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid435_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_copy436_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_copy436_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid437_In0_c0 <= "" & bh7_w51_9_c0 & bh7_w51_8_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid437_In1_c0 <= "" & bh7_w52_10_c0 & bh7_w52_9_c0;
   bh7_w51_10_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0(0);
   bh7_w52_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0(1);
   bh7_w53_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid437: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid437_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid437_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_copy438_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_copy438_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid439_In0_c0 <= "" & bh7_w53_11_c0 & bh7_w53_10_c0 & bh7_w53_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid439_In1_c0 <= "" & bh7_w54_12_c0 & bh7_w54_11_c0;
   bh7_w53_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0(0);
   bh7_w54_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0(1);
   bh7_w55_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid439: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid439_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid439_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_copy440_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_copy440_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid441_In0_c0 <= "" & bh7_w55_10_c0 & bh7_w55_12_c0 & bh7_w55_11_c0;
   bh7_w55_14_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_c0(0);
   bh7_w56_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid441: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid441_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_copy442_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_copy442_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid443_In0_c0 <= "" & bh7_w56_8_c0 & bh7_w56_11_c0 & bh7_w56_10_c0 & bh7_w56_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid443_In1_c0 <= "" & "0";
   bh7_w56_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0(0);
   bh7_w57_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0(1);
   bh7_w58_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid443: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid443_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid443_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_copy444_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_copy444_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid445_In0_c0 <= "" & bh7_w57_12_c0 & bh7_w57_13_c0 & bh7_w57_11_c0;
   bh7_w57_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_c0(0);
   bh7_w58_14_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid445: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid445_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_copy446_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_copy446_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid447_In0_c0 <= "" & bh7_w58_10_c0 & bh7_w58_12_c0 & bh7_w58_11_c0;
   bh7_w58_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_c0(0);
   bh7_w59_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid447: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid447_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_copy448_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_copy448_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid449_In0_c0 <= "" & bh7_w59_8_c0 & bh7_w59_11_c0 & bh7_w59_10_c0 & bh7_w59_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid449_In1_c0 <= "" & "0";
   bh7_w59_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0(0);
   bh7_w60_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0(1);
   bh7_w61_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid449: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid449_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid449_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_copy450_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_copy450_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid451_In0_c0 <= "" & bh7_w60_12_c0 & bh7_w60_13_c0 & bh7_w60_11_c0;
   bh7_w60_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_c0(0);
   bh7_w61_14_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid451: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid451_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_copy452_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_copy452_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid453_In0_c0 <= "" & bh7_w61_10_c0 & bh7_w61_12_c0 & bh7_w61_11_c0;
   bh7_w61_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_c0(0);
   bh7_w62_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid453: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid453_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_copy454_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_copy454_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid455_In0_c0 <= "" & bh7_w62_8_c0 & bh7_w62_11_c0 & bh7_w62_10_c0 & bh7_w62_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid455_In1_c0 <= "" & "0";
   bh7_w62_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0(0);
   bh7_w63_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0(1);
   bh7_w64_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid455: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid455_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid455_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_copy456_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_copy456_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid457_In0_c0 <= "" & bh7_w63_12_c0 & bh7_w63_13_c0 & bh7_w63_11_c0;
   bh7_w63_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_c0(0);
   bh7_w64_14_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid457: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid457_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_copy458_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_copy458_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid459_In0_c0 <= "" & bh7_w64_10_c0 & bh7_w64_12_c0 & bh7_w64_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid459_In1_c0 <= "" & bh7_w65_11_c0 & bh7_w65_10_c0;
   bh7_w64_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0(0);
   bh7_w65_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0(1);
   bh7_w66_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid459: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid459_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid459_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_copy460_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_copy460_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid461_In0_c0 <= "" & bh7_w66_9_c0 & bh7_w66_12_c0 & bh7_w66_11_c0 & bh7_w66_10_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid461_In1_c0 <= "" & "0";
   bh7_w66_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0(0);
   bh7_w67_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0(1);
   bh7_w68_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid461: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid461_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid461_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_copy462_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_copy462_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid463_In0_c0 <= "" & bh7_w67_11_c0 & bh7_w67_10_c0 & bh7_w67_9_c0;
   bh7_w67_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_c0(0);
   bh7_w68_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid463: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid463_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_copy464_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_copy464_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid465_In0_c0 <= "" & bh7_w68_11_c0 & bh7_w68_10_c0 & bh7_w68_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid465_In1_c0 <= "" & bh7_w69_11_c0 & bh7_w69_10_c0;
   bh7_w68_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0(0);
   bh7_w69_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0(1);
   bh7_w70_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid465: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid465_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid465_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_copy466_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_copy466_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid467_In0_c0 <= "" & bh7_w70_11_c0 & bh7_w70_10_c0 & bh7_w70_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid467_In1_c0 <= "" & bh7_w71_11_c0 & bh7_w71_10_c0;
   bh7_w70_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0(0);
   bh7_w71_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0(1);
   bh7_w72_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid467: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid467_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid467_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_copy468_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_copy468_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid469_In0_c0 <= "" & bh7_w72_11_c0 & bh7_w72_10_c0 & bh7_w72_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid469_In1_c0 <= "" & bh7_w73_11_c0 & bh7_w73_10_c0;
   bh7_w72_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0(0);
   bh7_w73_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0(1);
   bh7_w74_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid469: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid469_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid469_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_copy470_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_copy470_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid471_In0_c0 <= "" & bh7_w74_11_c0 & bh7_w74_10_c0 & bh7_w74_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid471_In1_c0 <= "" & bh7_w75_10_c0 & bh7_w75_9_c0;
   bh7_w74_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0(0);
   bh7_w75_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0(1);
   bh7_w76_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid471: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid471_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid471_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_copy472_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_copy472_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid473_In0_c0 <= "" & bh7_w76_10_c0 & bh7_w76_9_c0 & bh7_w76_8_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid473_In1_c0 <= "" & bh7_w77_10_c0 & bh7_w77_9_c0;
   bh7_w76_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0(0);
   bh7_w77_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0(1);
   bh7_w78_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid473: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid473_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid473_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_copy474_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_copy474_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid475_In0_c0 <= "" & bh7_w78_10_c0 & bh7_w78_9_c0 & bh7_w78_8_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid475_In1_c0 <= "" & bh7_w79_10_c0 & bh7_w79_9_c0;
   bh7_w78_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0(0);
   bh7_w79_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0(1);
   bh7_w80_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid475: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid475_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid475_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_copy476_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_copy476_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid477_In0_c0 <= "" & bh7_w80_10_c0 & bh7_w80_9_c0 & bh7_w80_8_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid477_In1_c0 <= "" & bh7_w81_10_c0 & bh7_w81_9_c0;
   bh7_w80_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0(0);
   bh7_w81_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0(1);
   bh7_w82_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid477: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid477_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid477_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_copy478_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_copy478_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid479_In0_c0 <= "" & bh7_w82_7_c0 & bh7_w82_10_c0 & bh7_w82_9_c0 & bh7_w82_8_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid479_In1_c0 <= "" & "0";
   bh7_w82_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0(0);
   bh7_w83_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0(1);
   bh7_w84_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid479: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid479_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid479_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_copy480_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_copy480_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid481_In0_c0 <= "" & bh7_w83_9_c0 & bh7_w83_8_c0 & bh7_w83_7_c0;
   bh7_w83_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_c0(0);
   bh7_w84_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid481: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid481_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_copy482_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_copy482_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid483_In0_c0 <= "" & bh7_w84_9_c0 & bh7_w84_8_c0 & bh7_w84_7_c0;
   bh7_w84_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_c0(0);
   bh7_w85_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid483: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid483_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_copy484_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_copy484_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid485_In0_c0 <= "" & bh7_w85_7_c0 & bh7_w85_10_c0 & bh7_w85_9_c0 & bh7_w85_8_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid485_In1_c0 <= "" & "0";
   bh7_w85_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0(0);
   bh7_w86_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0(1);
   bh7_w87_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid485: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid485_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid485_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_copy486_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_copy486_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid487_In0_c0 <= "" & bh7_w86_8_c0 & bh7_w86_7_c0 & bh7_w86_6_c0;
   bh7_w86_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_c0(0);
   bh7_w87_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid487: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid487_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_copy488_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_copy488_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid489_In0_c0 <= "" & bh7_w87_8_c0 & bh7_w87_9_c0 & bh7_w87_7_c0;
   bh7_w87_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_c0(0);
   bh7_w88_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid489: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid489_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_copy490_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_copy490_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid491_In0_c0 <= "" & bh7_w88_7_c0 & bh7_w88_8_c0 & bh7_w88_10_c0 & bh7_w88_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid491_In1_c0 <= "" & "0";
   bh7_w88_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0(0);
   bh7_w89_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0(1);
   bh7_w90_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid491: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid491_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid491_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_copy492_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_copy492_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid493_In0_c0 <= "" & bh7_w89_8_c0 & bh7_w89_7_c0 & bh7_w89_6_c0;
   bh7_w89_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_c0(0);
   bh7_w90_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid493: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid493_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_copy494_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_copy494_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid495_In0_c0 <= "" & bh7_w90_8_c0 & bh7_w90_9_c0 & bh7_w90_7_c0;
   bh7_w90_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_c0(0);
   bh7_w91_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid495: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid495_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_copy496_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_copy496_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid497_In0_c0 <= "" & bh7_w91_7_c0 & bh7_w91_8_c0 & bh7_w91_10_c0 & bh7_w91_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid497_In1_c0 <= "" & "0";
   bh7_w91_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0(0);
   bh7_w92_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0(1);
   bh7_w93_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid497: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid497_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid497_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_copy498_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_copy498_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid499_In0_c0 <= "" & bh7_w92_8_c0 & bh7_w92_7_c0 & bh7_w92_6_c0;
   bh7_w92_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_c0(0);
   bh7_w93_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid499: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid499_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_copy500_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_copy500_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid501_In0_c0 <= "" & bh7_w93_8_c0 & bh7_w93_9_c0 & bh7_w93_7_c0;
   bh7_w93_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_c0(0);
   bh7_w94_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid501: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid501_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_copy502_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_copy502_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid503_In0_c0 <= "" & bh7_w94_7_c0 & bh7_w94_8_c0 & bh7_w94_10_c0 & bh7_w94_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid503_In1_c0 <= "" & "0";
   bh7_w94_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0(0);
   bh7_w95_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0(1);
   bh7_w96_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid503: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid503_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid503_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_copy504_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_copy504_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid505_In0_c0 <= "" & bh7_w95_8_c0 & bh7_w95_7_c0 & bh7_w95_6_c0;
   bh7_w95_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_c0(0);
   bh7_w96_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid505: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid505_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_copy506_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_copy506_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid507_In0_c0 <= "" & bh7_w96_8_c0 & bh7_w96_9_c0 & bh7_w96_7_c0;
   bh7_w96_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_c0(0);
   bh7_w97_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid507: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid507_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_copy508_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_copy508_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid509_In0_c0 <= "" & bh7_w97_7_c0 & bh7_w97_8_c0 & bh7_w97_10_c0 & bh7_w97_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid509_In1_c0 <= "" & "0";
   bh7_w97_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0(0);
   bh7_w98_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0(1);
   bh7_w99_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid509: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid509_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid509_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_copy510_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_copy510_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid511_In0_c0 <= "" & bh7_w98_8_c0 & bh7_w98_7_c0 & bh7_w98_6_c0;
   bh7_w98_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_c0(0);
   bh7_w99_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid511: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid511_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_copy512_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_copy512_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid513_In0_c0 <= "" & bh7_w99_7_c0 & bh7_w99_8_c0 & bh7_w99_6_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid513_In1_c0 <= "" & bh7_w100_6_c0 & bh7_w100_8_c0;
   bh7_w99_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0(0);
   bh7_w100_9_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0(1);
   bh7_w101_6_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid513: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid513_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid513_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_copy514_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_copy514_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid515_In0_c0 <= "" & bh7_w101_5_c0 & bh7_w101_4_c0 & bh7_w101_3_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid515_In1_c0 <= "" & bh7_w102_6_c0 & bh7_w102_5_c0;
   bh7_w101_7_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0(0);
   bh7_w102_7_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0(1);
   bh7_w103_3_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid515: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid515_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid515_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_copy516_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_copy516_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid517_In0_c0 <= "" & bh7_w103_1_c0 & bh7_w103_2_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid517_In1_c0 <= "" & bh7_w104_0_c0 & bh7_w104_1_c0;
   bh7_w103_4_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0(0);
   bh7_w104_2_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0(1);
   bh7_w105_1_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid517: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid517_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid517_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_copy518_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_copy518_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid519_In0_c0 <= "" & bh7_w53_13_c0 & bh7_w53_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid519_In1_c0 <= "" & bh7_w54_13_c0 & bh7_w54_14_c0;
   bh7_w53_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0(0);
   bh7_w54_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0(1);
   bh7_w55_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid519: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid519_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid519_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_copy520_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_copy520_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid521_In0_c0 <= "" & bh7_w55_13_c0 & bh7_w55_14_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid521_In1_c0 <= "" & bh7_w56_13_c0 & bh7_w56_12_c0;
   bh7_w55_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0(0);
   bh7_w56_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0(1);
   bh7_w57_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid521: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid521_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid521_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_copy522_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_copy522_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid523_In0_c0 <= "" & bh7_w57_14_c0 & bh7_w57_15_c0 & "0";
   bh7_w57_17_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_c0(0);
   bh7_w58_16_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid523: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid523_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_copy524_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_copy524_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid525_In0_c0 <= "" & bh7_w58_13_c0 & bh7_w58_15_c0 & bh7_w58_14_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid525_In1_c0 <= "" & bh7_w59_13_c0 & bh7_w59_12_c0;
   bh7_w58_17_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0(0);
   bh7_w59_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0(1);
   bh7_w60_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid525: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid525_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid525_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_copy526_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_copy526_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid527_In0_c0 <= "" & bh7_w60_14_c0 & bh7_w60_15_c0 & "0";
   bh7_w60_17_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_c0(0);
   bh7_w61_16_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid527: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid527_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_copy528_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_copy528_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid529_In0_c0 <= "" & bh7_w61_13_c0 & bh7_w61_15_c0 & bh7_w61_14_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid529_In1_c0 <= "" & bh7_w62_13_c0 & bh7_w62_12_c0;
   bh7_w61_17_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0(0);
   bh7_w62_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0(1);
   bh7_w63_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid529: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid529_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid529_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_copy530_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_copy530_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid531_In0_c0 <= "" & bh7_w63_14_c0 & bh7_w63_15_c0 & "0";
   bh7_w63_17_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_c0(0);
   bh7_w64_16_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid531: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid531_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_copy532_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_copy532_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid533_In0_c0 <= "" & bh7_w64_13_c0 & bh7_w64_15_c0 & bh7_w64_14_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid533_In1_c0 <= "" & bh7_w65_9_c0 & bh7_w65_12_c0;
   bh7_w64_17_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0(0);
   bh7_w65_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0(1);
   bh7_w66_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid533: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid533_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid533_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_copy534_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_copy534_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid535_In0_c0 <= "" & bh7_w66_14_c0 & bh7_w66_13_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid535_In1_c0 <= "" & bh7_w67_12_c0 & bh7_w67_13_c0;
   bh7_w66_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0(0);
   bh7_w67_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0(1);
   bh7_w68_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid535: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid535_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid535_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_copy536_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_copy536_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid537_In0_c0 <= "" & bh7_w68_12_c0 & bh7_w68_14_c0 & bh7_w68_13_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid537_In1_c0 <= "" & bh7_w69_9_c0 & bh7_w69_12_c0;
   bh7_w68_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0(0);
   bh7_w69_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0(1);
   bh7_w70_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid537: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid537_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid537_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_copy538_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_copy538_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid539_In0_c0 <= "" & bh7_w70_13_c0 & bh7_w70_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid539_In1_c0 <= "" & bh7_w71_9_c0 & bh7_w71_12_c0;
   bh7_w70_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0(0);
   bh7_w71_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0(1);
   bh7_w72_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid539: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid539_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid539_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_copy540_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_copy540_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid541_In0_c0 <= "" & bh7_w72_13_c0 & bh7_w72_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid541_In1_c0 <= "" & bh7_w73_9_c0 & bh7_w73_12_c0;
   bh7_w72_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0(0);
   bh7_w73_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0(1);
   bh7_w74_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid541: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid541_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid541_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_copy542_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_copy542_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid543_In0_c0 <= "" & bh7_w74_13_c0 & bh7_w74_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid543_In1_c0 <= "" & bh7_w75_8_c0 & bh7_w75_11_c0;
   bh7_w74_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0(0);
   bh7_w75_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0(1);
   bh7_w76_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid543: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid543_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid543_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_copy544_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_copy544_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid545_In0_c0 <= "" & bh7_w76_12_c0 & bh7_w76_11_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid545_In1_c0 <= "" & bh7_w77_8_c0 & bh7_w77_11_c0;
   bh7_w76_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0(0);
   bh7_w77_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0(1);
   bh7_w78_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid545: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid545_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid545_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_copy546_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_copy546_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid547_In0_c0 <= "" & bh7_w78_12_c0 & bh7_w78_11_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid547_In1_c0 <= "" & bh7_w79_8_c0 & bh7_w79_11_c0;
   bh7_w78_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0(0);
   bh7_w79_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0(1);
   bh7_w80_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid547: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid547_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid547_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_copy548_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_copy548_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid549_In0_c0 <= "" & bh7_w80_12_c0 & bh7_w80_11_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid549_In1_c0 <= "" & bh7_w81_8_c0 & bh7_w81_11_c0;
   bh7_w80_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0(0);
   bh7_w81_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0(1);
   bh7_w82_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid549: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid549_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid549_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_copy550_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_copy550_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid551_In0_c0 <= "" & bh7_w82_12_c0 & bh7_w82_11_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid551_In1_c0 <= "" & bh7_w83_10_c0 & bh7_w83_11_c0;
   bh7_w82_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0(0);
   bh7_w83_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0(1);
   bh7_w84_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid551: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid551_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid551_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_copy552_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_copy552_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid553_In0_c0 <= "" & bh7_w84_10_c0 & bh7_w84_12_c0 & bh7_w84_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid553_In1_c0 <= "" & bh7_w85_12_c0 & bh7_w85_11_c0;
   bh7_w84_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0(0);
   bh7_w85_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0(1);
   bh7_w86_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid553: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid553_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid553_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_copy554_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_copy554_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid555_In0_c0 <= "" & bh7_w86_9_c0 & bh7_w86_10_c0 & "0";
   bh7_w86_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_c0(0);
   bh7_w87_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid555: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid555_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_copy556_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_copy556_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid557_In0_c0 <= "" & bh7_w87_10_c0 & bh7_w87_12_c0 & bh7_w87_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid557_In1_c0 <= "" & bh7_w88_12_c0 & bh7_w88_11_c0;
   bh7_w87_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0(0);
   bh7_w88_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0(1);
   bh7_w89_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid557: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid557_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid557_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_copy558_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_copy558_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid559_In0_c0 <= "" & bh7_w89_9_c0 & bh7_w89_10_c0 & "0";
   bh7_w89_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_c0(0);
   bh7_w90_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid559: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid559_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_copy560_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_copy560_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid561_In0_c0 <= "" & bh7_w90_10_c0 & bh7_w90_12_c0 & bh7_w90_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid561_In1_c0 <= "" & bh7_w91_12_c0 & bh7_w91_11_c0;
   bh7_w90_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0(0);
   bh7_w91_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0(1);
   bh7_w92_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid561: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid561_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid561_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_copy562_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_copy562_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid563_In0_c0 <= "" & bh7_w92_9_c0 & bh7_w92_10_c0 & "0";
   bh7_w92_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_c0(0);
   bh7_w93_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid563: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid563_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_copy564_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_copy564_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid565_In0_c0 <= "" & bh7_w93_10_c0 & bh7_w93_12_c0 & bh7_w93_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid565_In1_c0 <= "" & bh7_w94_12_c0 & bh7_w94_11_c0;
   bh7_w93_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0(0);
   bh7_w94_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0(1);
   bh7_w95_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid565: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid565_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid565_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_copy566_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_copy566_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid567_In0_c0 <= "" & bh7_w95_9_c0 & bh7_w95_10_c0 & "0";
   bh7_w95_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_c0(0);
   bh7_w96_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid567: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid567_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_copy568_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_copy568_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid569_In0_c0 <= "" & bh7_w96_10_c0 & bh7_w96_12_c0 & bh7_w96_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid569_In1_c0 <= "" & bh7_w97_12_c0 & bh7_w97_11_c0;
   bh7_w96_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0(0);
   bh7_w97_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0(1);
   bh7_w98_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid569: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid569_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid569_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_copy570_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_copy570_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid571_In0_c0 <= "" & bh7_w98_9_c0 & bh7_w98_10_c0 & "0";
   bh7_w98_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_c0(0);
   bh7_w99_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid571: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid571_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_copy572_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_copy572_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid573_In0_c0 <= "" & bh7_w99_9_c0 & bh7_w99_11_c0 & bh7_w99_10_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid573_In1_c0 <= "" & bh7_w100_7_c0 & bh7_w100_9_c0;
   bh7_w99_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0(0);
   bh7_w100_10_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0(1);
   bh7_w101_8_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid573: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid573_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid573_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_copy574_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_copy574_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid575_In0_c0 <= "" & bh7_w101_7_c0 & bh7_w101_6_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid575_In1_c0 <= "" & bh7_w102_4_c0 & bh7_w102_7_c0;
   bh7_w101_9_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0(0);
   bh7_w102_8_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0(1);
   bh7_w103_5_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid575: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid575_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid575_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_copy576_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_copy576_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid577_In0_c0 <= "" & bh7_w103_4_c0 & bh7_w103_3_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid577_In1_c0 <= "" & bh7_w104_2_c0;
   bh7_w103_6_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0(0);
   bh7_w104_3_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0(1);
   bh7_w105_2_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid577: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid577_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid577_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_copy578_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_copy578_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid579_In0_c0 <= "" & bh7_w105_0_c0 & bh7_w105_1_c0 & "0";
   bh7_w105_3_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_c0(0);
   Compressor_3_2_Freq300_uid432_uid579: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid579_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_copy580_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_copy580_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid581_In0_c0 <= "" & bh7_w55_16_c0 & bh7_w55_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid581_In1_c0 <= "" & bh7_w56_14_c0;
   bh7_w55_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0(0);
   bh7_w56_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0(1);
   bh7_w57_18_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid581: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid581_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid581_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_copy582_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_copy582_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid583_In0_c0 <= "" & bh7_w57_16_c0 & bh7_w57_17_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid583_In1_c0 <= "" & bh7_w58_16_c0 & bh7_w58_17_c0;
   bh7_w57_19_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0(0);
   bh7_w58_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0(1);
   bh7_w59_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid583: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid583_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid583_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_copy584_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_copy584_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid585_In0_c0 <= "" & bh7_w60_16_c0 & bh7_w60_17_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid585_In1_c0 <= "" & bh7_w61_16_c0 & bh7_w61_17_c0;
   bh7_w60_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0(0);
   bh7_w61_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0(1);
   bh7_w62_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid585: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid585_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid585_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_copy586_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_copy586_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid587_In0_c0 <= "" & bh7_w63_16_c0 & bh7_w63_17_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid587_In1_c0 <= "" & bh7_w64_16_c0 & bh7_w64_17_c0;
   bh7_w63_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0(0);
   bh7_w64_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0(1);
   bh7_w65_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid587: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid587_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid587_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_copy588_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_copy588_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid589_In0_c0 <= "" & bh7_w66_15_c0 & bh7_w66_16_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid589_In1_c0 <= "" & bh7_w67_14_c0;
   bh7_w66_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0(0);
   bh7_w67_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0(1);
   bh7_w68_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid589: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid589_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid589_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_copy590_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_copy590_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid591_In0_c0 <= "" & bh7_w68_15_c0 & bh7_w68_16_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid591_In1_c0 <= "" & bh7_w69_13_c0;
   bh7_w68_18_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0(0);
   bh7_w69_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0(1);
   bh7_w70_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid591: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid591_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid591_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_copy592_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_copy592_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid593_In0_c0 <= "" & bh7_w70_14_c0 & bh7_w70_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid593_In1_c0 <= "" & bh7_w71_13_c0;
   bh7_w70_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0(0);
   bh7_w71_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0(1);
   bh7_w72_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid593: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid593_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid593_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_copy594_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_copy594_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid595_In0_c0 <= "" & bh7_w72_15_c0 & bh7_w72_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid595_In1_c0 <= "" & bh7_w73_13_c0;
   bh7_w72_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0(0);
   bh7_w73_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0(1);
   bh7_w74_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid595: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid595_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid595_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_copy596_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_copy596_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid597_In0_c0 <= "" & bh7_w74_15_c0 & bh7_w74_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid597_In1_c0 <= "" & bh7_w75_12_c0;
   bh7_w74_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0(0);
   bh7_w75_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0(1);
   bh7_w76_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid597: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid597_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid597_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_copy598_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_copy598_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid599_In0_c0 <= "" & bh7_w76_14_c0 & bh7_w76_13_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid599_In1_c0 <= "" & bh7_w77_12_c0;
   bh7_w76_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0(0);
   bh7_w77_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0(1);
   bh7_w78_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid599: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid599_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid599_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_copy600_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_copy600_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid601_In0_c0 <= "" & bh7_w78_14_c0 & bh7_w78_13_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid601_In1_c0 <= "" & bh7_w79_12_c0;
   bh7_w78_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0(0);
   bh7_w79_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0(1);
   bh7_w80_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid601: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid601_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid601_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_copy602_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_copy602_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid603_In0_c0 <= "" & bh7_w80_14_c0 & bh7_w80_13_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid603_In1_c0 <= "" & bh7_w81_12_c0;
   bh7_w80_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0(0);
   bh7_w81_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0(1);
   bh7_w82_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid603: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid603_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid603_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_copy604_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_copy604_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid605_In0_c0 <= "" & bh7_w82_14_c0 & bh7_w82_13_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid605_In1_c0 <= "" & bh7_w83_12_c0;
   bh7_w82_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0(0);
   bh7_w83_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0(1);
   bh7_w84_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid605: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid605_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid605_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_copy606_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_copy606_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid607_In0_c0 <= "" & bh7_w84_13_c0 & bh7_w84_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid607_In1_c0 <= "" & bh7_w85_13_c0;
   bh7_w84_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0(0);
   bh7_w85_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0(1);
   bh7_w86_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid607: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid607_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid607_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_copy608_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_copy608_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid609_In0_c0 <= "" & bh7_w86_11_c0 & bh7_w86_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid609_In1_c0 <= "" & bh7_w87_13_c0 & bh7_w87_14_c0;
   bh7_w86_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0(0);
   bh7_w87_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0(1);
   bh7_w88_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid609: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid609_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid609_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_copy610_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_copy610_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid611_In0_c0 <= "" & bh7_w89_11_c0 & bh7_w89_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid611_In1_c0 <= "" & bh7_w90_13_c0 & bh7_w90_14_c0;
   bh7_w89_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0(0);
   bh7_w90_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0(1);
   bh7_w91_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid611: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid611_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid611_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_copy612_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_copy612_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid613_In0_c0 <= "" & bh7_w92_11_c0 & bh7_w92_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid613_In1_c0 <= "" & bh7_w93_13_c0 & bh7_w93_14_c0;
   bh7_w92_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0(0);
   bh7_w93_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0(1);
   bh7_w94_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid613: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid613_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid613_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_copy614_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_copy614_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid615_In0_c0 <= "" & bh7_w95_11_c0 & bh7_w95_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid615_In1_c0 <= "" & bh7_w96_13_c0 & bh7_w96_14_c0;
   bh7_w95_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0(0);
   bh7_w96_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0(1);
   bh7_w97_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid615: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid615_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid615_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_copy616_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_copy616_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid617_In0_c0 <= "" & bh7_w98_11_c0 & bh7_w98_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid617_In1_c0 <= "" & bh7_w99_12_c0 & bh7_w99_13_c0;
   bh7_w98_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0(0);
   bh7_w99_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0(1);
   bh7_w100_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid617: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid617_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid617_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_copy618_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_copy618_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid619_In0_c0 <= "" & bh7_w101_8_c0 & bh7_w101_9_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid619_In1_c0 <= "" & bh7_w102_8_c0;
   bh7_w101_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0(0);
   bh7_w102_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0(1);
   bh7_w103_7_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid619: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid619_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid619_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_copy620_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_copy620_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid621_In0_c0 <= "" & bh7_w103_6_c0 & bh7_w103_5_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid621_In1_c0 <= "" & bh7_w104_3_c0;
   bh7_w103_8_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0(0);
   bh7_w104_4_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0(1);
   bh7_w105_4_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid621: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid621_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid621_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_copy622_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_copy622_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid623_In0_c0 <= "" & bh7_w105_3_c0 & bh7_w105_2_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid623_In1_c0 <= "" & "0";
   bh7_w105_5_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_c0(0);
   Compressor_14_3_Freq300_uid326_uid623: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid623_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid623_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_copy624_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_copy624_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid625_In0_c0 <= "" & bh7_w57_18_c0 & bh7_w57_19_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid625_In1_c0 <= "" & bh7_w58_18_c0;
   bh7_w57_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1(0);
   bh7_w58_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1(1);
   bh7_w59_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid625: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid625_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid625_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid627_In0_c0 <= "" & bh7_w59_14_c0 & bh7_w59_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid627_In1_c0 <= "" & bh7_w60_18_c0;
   bh7_w59_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1(0);
   bh7_w60_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1(1);
   bh7_w61_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid627: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid627_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid627_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid629_In0_c0 <= "" & bh7_w62_14_c0 & bh7_w62_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid629_In1_c0 <= "" & bh7_w63_18_c0;
   bh7_w62_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1(0);
   bh7_w63_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1(1);
   bh7_w64_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid629: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid629_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid629_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid631_In0_c0 <= "" & bh7_w65_13_c0 & bh7_w65_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid631_In1_c0 <= "" & bh7_w66_17_c0;
   bh7_w65_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1(0);
   bh7_w66_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1(1);
   bh7_w67_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid631: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid631_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid631_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid633_In0_c0 <= "" & bh7_w68_17_c0 & bh7_w68_18_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid633_In1_c0 <= "" & bh7_w69_14_c0;
   bh7_w68_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1(0);
   bh7_w69_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1(1);
   bh7_w70_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid633: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid633_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid633_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid635_In0_c0 <= "" & bh7_w70_16_c0 & bh7_w70_17_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid635_In1_c0 <= "" & bh7_w71_14_c0;
   bh7_w70_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1(0);
   bh7_w71_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1(1);
   bh7_w72_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid635: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid635_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid635_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid637_In0_c0 <= "" & bh7_w72_16_c0 & bh7_w72_17_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid637_In1_c0 <= "" & bh7_w73_14_c0;
   bh7_w72_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1(0);
   bh7_w73_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1(1);
   bh7_w74_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid637: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid637_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid637_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid639_In0_c0 <= "" & bh7_w74_17_c0 & bh7_w74_16_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid639_In1_c0 <= "" & bh7_w75_13_c0;
   bh7_w74_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1(0);
   bh7_w75_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1(1);
   bh7_w76_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid639: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid639_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid639_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid641_In0_c0 <= "" & bh7_w76_16_c0 & bh7_w76_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid641_In1_c0 <= "" & bh7_w77_13_c0;
   bh7_w76_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1(0);
   bh7_w77_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1(1);
   bh7_w78_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid641: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid641_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid641_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid643_In0_c0 <= "" & bh7_w78_16_c0 & bh7_w78_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid643_In1_c0 <= "" & bh7_w79_13_c0;
   bh7_w78_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1(0);
   bh7_w79_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1(1);
   bh7_w80_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid643: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid643_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid643_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid645_In0_c0 <= "" & bh7_w80_16_c0 & bh7_w80_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid645_In1_c0 <= "" & bh7_w81_13_c0;
   bh7_w80_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1(0);
   bh7_w81_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1(1);
   bh7_w82_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid645: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid645_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid645_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid647_In0_c0 <= "" & bh7_w82_16_c0 & bh7_w82_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid647_In1_c0 <= "" & bh7_w83_13_c0;
   bh7_w82_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1(0);
   bh7_w83_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1(1);
   bh7_w84_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid647: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid647_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid647_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid649_In0_c0 <= "" & bh7_w84_15_c0 & bh7_w84_16_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid649_In1_c0 <= "" & bh7_w85_14_c0;
   bh7_w84_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1(0);
   bh7_w85_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1(1);
   bh7_w86_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid649: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid649_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid649_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid651_In0_c0 <= "" & bh7_w86_13_c0 & bh7_w86_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid651_In1_c0 <= "" & bh7_w87_15_c0;
   bh7_w86_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1(0);
   bh7_w87_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1(1);
   bh7_w88_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid651: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid651_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid651_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid653_In0_c0 <= "" & bh7_w88_13_c0 & bh7_w88_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid653_In1_c0 <= "" & bh7_w89_13_c0;
   bh7_w88_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1(0);
   bh7_w89_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1(1);
   bh7_w90_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid653: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid653_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid653_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid655_In0_c0 <= "" & bh7_w91_13_c0 & bh7_w91_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid655_In1_c0 <= "" & bh7_w92_13_c0;
   bh7_w91_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1(0);
   bh7_w92_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1(1);
   bh7_w93_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid655: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid655_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid655_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid657_In0_c0 <= "" & bh7_w94_13_c0 & bh7_w94_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid657_In1_c0 <= "" & bh7_w95_13_c0;
   bh7_w94_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1(0);
   bh7_w95_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1(1);
   bh7_w96_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid657: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid657_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid657_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid659_In0_c0 <= "" & bh7_w97_13_c0 & bh7_w97_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid659_In1_c0 <= "" & bh7_w98_13_c0;
   bh7_w97_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1(0);
   bh7_w98_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1(1);
   bh7_w99_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid659: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid659_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid659_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid661_In0_c0 <= "" & bh7_w100_10_c0 & bh7_w100_11_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid661_In1_c0 <= "" & bh7_w101_10_c0;
   bh7_w100_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1(0);
   bh7_w101_11_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1(1);
   bh7_w102_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid661: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid661_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid661_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid663_In0_c0 <= "" & bh7_w103_7_c0 & bh7_w103_8_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid663_In1_c0 <= "" & bh7_w104_4_c0;
   bh7_w103_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1(0);
   bh7_w104_5_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1(1);
   bh7_w105_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid663: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid663_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid663_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid665_In0_c0 <= "" & bh7_w105_5_c0 & bh7_w105_4_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid665_In1_c0 <= "" & "0";
   bh7_w105_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_c1(0);
   Compressor_14_3_Freq300_uid326_uid665: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid665_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid665_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid667_In0_c0 <= "" & bh7_w17_0_c0 & bh7_w17_1_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid667_In1_c0 <= "" & bh7_w18_0_c0 & bh7_w18_1_c0;
   bh7_w17_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1(0);
   bh7_w18_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1(1);
   bh7_w19_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid667: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid667_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid667_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid669_In0_c0 <= "" & bh7_w19_0_c0 & bh7_w19_1_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid669_In1_c0 <= "" & bh7_w20_0_c0 & bh7_w20_1_c0;
   bh7_w19_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1(0);
   bh7_w20_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1(1);
   bh7_w21_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid669: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid669_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid669_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid671_In0_c0 <= "" & bh7_w21_0_c0 & bh7_w21_1_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid671_In1_c0 <= "" & bh7_w22_0_c0 & bh7_w22_1_c0;
   bh7_w21_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1(0);
   bh7_w22_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1(1);
   bh7_w23_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid671: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid671_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid671_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid673_In0_c0 <= "" & bh7_w23_0_c0 & bh7_w23_1_c0 & "0";
   bh7_w23_3_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_c1(0);
   bh7_w24_3_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid673: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid673_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid675_In0_c0 <= "" & bh7_w24_0_c0 & bh7_w24_1_c0 & bh7_w24_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid675_In1_c0 <= "" & bh7_w25_0_c0 & bh7_w25_1_c0;
   bh7_w24_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1(0);
   bh7_w25_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1(1);
   bh7_w26_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid675: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid675_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid675_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid677_In0_c0 <= "" & bh7_w26_0_c0 & bh7_w26_1_c0 & bh7_w26_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid677_In1_c0 <= "" & bh7_w27_0_c0 & bh7_w27_1_c0;
   bh7_w26_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1(0);
   bh7_w27_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1(1);
   bh7_w28_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid677: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid677_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid677_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid679_In0_c0 <= "" & bh7_w28_0_c0 & bh7_w28_1_c0 & bh7_w28_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid679_In1_c0 <= "" & bh7_w29_0_c0 & bh7_w29_1_c0;
   bh7_w28_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1(0);
   bh7_w29_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1(1);
   bh7_w30_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid679: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid679_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid679_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid681_In0_c0 <= "" & bh7_w30_0_c0 & bh7_w30_1_c0 & bh7_w30_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid681_In1_c0 <= "" & bh7_w31_0_c0 & bh7_w31_1_c0;
   bh7_w30_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1(0);
   bh7_w31_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1(1);
   bh7_w32_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid681: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid681_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid681_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid683_In0_c0 <= "" & bh7_w32_0_c0 & bh7_w32_1_c0 & bh7_w32_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid683_In1_c0 <= "" & bh7_w33_0_c0 & bh7_w33_1_c0;
   bh7_w32_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1(0);
   bh7_w33_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1(1);
   bh7_w34_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid683: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid683_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid683_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid685_In0_c0 <= "" & bh7_w34_0_c0 & bh7_w34_1_c0 & bh7_w34_2_c0 & bh7_w34_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid685_In1_c0 <= "" & bh7_w35_0_c0;
   bh7_w34_5_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1(0);
   bh7_w35_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1(1);
   bh7_w36_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid685: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid685_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid685_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid687_In0_c0 <= "" & bh7_w35_1_c0 & bh7_w35_2_c0 & bh7_w35_3_c0;
   bh7_w35_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_c1(0);
   bh7_w36_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid687: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid687_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid689_In0_c0 <= "" & bh7_w36_0_c0 & bh7_w36_1_c0 & bh7_w36_2_c0 & bh7_w36_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid689_In1_c0 <= "" & bh7_w37_0_c0;
   bh7_w36_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1(0);
   bh7_w37_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1(1);
   bh7_w38_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid689: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid689_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid689_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid691_In0_c0 <= "" & bh7_w37_1_c0 & bh7_w37_2_c0 & bh7_w37_3_c0;
   bh7_w37_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_c1(0);
   bh7_w38_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid691: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid691_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid693_In0_c0 <= "" & bh7_w38_0_c0 & bh7_w38_1_c0 & bh7_w38_2_c0 & bh7_w38_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid693_In1_c0 <= "" & bh7_w39_0_c0;
   bh7_w38_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1(0);
   bh7_w39_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1(1);
   bh7_w40_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid693: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid693_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid693_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid695_In0_c0 <= "" & bh7_w39_1_c0 & bh7_w39_2_c0 & bh7_w39_3_c0;
   bh7_w39_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_c1(0);
   bh7_w40_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid695: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid695_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid697_In0_c0 <= "" & bh7_w40_0_c0 & bh7_w40_1_c0 & bh7_w40_2_c0 & bh7_w40_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid697_In1_c0 <= "" & bh7_w41_0_c0;
   bh7_w40_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1(0);
   bh7_w41_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1(1);
   bh7_w42_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid697: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid697_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid697_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid699_In0_c0 <= "" & bh7_w41_1_c0 & bh7_w41_2_c0 & bh7_w41_3_c0;
   bh7_w41_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_c1(0);
   bh7_w42_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid699: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid699_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid701_In0_c0 <= "" & bh7_w42_0_c0 & bh7_w42_1_c0 & bh7_w42_2_c0 & bh7_w42_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid701_In1_c0 <= "" & bh7_w43_0_c0;
   bh7_w42_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1(0);
   bh7_w43_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1(1);
   bh7_w44_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid701: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid701_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid701_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid703_In0_c0 <= "" & bh7_w43_1_c0 & bh7_w43_2_c0 & bh7_w43_3_c0;
   bh7_w43_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_c1(0);
   bh7_w44_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid703: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid703_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid705_In0_c0 <= "" & bh7_w44_0_c0 & bh7_w44_1_c0 & bh7_w44_2_c0 & bh7_w44_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid705_In1_c0 <= "" & bh7_w45_0_c0;
   bh7_w44_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1(0);
   bh7_w45_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1(1);
   bh7_w46_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid705: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid705_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid705_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid707_In0_c0 <= "" & bh7_w45_1_c0 & bh7_w45_2_c0 & bh7_w45_3_c0;
   bh7_w45_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_c1(0);
   bh7_w46_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid707: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid707_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid709_In0_c0 <= "" & bh7_w46_0_c0 & bh7_w46_1_c0 & bh7_w46_2_c0 & bh7_w46_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid709_In1_c0 <= "" & bh7_w47_0_c0;
   bh7_w46_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1(0);
   bh7_w47_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1(1);
   bh7_w48_5_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid709: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid709_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid709_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid711_In0_c0 <= "" & bh7_w47_1_c0 & bh7_w47_2_c0 & bh7_w47_3_c0;
   bh7_w47_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_c1(0);
   bh7_w48_6_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid711: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid711_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid713_In0_c0 <= "" & bh7_w48_4_c0 & bh7_w48_0_c0 & bh7_w48_1_c0 & bh7_w48_2_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid713_In1_c0 <= "" & bh7_w49_5_c0;
   bh7_w48_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1(0);
   bh7_w49_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1(1);
   bh7_w50_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid713: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid713_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid713_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid715_In0_c0 <= "" & bh7_w49_0_c0 & bh7_w49_1_c0 & bh7_w49_2_c0 & bh7_w49_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid715_In1_c0 <= "" & bh7_w50_6_c0;
   bh7_w49_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1(0);
   bh7_w50_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1(1);
   bh7_w51_11_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid715: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid715_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid715_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid717_In0_c0 <= "" & bh7_w50_0_c0 & bh7_w50_1_c0 & bh7_w50_2_c0 & bh7_w50_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid717_In1_c0 <= "" & bh7_w51_10_c0;
   bh7_w50_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1(0);
   bh7_w51_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1(1);
   bh7_w52_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid717: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid717_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid717_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid719_In0_c0 <= "" & bh7_w51_0_c0 & bh7_w51_1_c0 & bh7_w51_3_c0 & bh7_w51_4_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid719_In1_c0 <= "" & bh7_w52_11_c0;
   bh7_w51_13_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1(0);
   bh7_w52_13_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1(1);
   bh7_w53_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid719: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid719_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid719_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid721_In0_c0 <= "" & bh7_w52_0_c0 & bh7_w52_1_c0 & bh7_w52_3_c0 & bh7_w52_4_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid721_In1_c0 <= "" & bh7_w53_14_c0;
   bh7_w52_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1(0);
   bh7_w53_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1(1);
   bh7_w54_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid721: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid721_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid721_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid723_In0_c0 <= "" & bh7_w53_0_c0 & bh7_w53_1_c0 & bh7_w53_3_c0 & bh7_w53_4_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid723_In1_c0 <= "" & bh7_w54_15_c0;
   bh7_w53_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1(0);
   bh7_w54_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1(1);
   bh7_w55_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid723: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid723_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid723_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid725_In0_c0 <= "" & bh7_w54_0_c0 & bh7_w54_1_c0 & bh7_w54_4_c0 & bh7_w54_5_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid725_In1_c0 <= "" & bh7_w55_17_c0;
   bh7_w54_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1(0);
   bh7_w55_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1(1);
   bh7_w56_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid725: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid725_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid725_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid727_In0_c0 <= "" & bh7_w55_0_c0 & bh7_w55_1_c0 & bh7_w55_4_c0 & bh7_w55_5_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid727_In1_c0 <= "" & bh7_w56_15_c0;
   bh7_w55_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1(0);
   bh7_w56_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1(1);
   bh7_w57_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid727: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid727_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid727_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c0 <= "" & bh7_w56_0_c0 & bh7_w56_1_c0 & bh7_w56_3_c0 & bh7_w56_4_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid729_In1_c1 <= "" & bh7_w57_20_c1;
   bh7_w56_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1(0);
   bh7_w57_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1(1);
   bh7_w58_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid729: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid729_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_copy730_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_copy730_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c0 <= "" & bh7_w57_0_c0 & bh7_w57_1_c0 & bh7_w57_4_c0 & bh7_w57_5_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid731_In1_c1 <= "" & bh7_w58_19_c1;
   bh7_w57_23_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1(0);
   bh7_w58_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1(1);
   bh7_w59_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid731: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid731_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_copy732_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_copy732_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid733_In0_c0 <= "" & bh7_w58_0_c0 & bh7_w58_3_c0 & bh7_w58_4_c0;
   bh7_w58_22_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_c1(0);
   bh7_w59_19_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid733: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid733_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid735_In0_c1 <= "" & bh7_w59_16_c1 & bh7_w59_17_c1 & bh7_w59_0_c1 & bh7_w59_2_c1 & bh7_w59_3_c1 & bh7_w59_4_c1;
   bh7_w59_20_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1(0);
   bh7_w60_20_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1(1);
   bh7_w61_20_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1(2);
   Compressor_6_3_Freq300_uid334_uid735: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid735_In0_c1,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_copy736_c1);
   Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_copy736_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid737_In0_c1 <= "" & bh7_w60_19_c1 & bh7_w60_0_c1 & bh7_w60_3_c1 & bh7_w60_4_c1 & bh7_w60_5_c1;
   bh7_w60_21_c1 <= Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1(0);
   bh7_w61_21_c1 <= Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1(1);
   bh7_w62_17_c1 <= Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1(2);
   Compressor_5_3_Freq300_uid400_uid737: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid737_In0_c1,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_copy738_c1);
   Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1 <= Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_copy738_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid739_In0_c1 <= "" & bh7_w61_18_c1 & bh7_w61_19_c1 & bh7_w61_0_c1 & bh7_w61_3_c1 & bh7_w61_4_c1 & bh7_w61_5_c1;
   bh7_w61_22_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1(0);
   bh7_w62_18_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1(1);
   bh7_w63_20_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1(2);
   Compressor_6_3_Freq300_uid334_uid739: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid739_In0_c1,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_copy740_c1);
   Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_copy740_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid741_In0_c1 <= "" & bh7_w62_16_c1 & bh7_w62_0_c1 & bh7_w62_2_c1 & bh7_w62_3_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid741_In1_c1 <= "" & bh7_w63_19_c1;
   bh7_w62_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1(0);
   bh7_w63_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1(1);
   bh7_w64_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid741: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid741_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid741_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_copy742_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_copy742_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid743_In0_c0 <= "" & bh7_w63_0_c0 & bh7_w63_3_c0 & bh7_w63_4_c0;
   bh7_w63_22_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_c1(0);
   bh7_w64_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid743: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid743_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid745_In0_c1 <= "" & bh7_w64_18_c1 & bh7_w64_19_c1 & bh7_w64_0_c1 & bh7_w64_3_c1 & bh7_w64_4_c1 & bh7_w64_5_c1;
   bh7_w64_22_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1(0);
   bh7_w65_16_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1(1);
   bh7_w66_19_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1(2);
   Compressor_6_3_Freq300_uid334_uid745: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid745_In0_c1,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_copy746_c1);
   Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_copy746_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid747_In0_c1 <= "" & bh7_w65_15_c1 & bh7_w65_0_c1 & bh7_w65_2_c1 & bh7_w65_3_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid747_In1_c1 <= "" & bh7_w66_18_c1;
   bh7_w65_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1(0);
   bh7_w66_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1(1);
   bh7_w67_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid747: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid747_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid747_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_copy748_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_copy748_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid749_In0_c0 <= "" & bh7_w66_0_c0 & bh7_w66_3_c0 & bh7_w66_4_c0;
   bh7_w66_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_c1(0);
   bh7_w67_18_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid749: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid749_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid751_In0_c1 <= "" & bh7_w67_15_c1 & bh7_w67_16_c1 & bh7_w67_0_c1 & bh7_w67_3_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid751_In1_c1 <= "" & bh7_w68_19_c1;
   bh7_w67_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1(0);
   bh7_w68_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1(1);
   bh7_w69_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid751: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid751_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid751_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_copy752_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_copy752_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid753_In0_c0 <= "" & bh7_w68_0_c0 & bh7_w68_2_c0 & bh7_w68_3_c0;
   bh7_w68_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_c1(0);
   bh7_w69_17_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid753: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid753_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid755_In0_c1 <= "" & bh7_w69_15_c1 & bh7_w69_0_c1 & bh7_w69_3_c1 & bh7_w69_4_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid755_In1_c1 <= "" & bh7_w70_18_c1;
   bh7_w69_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1(0);
   bh7_w70_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1(1);
   bh7_w71_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid755: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid755_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid755_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_copy756_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_copy756_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid757_In0_c1 <= "" & bh7_w70_19_c1 & bh7_w70_0_c1 & bh7_w70_3_c1 & bh7_w70_4_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid757_In1_c1 <= "" & bh7_w71_15_c1;
   bh7_w70_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1(0);
   bh7_w71_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1(1);
   bh7_w72_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid757: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid757_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid757_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_copy758_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_copy758_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid759_In0_c0 <= "" & bh7_w71_0_c0 & bh7_w71_2_c0 & bh7_w71_3_c0;
   bh7_w71_18_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_c1(0);
   bh7_w72_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid759: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid759_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid761_In0_c1 <= "" & bh7_w72_18_c1 & bh7_w72_19_c1 & bh7_w72_0_c1 & bh7_w72_3_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid761_In1_c1 <= "" & bh7_w73_15_c1;
   bh7_w72_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1(0);
   bh7_w73_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1(1);
   bh7_w74_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid761: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid761_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid761_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_copy762_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_copy762_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid763_In0_c0 <= "" & bh7_w73_0_c0 & bh7_w73_3_c0 & bh7_w73_4_c0;
   bh7_w73_17_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_c1(0);
   bh7_w74_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid763: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid763_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid765_In0_c1 <= "" & bh7_w74_18_c1 & bh7_w74_0_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c0 <= "" & bh7_w75_1_c0;
   bh7_w74_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1(0);
   bh7_w75_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1(1);
   bh7_w76_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid765: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid765_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_copy766_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_copy766_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid767_In0_c1 <= "" & bh7_w74_2_c1 & bh7_w74_3_c1 & bh7_w74_19_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid767_In1_c1 <= "" & bh7_w75_2_c1 & bh7_w75_14_c1;
   bh7_w74_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1(0);
   bh7_w75_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1(1);
   bh7_w76_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid767: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid767_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid767_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_copy768_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_copy768_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid769_In0_c1 <= "" & bh7_w76_1_c1 & bh7_w76_2_c1 & bh7_w76_18_c1 & bh7_w76_17_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c0 <= "" & "0";
   bh7_w76_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1(0);
   bh7_w77_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1(1);
   bh7_w78_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid769: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid769_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_copy770_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_copy770_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid771_In0_c1 <= "" & bh7_w77_0_c1 & bh7_w77_1_c1 & bh7_w77_14_c1;
   bh7_w77_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_c1(0);
   bh7_w78_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid771: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid771_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_copy772_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_copy772_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid773_In0_c1 <= "" & bh7_w78_0_c1 & bh7_w78_1_c1 & bh7_w78_18_c1 & bh7_w78_17_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c0 <= "" & "0";
   bh7_w78_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1(0);
   bh7_w79_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1(1);
   bh7_w80_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid773: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid773_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_copy774_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_copy774_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid775_In0_c1 <= "" & bh7_w79_0_c1 & bh7_w79_1_c1 & bh7_w79_14_c1;
   bh7_w79_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_c1(0);
   bh7_w80_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid775: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid775_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_copy776_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_copy776_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid777_In0_c1 <= "" & bh7_w80_0_c1 & bh7_w80_1_c1 & bh7_w80_18_c1 & bh7_w80_17_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c0 <= "" & "0";
   bh7_w80_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1(0);
   bh7_w81_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1(1);
   bh7_w82_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid777: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid777_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_copy778_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_copy778_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid779_In0_c1 <= "" & bh7_w81_0_c1 & bh7_w81_1_c1 & bh7_w81_14_c1;
   bh7_w81_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_c1(0);
   bh7_w82_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid779: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid779_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_copy780_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_copy780_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid781_In0_c1 <= "" & bh7_w82_18_c1 & bh7_w82_0_c1 & bh7_w82_17_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid781_In1_c1 <= "" & bh7_w83_14_c1 & bh7_w83_0_c1;
   bh7_w82_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1(0);
   bh7_w83_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1(1);
   bh7_w84_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid781: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid781_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid781_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_copy782_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_copy782_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid783_In0_c1 <= "" & bh7_w84_17_c1 & bh7_w84_18_c1 & bh7_w84_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid783_In1_c1 <= "" & bh7_w85_15_c1 & bh7_w85_0_c1;
   bh7_w84_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1(0);
   bh7_w85_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1(1);
   bh7_w86_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid783: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid783_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid783_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_copy784_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_copy784_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid785_In0_c1 <= "" & bh7_w86_15_c1 & bh7_w86_16_c1 & bh7_w86_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid785_In1_c1 <= "" & bh7_w87_16_c1 & bh7_w87_0_c1;
   bh7_w86_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1(0);
   bh7_w87_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1(1);
   bh7_w88_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid785: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid785_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid785_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_copy786_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_copy786_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid787_In0_c1 <= "" & bh7_w88_15_c1 & bh7_w88_16_c1 & bh7_w88_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid787_In1_c1 <= "" & bh7_w89_14_c1 & bh7_w89_0_c1;
   bh7_w88_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1(0);
   bh7_w89_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1(1);
   bh7_w90_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid787: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid787_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid787_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_copy788_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_copy788_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid789_In0_c1 <= "" & bh7_w90_15_c1 & bh7_w90_16_c1 & bh7_w90_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid789_In1_c1 <= "" & bh7_w91_15_c1 & bh7_w91_0_c1;
   bh7_w90_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1(0);
   bh7_w91_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1(1);
   bh7_w92_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid789: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid789_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid789_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_copy790_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_copy790_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid791_In0_c1 <= "" & bh7_w92_14_c1 & bh7_w92_0_c1 & "0";
   bh7_w92_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_c1(0);
   bh7_w93_17_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid791: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid791_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_copy792_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_copy792_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid793_In0_c1 <= "" & bh7_w93_15_c1 & bh7_w93_16_c1 & bh7_w93_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid793_In1_c1 <= "" & bh7_w94_15_c1 & bh7_w94_0_c1;
   bh7_w93_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1(0);
   bh7_w94_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1(1);
   bh7_w95_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid793: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid793_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid793_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_copy794_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_copy794_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid795_In0_c1 <= "" & bh7_w95_14_c1 & bh7_w95_0_c1 & "0";
   bh7_w95_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_c1(0);
   bh7_w96_17_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid795: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid795_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_copy796_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_copy796_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid797_In0_c1 <= "" & bh7_w96_15_c1 & bh7_w96_16_c1 & bh7_w96_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid797_In1_c1 <= "" & bh7_w97_15_c1 & bh7_w97_0_c1;
   bh7_w96_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1(0);
   bh7_w97_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1(1);
   bh7_w98_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid797: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid797_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid797_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_copy798_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_copy798_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid799_In0_c1 <= "" & bh7_w98_14_c1 & bh7_w98_0_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid799_In1_c1 <= "" & bh7_w99_14_c1 & bh7_w99_15_c1;
   bh7_w98_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1(0);
   bh7_w99_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1(1);
   bh7_w100_13_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid799: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid799_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid799_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_copy800_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_copy800_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid801_In0_c1 <= "" & bh7_w102_9_c1 & bh7_w102_10_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid801_In1_c1 <= "" & bh7_w103_9_c1;
   bh7_w102_11_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1(0);
   bh7_w103_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1(1);
   bh7_w104_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid801: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid801_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid801_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_copy802_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_copy802_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid803_In0_c1 <= "" & bh7_w105_6_c1 & bh7_w105_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c0 <= "" & "0";
   bh7_w105_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_c1(0);
   Compressor_14_3_Freq300_uid326_uid803: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid803_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_copy804_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_copy804_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid805_In0_c1 <= "" & bh7_w19_3_c1 & bh7_w19_2_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid805_In1_c1 <= "" & bh7_w20_2_c1;
   bh7_w19_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1(0);
   bh7_w20_3_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1(1);
   bh7_w21_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid805: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid805_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid805_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_copy806_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_copy806_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid807_In0_c1 <= "" & bh7_w21_3_c1 & bh7_w21_2_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid807_In1_c1 <= "" & bh7_w22_2_c1;
   bh7_w21_5_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1(0);
   bh7_w22_3_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1(1);
   bh7_w23_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid807: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid807_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid807_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_copy808_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_copy808_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid809_In0_c1 <= "" & bh7_w23_3_c1 & bh7_w23_2_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid809_In1_c1 <= "" & bh7_w24_4_c1 & bh7_w24_3_c1;
   bh7_w23_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1(0);
   bh7_w24_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1(1);
   bh7_w25_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid809: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid809_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid809_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_copy810_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_copy810_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid811_In0_c1 <= "" & bh7_w25_2_c1 & bh7_w25_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid811_In1_c1 <= "" & bh7_w26_4_c1 & bh7_w26_3_c1;
   bh7_w25_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1(0);
   bh7_w26_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1(1);
   bh7_w27_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid811: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid811_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid811_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_copy812_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_copy812_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid813_In0_c1 <= "" & bh7_w27_2_c1 & bh7_w27_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid813_In1_c1 <= "" & bh7_w28_4_c1 & bh7_w28_3_c1;
   bh7_w27_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1(0);
   bh7_w28_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1(1);
   bh7_w29_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid813: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid813_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid813_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_copy814_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_copy814_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid815_In0_c1 <= "" & bh7_w29_2_c1 & bh7_w29_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid815_In1_c1 <= "" & bh7_w30_4_c1 & bh7_w30_3_c1;
   bh7_w29_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1(0);
   bh7_w30_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1(1);
   bh7_w31_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid815: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid815_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid815_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_copy816_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_copy816_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid817_In0_c1 <= "" & bh7_w31_2_c1 & bh7_w31_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid817_In1_c1 <= "" & bh7_w32_4_c1 & bh7_w32_3_c1;
   bh7_w31_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1(0);
   bh7_w32_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1(1);
   bh7_w33_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid817: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid817_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid817_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_copy818_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_copy818_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid819_In0_c1 <= "" & bh7_w33_2_c1 & bh7_w33_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid819_In1_c1 <= "" & bh7_w34_5_c1 & bh7_w34_4_c1;
   bh7_w33_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1(0);
   bh7_w34_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1(1);
   bh7_w35_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid819: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid819_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid819_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_copy820_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_copy820_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid821_In0_c1 <= "" & bh7_w35_5_c1 & bh7_w35_4_c1 & "0";
   bh7_w35_7_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_c1(0);
   bh7_w36_7_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid821: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid821_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_copy822_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_copy822_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid823_In0_c1 <= "" & bh7_w36_6_c1 & bh7_w36_5_c1 & bh7_w36_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid823_In1_c1 <= "" & bh7_w37_5_c1 & bh7_w37_4_c1;
   bh7_w36_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1(0);
   bh7_w37_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1(1);
   bh7_w38_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid823: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid823_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid823_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_copy824_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_copy824_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid825_In0_c1 <= "" & bh7_w38_6_c1 & bh7_w38_5_c1 & bh7_w38_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid825_In1_c1 <= "" & bh7_w39_5_c1 & bh7_w39_4_c1;
   bh7_w38_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1(0);
   bh7_w39_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1(1);
   bh7_w40_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid825: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid825_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid825_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_copy826_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_copy826_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid827_In0_c1 <= "" & bh7_w40_6_c1 & bh7_w40_5_c1 & bh7_w40_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid827_In1_c1 <= "" & bh7_w41_5_c1 & bh7_w41_4_c1;
   bh7_w40_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1(0);
   bh7_w41_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1(1);
   bh7_w42_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid827: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid827_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid827_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_copy828_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_copy828_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid829_In0_c1 <= "" & bh7_w42_6_c1 & bh7_w42_5_c1 & bh7_w42_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid829_In1_c1 <= "" & bh7_w43_5_c1 & bh7_w43_4_c1;
   bh7_w42_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1(0);
   bh7_w43_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1(1);
   bh7_w44_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid829: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid829_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid829_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_copy830_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_copy830_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid831_In0_c1 <= "" & bh7_w44_6_c1 & bh7_w44_5_c1 & bh7_w44_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid831_In1_c1 <= "" & bh7_w45_5_c1 & bh7_w45_4_c1;
   bh7_w44_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1(0);
   bh7_w45_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1(1);
   bh7_w46_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid831: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid831_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid831_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_copy832_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_copy832_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid833_In0_c1 <= "" & bh7_w46_6_c1 & bh7_w46_5_c1 & bh7_w46_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid833_In1_c1 <= "" & bh7_w47_5_c1 & bh7_w47_4_c1;
   bh7_w46_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1(0);
   bh7_w47_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1(1);
   bh7_w48_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid833: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid833_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid833_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_copy834_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_copy834_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid835_In0_c1 <= "" & bh7_w48_3_c1 & bh7_w48_7_c1 & bh7_w48_6_c1 & bh7_w48_5_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid835_In1_c1 <= "" & bh7_w49_7_c1;
   bh7_w48_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1(0);
   bh7_w49_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1(1);
   bh7_w50_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid835: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid835_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid835_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_copy836_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_copy836_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid837_In0_c1 <= "" & bh7_w50_9_c1 & bh7_w50_8_c1 & bh7_w50_7_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid837_In1_c1 <= "" & bh7_w51_13_c1 & bh7_w51_12_c1;
   bh7_w50_11_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1(0);
   bh7_w51_14_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1(1);
   bh7_w52_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid837: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid837_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid837_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_copy838_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_copy838_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid839_In0_c1 <= "" & bh7_w52_14_c1 & bh7_w52_13_c1 & bh7_w52_12_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid839_In1_c1 <= "" & bh7_w53_17_c1 & bh7_w53_16_c1;
   bh7_w52_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1(0);
   bh7_w53_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1(1);
   bh7_w54_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid839: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid839_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid839_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_copy840_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_copy840_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid841_In0_c1 <= "" & bh7_w54_18_c1 & bh7_w54_17_c1 & bh7_w54_16_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid841_In1_c1 <= "" & bh7_w55_19_c1 & bh7_w55_20_c1;
   bh7_w54_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1(0);
   bh7_w55_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1(1);
   bh7_w56_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid841: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid841_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid841_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_copy842_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_copy842_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid843_In0_c1 <= "" & bh7_w56_16_c1 & bh7_w56_17_c1 & bh7_w56_18_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid843_In1_c1 <= "" & bh7_w57_21_c1 & bh7_w57_22_c1;
   bh7_w56_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1(0);
   bh7_w57_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1(1);
   bh7_w58_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid843: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid843_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid843_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_copy844_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_copy844_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid845_In0_c1 <= "" & bh7_w58_20_c1 & bh7_w58_21_c1 & bh7_w58_5_c1 & bh7_w58_22_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c0 <= "" & "0";
   bh7_w58_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1(0);
   bh7_w59_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1(1);
   bh7_w60_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid845: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid845_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_copy846_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_copy846_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid847_In0_c1 <= "" & bh7_w59_18_c1 & bh7_w59_20_c1 & bh7_w59_19_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid847_In1_c1 <= "" & bh7_w60_20_c1 & bh7_w60_21_c1;
   bh7_w59_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1(0);
   bh7_w60_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1(1);
   bh7_w61_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid847: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid847_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid847_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_copy848_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_copy848_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid849_In0_c1 <= "" & bh7_w61_20_c1 & bh7_w61_21_c1 & bh7_w61_22_c1;
   bh7_w61_24_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_c1(0);
   bh7_w62_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid849: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid849_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_copy850_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_copy850_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid851_In0_c1 <= "" & bh7_w62_17_c1 & bh7_w62_18_c1 & bh7_w62_19_c1 & bh7_w62_4_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid851_In1_c1 <= "" & bh7_w63_20_c1;
   bh7_w62_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1(0);
   bh7_w63_23_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1(1);
   bh7_w64_23_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid851: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid851_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid851_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_copy852_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_copy852_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid853_In0_c1 <= "" & bh7_w63_21_c1 & bh7_w63_5_c1 & bh7_w63_22_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c0 <= "" & "0" & "0";
   bh7_w63_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1(0);
   bh7_w64_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1(1);
   bh7_w65_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid853: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid853_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_copy854_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_copy854_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid855_In0_c1 <= "" & bh7_w64_20_c1 & bh7_w64_22_c1 & bh7_w64_21_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid855_In1_c1 <= "" & bh7_w65_16_c1 & bh7_w65_17_c1;
   bh7_w64_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1(0);
   bh7_w65_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1(1);
   bh7_w66_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid855: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid855_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid855_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_copy856_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_copy856_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid857_In0_c1 <= "" & bh7_w66_19_c1 & bh7_w66_20_c1 & bh7_w66_21_c1;
   bh7_w66_23_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_c1(0);
   bh7_w67_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid857: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid857_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_copy858_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_copy858_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid859_In0_c1 <= "" & bh7_w67_17_c1 & bh7_w67_19_c1 & bh7_w67_4_c1 & bh7_w67_18_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid859_In1_c1 <= "" & bh7_w68_20_c1;
   bh7_w67_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1(0);
   bh7_w68_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1(1);
   bh7_w69_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid859: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid859_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid859_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_copy860_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_copy860_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid861_In0_c1 <= "" & bh7_w69_16_c1 & bh7_w69_18_c1 & bh7_w69_17_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid861_In1_c1 <= "" & bh7_w70_20_c1 & bh7_w70_21_c1;
   bh7_w69_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1(0);
   bh7_w70_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1(1);
   bh7_w71_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid861: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid861_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid861_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_copy862_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_copy862_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid863_In0_c1 <= "" & bh7_w71_16_c1 & bh7_w71_17_c1 & bh7_w71_18_c1;
   bh7_w71_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_c1(0);
   bh7_w72_23_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid863: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid863_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_copy864_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_copy864_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid865_In0_c1 <= "" & bh7_w72_20_c1 & bh7_w72_22_c1 & bh7_w72_4_c1 & bh7_w72_21_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid865_In1_c1 <= "" & bh7_w73_16_c1;
   bh7_w72_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1(0);
   bh7_w73_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1(1);
   bh7_w74_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid865: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid865_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid865_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_copy866_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_copy866_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid867_In0_c1 <= "" & bh7_w74_20_c1 & bh7_w74_22_c1 & bh7_w74_21_c1 & bh7_w74_23_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid867_In1_c1 <= "" & bh7_w75_15_c1;
   bh7_w74_25_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1(0);
   bh7_w75_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1(1);
   bh7_w76_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid867: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid867_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid867_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_copy868_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_copy868_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid869_In0_c1 <= "" & bh7_w76_19_c1 & bh7_w76_21_c1 & bh7_w76_20_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid869_In1_c1 <= "" & bh7_w77_15_c1 & bh7_w77_16_c1;
   bh7_w76_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1(0);
   bh7_w77_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1(1);
   bh7_w78_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid869: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid869_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid869_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_copy870_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_copy870_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid871_In0_c1 <= "" & bh7_w78_19_c1 & bh7_w78_21_c1 & bh7_w78_20_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid871_In1_c1 <= "" & bh7_w79_15_c1 & bh7_w79_16_c1;
   bh7_w78_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1(0);
   bh7_w79_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1(1);
   bh7_w80_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid871: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid871_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid871_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_copy872_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_copy872_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid873_In0_c1 <= "" & bh7_w80_19_c1 & bh7_w80_21_c1 & bh7_w80_20_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid873_In1_c1 <= "" & bh7_w81_15_c1 & bh7_w81_16_c1;
   bh7_w80_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1(0);
   bh7_w81_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1(1);
   bh7_w82_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid873: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid873_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid873_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_copy874_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_copy874_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid875_In0_c1 <= "" & bh7_w82_19_c1 & bh7_w82_21_c1 & bh7_w82_20_c1;
   bh7_w82_23_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_c1(0);
   bh7_w83_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid875: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid875_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_copy876_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_copy876_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid877_In0_c1 <= "" & bh7_w84_19_c1 & bh7_w84_20_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid877_In1_c1 <= "" & bh7_w85_16_c1;
   bh7_w84_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1(0);
   bh7_w85_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1(1);
   bh7_w86_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid877: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid877_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid877_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_copy878_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_copy878_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid879_In0_c1 <= "" & bh7_w86_17_c1 & bh7_w86_18_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid879_In1_c1 <= "" & bh7_w87_17_c1;
   bh7_w86_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1(0);
   bh7_w87_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1(1);
   bh7_w88_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid879: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid879_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid879_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_copy880_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_copy880_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid881_In0_c1 <= "" & bh7_w88_17_c1 & bh7_w88_18_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid881_In1_c1 <= "" & bh7_w89_15_c1;
   bh7_w88_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1(0);
   bh7_w89_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1(1);
   bh7_w90_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid881: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid881_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid881_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_copy882_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_copy882_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid883_In0_c1 <= "" & bh7_w90_17_c1 & bh7_w90_18_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid883_In1_c1 <= "" & bh7_w91_16_c1;
   bh7_w90_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1(0);
   bh7_w91_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1(1);
   bh7_w92_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid883: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid883_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid883_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_copy884_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_copy884_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid885_In0_c1 <= "" & bh7_w92_15_c1 & bh7_w92_16_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid885_In1_c1 <= "" & bh7_w93_17_c1 & bh7_w93_18_c1;
   bh7_w92_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1(0);
   bh7_w93_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1(1);
   bh7_w94_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid885: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid885_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid885_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_copy886_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_copy886_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid887_In0_c1 <= "" & bh7_w95_15_c1 & bh7_w95_16_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid887_In1_c1 <= "" & bh7_w96_17_c1 & bh7_w96_18_c1;
   bh7_w95_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1(0);
   bh7_w96_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1(1);
   bh7_w97_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid887: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid887_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid887_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_copy888_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_copy888_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid889_In0_c1 <= "" & bh7_w98_15_c1 & bh7_w98_16_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid889_In1_c1 <= "" & bh7_w99_16_c1;
   bh7_w98_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1(0);
   bh7_w99_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1(1);
   bh7_w100_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid889: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid889_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid889_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_copy890_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_copy890_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid891_In0_c1 <= "" & bh7_w100_12_c1 & bh7_w100_13_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid891_In1_c1 <= "" & bh7_w101_11_c1;
   bh7_w100_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1(0);
   bh7_w101_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1(1);
   bh7_w102_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid891: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid891_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid891_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_copy892_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_copy892_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid893_In0_c1 <= "" & bh7_w104_5_c1 & bh7_w104_6_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid893_In1_c1 <= "" & bh7_w105_8_c1;
   bh7_w104_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_c1(0);
   bh7_w105_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_c1(1);
   Compressor_14_3_Freq300_uid326_uid893: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid893_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid893_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_copy894_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_copy894_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid895_In0_c1 <= "" & bh7_w21_5_c1 & bh7_w21_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid895_In1_c1 <= "" & bh7_w22_3_c1;
   bh7_w21_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1(0);
   bh7_w22_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1(1);
   bh7_w23_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid895: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid895_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid895_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_copy896_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_copy896_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid897_In0_c1 <= "" & bh7_w23_5_c1 & bh7_w23_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid897_In1_c1 <= "" & bh7_w24_5_c1;
   bh7_w23_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1(0);
   bh7_w24_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1(1);
   bh7_w25_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid897: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid897_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid897_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_copy898_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_copy898_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid899_In0_c1 <= "" & bh7_w25_5_c1 & bh7_w25_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid899_In1_c1 <= "" & bh7_w26_5_c1;
   bh7_w25_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1(0);
   bh7_w26_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1(1);
   bh7_w27_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid899: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid899_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid899_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_copy900_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_copy900_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid901_In0_c1 <= "" & bh7_w27_5_c1 & bh7_w27_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid901_In1_c1 <= "" & bh7_w28_5_c1;
   bh7_w27_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1(0);
   bh7_w28_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1(1);
   bh7_w29_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid901: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid901_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid901_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_copy902_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_copy902_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid903_In0_c1 <= "" & bh7_w29_5_c1 & bh7_w29_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid903_In1_c1 <= "" & bh7_w30_5_c1;
   bh7_w29_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1(0);
   bh7_w30_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1(1);
   bh7_w31_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid903: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid903_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid903_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_copy904_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_copy904_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid905_In0_c1 <= "" & bh7_w31_5_c1 & bh7_w31_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid905_In1_c1 <= "" & bh7_w32_5_c1;
   bh7_w31_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1(0);
   bh7_w32_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1(1);
   bh7_w33_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid905: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid905_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid905_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_copy906_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_copy906_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid907_In0_c1 <= "" & bh7_w33_5_c1 & bh7_w33_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid907_In1_c1 <= "" & bh7_w34_6_c1;
   bh7_w33_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1(0);
   bh7_w34_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1(1);
   bh7_w35_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid907: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid907_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid907_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_copy908_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_copy908_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid909_In0_c1 <= "" & bh7_w35_7_c1 & bh7_w35_6_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid909_In1_c1 <= "" & bh7_w36_8_c1 & bh7_w36_7_c1;
   bh7_w35_9_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1(0);
   bh7_w36_9_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1(1);
   bh7_w37_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid909: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid909_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid909_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_copy910_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_copy910_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid911_In0_c1 <= "" & bh7_w38_8_c1 & bh7_w38_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid911_In1_c1 <= "" & bh7_w39_6_c1;
   bh7_w38_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1(0);
   bh7_w39_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1(1);
   bh7_w40_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid911: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid911_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid911_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_copy912_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_copy912_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid913_In0_c1 <= "" & bh7_w40_8_c1 & bh7_w40_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid913_In1_c1 <= "" & bh7_w41_6_c1;
   bh7_w40_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1(0);
   bh7_w41_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1(1);
   bh7_w42_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid913: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid913_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid913_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_copy914_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_copy914_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid915_In0_c1 <= "" & bh7_w42_8_c1 & bh7_w42_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid915_In1_c1 <= "" & bh7_w43_6_c1;
   bh7_w42_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1(0);
   bh7_w43_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1(1);
   bh7_w44_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid915: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid915_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid915_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_copy916_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_copy916_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid917_In0_c1 <= "" & bh7_w44_8_c1 & bh7_w44_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid917_In1_c1 <= "" & bh7_w45_6_c1;
   bh7_w44_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1(0);
   bh7_w45_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1(1);
   bh7_w46_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid917: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid917_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid917_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_copy918_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_copy918_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid919_In0_c1 <= "" & bh7_w46_8_c1 & bh7_w46_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid919_In1_c1 <= "" & bh7_w47_6_c1;
   bh7_w46_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1(0);
   bh7_w47_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1(1);
   bh7_w48_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid919: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid919_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid919_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_copy920_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_copy920_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid921_In0_c1 <= "" & bh7_w48_9_c1 & bh7_w48_8_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid921_In1_c1 <= "" & bh7_w49_6_c1 & bh7_w49_8_c1;
   bh7_w48_11_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1(0);
   bh7_w49_9_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1(1);
   bh7_w50_12_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid921: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid921_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid921_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_copy922_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_copy922_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid923_In0_c1 <= "" & bh7_w50_11_c1 & bh7_w50_10_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid923_In1_c1 <= "" & bh7_w51_11_c1 & bh7_w51_14_c1;
   bh7_w50_13_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1(0);
   bh7_w51_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1(1);
   bh7_w52_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid923: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid923_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid923_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_copy924_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_copy924_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid925_In0_c1 <= "" & bh7_w52_16_c1 & bh7_w52_15_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid925_In1_c1 <= "" & bh7_w53_15_c1 & bh7_w53_18_c1;
   bh7_w52_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1(0);
   bh7_w53_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1(1);
   bh7_w54_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid925: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid925_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid925_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_copy926_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_copy926_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid927_In0_c1 <= "" & bh7_w54_20_c1 & bh7_w54_19_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid927_In1_c1 <= "" & bh7_w55_21_c1 & bh7_w55_18_c1;
   bh7_w54_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1(0);
   bh7_w55_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1(1);
   bh7_w56_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid927: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid927_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid927_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_copy928_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_copy928_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid929_In0_c1 <= "" & bh7_w56_19_c1 & bh7_w56_20_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid929_In1_c1 <= "" & bh7_w57_23_c1 & bh7_w57_24_c1;
   bh7_w56_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1(0);
   bh7_w57_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1(1);
   bh7_w58_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid929: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid929_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid929_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_copy930_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_copy930_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid931_In0_c1 <= "" & bh7_w58_23_c1 & bh7_w58_24_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid931_In1_c1 <= "" & bh7_w59_21_c1 & bh7_w59_22_c1;
   bh7_w58_26_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1(0);
   bh7_w59_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1(1);
   bh7_w60_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid931: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid931_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid931_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_copy932_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_copy932_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid933_In0_c1 <= "" & bh7_w60_22_c1 & bh7_w60_23_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid933_In1_c1 <= "" & bh7_w61_23_c1 & bh7_w61_24_c1;
   bh7_w60_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1(0);
   bh7_w61_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1(1);
   bh7_w62_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid933: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid933_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid933_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_copy934_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_copy934_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid935_In0_c1 <= "" & bh7_w62_20_c1 & bh7_w62_21_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid935_In1_c1 <= "" & bh7_w63_23_c1 & bh7_w63_24_c1;
   bh7_w62_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1(0);
   bh7_w63_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1(1);
   bh7_w64_26_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid935: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid935_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid935_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_copy936_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_copy936_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid937_In0_c1 <= "" & bh7_w64_23_c1 & bh7_w64_24_c1 & bh7_w64_25_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid937_In1_c1 <= "" & bh7_w65_18_c1 & bh7_w65_19_c1;
   bh7_w64_27_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1(0);
   bh7_w65_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1(1);
   bh7_w66_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid937: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid937_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid937_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_copy938_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_copy938_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid939_In0_c1 <= "" & bh7_w66_22_c1 & bh7_w66_23_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid939_In1_c1 <= "" & bh7_w67_20_c1 & bh7_w67_21_c1;
   bh7_w66_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1(0);
   bh7_w67_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1(1);
   bh7_w68_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid939: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid939_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid939_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_copy940_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_copy940_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid941_In0_c1 <= "" & bh7_w68_22_c1 & bh7_w68_21_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid941_In1_c1 <= "" & bh7_w69_19_c1 & bh7_w69_20_c1;
   bh7_w68_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1(0);
   bh7_w69_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1(1);
   bh7_w70_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid941: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid941_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid941_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_copy942_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_copy942_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid943_In0_c1 <= "" & bh7_w71_19_c1 & bh7_w71_20_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid943_In1_c1 <= "" & bh7_w72_23_c1 & bh7_w72_24_c1;
   bh7_w71_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1(0);
   bh7_w72_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1(1);
   bh7_w73_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid943: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid943_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid943_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_copy944_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_copy944_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid945_In0_c1 <= "" & bh7_w73_18_c1 & bh7_w73_17_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid945_In1_c1 <= "" & bh7_w74_24_c1 & bh7_w74_25_c1;
   bh7_w73_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1(0);
   bh7_w74_26_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1(1);
   bh7_w75_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid945: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid945_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid945_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_copy946_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_copy946_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid947_In0_c1 <= "" & bh7_w75_17_c1 & bh7_w75_16_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid947_In1_c1 <= "" & bh7_w76_22_c1 & bh7_w76_23_c1;
   bh7_w75_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1(0);
   bh7_w76_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1(1);
   bh7_w77_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid947: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid947_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid947_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_copy948_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_copy948_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid949_In0_c1 <= "" & bh7_w78_22_c1 & bh7_w78_23_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid949_In1_c1 <= "" & bh7_w79_17_c1;
   bh7_w78_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1(0);
   bh7_w79_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1(1);
   bh7_w80_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid949: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid949_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid949_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_copy950_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_copy950_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid951_In0_c1 <= "" & bh7_w80_22_c1 & bh7_w80_23_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid951_In1_c1 <= "" & bh7_w81_17_c1;
   bh7_w80_25_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1(0);
   bh7_w81_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1(1);
   bh7_w82_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid951: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid951_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid951_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_copy952_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_copy952_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid953_In0_c1 <= "" & bh7_w82_22_c1 & bh7_w82_23_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid953_In1_c1 <= "" & bh7_w83_15_c1 & bh7_w83_16_c1;
   bh7_w82_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1(0);
   bh7_w83_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1(1);
   bh7_w84_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid953: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid953_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid953_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_copy954_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_copy954_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid955_In0_c1 <= "" & bh7_w86_19_c1 & bh7_w86_20_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid955_In1_c1 <= "" & bh7_w87_18_c1;
   bh7_w86_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1(0);
   bh7_w87_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1(1);
   bh7_w88_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid955: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid955_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid955_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_copy956_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_copy956_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid957_In0_c1 <= "" & bh7_w88_19_c1 & bh7_w88_20_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid957_In1_c1 <= "" & bh7_w89_16_c1;
   bh7_w88_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1(0);
   bh7_w89_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1(1);
   bh7_w90_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid957: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid957_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid957_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_copy958_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_copy958_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid959_In0_c1 <= "" & bh7_w90_19_c1 & bh7_w90_20_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid959_In1_c1 <= "" & bh7_w91_17_c1;
   bh7_w90_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1(0);
   bh7_w91_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1(1);
   bh7_w92_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid959: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid959_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid959_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_copy960_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_copy960_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid961_In0_c1 <= "" & bh7_w92_17_c1 & bh7_w92_18_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid961_In1_c1 <= "" & bh7_w93_19_c1;
   bh7_w92_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1(0);
   bh7_w93_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1(1);
   bh7_w94_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid961: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid961_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid961_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_copy962_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_copy962_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid963_In0_c1 <= "" & bh7_w94_16_c1 & bh7_w94_17_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid963_In1_c1 <= "" & bh7_w95_17_c1;
   bh7_w94_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1(0);
   bh7_w95_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1(1);
   bh7_w96_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid963: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid963_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid963_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_copy964_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_copy964_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid965_In0_c1 <= "" & bh7_w97_16_c1 & bh7_w97_17_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid965_In1_c1 <= "" & bh7_w98_17_c1;
   bh7_w97_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1(0);
   bh7_w98_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1(1);
   bh7_w99_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid965: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid965_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid965_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_copy966_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_copy966_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid967_In0_c1 <= "" & bh7_w100_14_c1 & bh7_w100_15_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid967_In1_c1 <= "" & bh7_w101_12_c1;
   bh7_w100_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1(0);
   bh7_w101_13_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1(1);
   bh7_w102_13_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid967: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid967_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid967_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_copy968_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_copy968_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid969_In0_c1 <= "" & bh7_w102_11_c1 & bh7_w102_12_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid969_In1_c1 <= "" & bh7_w103_10_c1;
   bh7_w102_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1(0);
   bh7_w103_11_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1(1);
   bh7_w104_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid969: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid969_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid969_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_copy970_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_copy970_c1; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh7_22_c1 <= bh7_w22_4_c1 & bh7_w21_6_c1 & bh7_w20_3_c1 & bh7_w19_4_c1 & bh7_w18_2_c1 & bh7_w17_2_c1 & bh7_w16_0_c1 & bh7_w15_0_c1 & bh7_w14_0_c1 & bh7_w13_0_c1 & bh7_w12_0_c1 & bh7_w11_0_c1 & bh7_w10_0_c1 & bh7_w9_0_c1 & bh7_w8_0_c1 & bh7_w7_0_c1 & bh7_w6_0_c1 & bh7_w5_0_c1 & bh7_w4_0_c1 & bh7_w3_0_c1 & bh7_w2_0_c1 & bh7_w1_0_c1 & bh7_w0_0_c1;

   bitheapFinalAdd_bh7_In0_c1 <= "0" & bh7_w105_9_c1 & bh7_w104_7_c1 & bh7_w103_11_c1 & bh7_w102_13_c1 & bh7_w101_13_c1 & bh7_w100_16_c1 & bh7_w99_17_c1 & bh7_w98_18_c1 & bh7_w97_18_c1 & bh7_w96_19_c1 & bh7_w95_18_c1 & bh7_w94_18_c1 & bh7_w93_20_c1 & bh7_w92_19_c1 & bh7_w91_18_c1 & bh7_w90_21_c1 & bh7_w89_17_c1 & bh7_w88_21_c1 & bh7_w87_19_c1 & bh7_w86_21_c1 & bh7_w85_17_c1 & bh7_w84_21_c1 & bh7_w83_17_c1 & bh7_w82_24_c1 & bh7_w81_18_c1 & bh7_w80_24_c1 & bh7_w79_18_c1 & bh7_w78_24_c1 & bh7_w77_17_c1 & bh7_w76_24_c1 & bh7_w75_18_c1 & bh7_w74_26_c1 & bh7_w73_19_c1 & bh7_w72_25_c1 & bh7_w71_21_c1 & bh7_w70_22_c1 & bh7_w69_21_c1 & bh7_w68_23_c1 & bh7_w67_22_c1 & bh7_w66_24_c1 & bh7_w65_20_c1 & bh7_w64_26_c1 & bh7_w63_25_c1 & bh7_w62_22_c1 & bh7_w61_25_c1 & bh7_w60_24_c1 & bh7_w59_23_c1 & bh7_w58_25_c1 & bh7_w57_25_c1 & bh7_w56_21_c1 & bh7_w55_22_c1 & bh7_w54_22_c1 & bh7_w53_19_c1 & bh7_w52_18_c1 & bh7_w51_15_c1 & bh7_w50_13_c1 & bh7_w49_9_c1 & bh7_w48_11_c1 & bh7_w47_7_c1 & bh7_w46_10_c1 & bh7_w45_7_c1 & bh7_w44_10_c1 & bh7_w43_7_c1 & bh7_w42_10_c1 & bh7_w41_7_c1 & bh7_w40_10_c1 & bh7_w39_7_c1 & bh7_w38_9_c1 & bh7_w37_6_c1 & bh7_w36_9_c1 & bh7_w35_9_c1 & bh7_w34_7_c1 & bh7_w33_7_c1 & bh7_w32_6_c1 & bh7_w31_7_c1 & bh7_w30_6_c1 & bh7_w29_7_c1 & bh7_w28_6_c1 & bh7_w27_7_c1 & bh7_w26_6_c1 & bh7_w25_7_c1 & bh7_w24_6_c1 & bh7_w23_7_c1;
   bitheapFinalAdd_bh7_In1_c1 <= "0" & "0" & bh7_w104_8_c1 & "0" & bh7_w102_14_c1 & "0" & "0" & bh7_w99_18_c1 & "0" & "0" & bh7_w96_20_c1 & "0" & bh7_w94_19_c1 & "0" & bh7_w92_20_c1 & "0" & bh7_w90_22_c1 & "0" & bh7_w88_22_c1 & "0" & "0" & "0" & bh7_w84_22_c1 & "0" & bh7_w82_25_c1 & "0" & bh7_w80_25_c1 & "0" & "0" & bh7_w77_18_c1 & "0" & bh7_w75_19_c1 & "0" & bh7_w73_20_c1 & "0" & "0" & bh7_w70_23_c1 & "0" & bh7_w68_24_c1 & "0" & bh7_w66_25_c1 & "0" & bh7_w64_27_c1 & "0" & bh7_w62_23_c1 & "0" & bh7_w60_25_c1 & "0" & bh7_w58_26_c1 & "0" & bh7_w56_22_c1 & "0" & bh7_w54_21_c1 & "0" & bh7_w52_17_c1 & "0" & bh7_w50_12_c1 & "0" & bh7_w48_10_c1 & "0" & bh7_w46_9_c1 & "0" & bh7_w44_9_c1 & "0" & bh7_w42_9_c1 & "0" & bh7_w40_9_c1 & "0" & "0" & bh7_w37_7_c1 & "0" & bh7_w35_8_c1 & "0" & bh7_w33_6_c1 & "0" & bh7_w31_6_c1 & "0" & bh7_w29_6_c1 & "0" & bh7_w27_6_c1 & "0" & bh7_w25_6_c1 & "0" & bh7_w23_6_c1;
   bitheapFinalAdd_bh7_Cin_c0 <= '0';

   bitheapFinalAdd_bh7: IntAdder_84_Freq300_uid972
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 Cin => bitheapFinalAdd_bh7_Cin_c0,
                 X => bitheapFinalAdd_bh7_In0_c1,
                 Y => bitheapFinalAdd_bh7_In1_c1,
                 R => bitheapFinalAdd_bh7_Out_c2);
   bitheapResult_bh7_c2 <= bitheapFinalAdd_bh7_Out_c2(82 downto 0) & tmp_bitheapResult_bh7_22_c2;
   R <= bitheapResult_bh7_c2(105 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_65_Freq300_uid975
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_65_Freq300_uid975 is
    port (clk, ce_1, ce_2, ce_3 : in std_logic;
          X : in  std_logic_vector(64 downto 0);
          Y : in  std_logic_vector(64 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(64 downto 0)   );
end entity;

architecture arch of IntAdder_65_Freq300_uid975 is
signal Cin_1_c2, Cin_1_c3 :  std_logic;
signal X_1_c2, X_1_c3 :  std_logic_vector(65 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3 :  std_logic_vector(65 downto 0);
signal S_1_c3 :  std_logic_vector(65 downto 0);
signal R_1_c3 :  std_logic_vector(64 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_1_c1 <= Y_1_c0;
            end if;
            if ce_2 = '1' then
               Y_1_c2 <= Y_1_c1;
            end if;
            if ce_3 = '1' then
               Cin_1_c3 <= Cin_1_c2;
               X_1_c3 <= X_1_c2;
               Y_1_c3 <= Y_1_c2;
            end if;
         end if;
      end process;
   Cin_1_c2 <= Cin;
   X_1_c2 <= '0' & X(64 downto 0);
   Y_1_c0 <= '0' & Y(64 downto 0);
   S_1_c3 <= X_1_c3 + Y_1_c3 + Cin_1_c3;
   R_1_c3 <= S_1_c3(64 downto 0);
   R <= R_1_c3 ;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointMultiplier
--                      (FPMult_11_52_uid2_Freq300_uid3)
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointMultiplier is
    port (clk, ce_1, ce_2, ce_3 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointMultiplier is
   component IntMultiplier_53x53_106_Freq300_uid5 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             Y : in  std_logic_vector(52 downto 0);
             R : out  std_logic_vector(105 downto 0)   );
   end component;

   component IntAdder_65_Freq300_uid975 is
      port ( clk, ce_1, ce_2, ce_3 : in std_logic;
             X : in  std_logic_vector(64 downto 0);
             Y : in  std_logic_vector(64 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(64 downto 0)   );
   end component;

signal sign_c0, sign_c1, sign_c2, sign_c3 :  std_logic;
signal expX_c0 :  std_logic_vector(10 downto 0);
signal expY_c0 :  std_logic_vector(10 downto 0);
signal expSumPreSub_c0 :  std_logic_vector(12 downto 0);
signal bias_c0 :  std_logic_vector(12 downto 0);
signal expSum_c0, expSum_c1, expSum_c2 :  std_logic_vector(12 downto 0);
signal sigX_c0 :  std_logic_vector(52 downto 0);
signal sigY_c0 :  std_logic_vector(52 downto 0);
signal sigProd_c2 :  std_logic_vector(105 downto 0);
signal excSel_c0 :  std_logic_vector(3 downto 0);
signal exc_c0, exc_c1, exc_c2, exc_c3 :  std_logic_vector(1 downto 0);
signal norm_c2 :  std_logic;
signal expPostNorm_c2 :  std_logic_vector(12 downto 0);
signal sigProdExt_c2 :  std_logic_vector(105 downto 0);
signal expSig_c2 :  std_logic_vector(64 downto 0);
signal sticky_c2 :  std_logic;
signal guard_c2 :  std_logic;
signal round_c2 :  std_logic;
signal expSigPostRound_c3 :  std_logic_vector(64 downto 0);
signal excPostNorm_c3 :  std_logic_vector(1 downto 0);
signal finalExc_c3 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               sign_c1 <= sign_c0;
               expSum_c1 <= expSum_c0;
               exc_c1 <= exc_c0;
            end if;
            if ce_2 = '1' then
               sign_c2 <= sign_c1;
               expSum_c2 <= expSum_c1;
               exc_c2 <= exc_c1;
            end if;
            if ce_3 = '1' then
               sign_c3 <= sign_c2;
               exc_c3 <= exc_c2;
            end if;
         end if;
      end process;
   sign_c0 <= X(63) xor Y(63);
   expX_c0 <= X(62 downto 52);
   expY_c0 <= Y(62 downto 52);
   expSumPreSub_c0 <= ("00" & expX_c0) + ("00" & expY_c0);
   bias_c0 <= CONV_STD_LOGIC_VECTOR(1023,13);
   expSum_c0 <= expSumPreSub_c0 - bias_c0;
   sigX_c0 <= "1" & X(51 downto 0);
   sigY_c0 <= "1" & Y(51 downto 0);
   SignificandMultiplication: IntMultiplier_53x53_106_Freq300_uid5
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => sigX_c0,
                 Y => sigY_c0,
                 R => sigProd_c2);
   excSel_c0 <= X(65 downto 64) & Y(65 downto 64);
   with excSel_c0  select  
   exc_c0 <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm_c2 <= sigProd_c2(105);
   -- exponent update
   expPostNorm_c2 <= expSum_c2 + ("000000000000" & norm_c2);
   -- significand normalization shift
   sigProdExt_c2 <= sigProd_c2(104 downto 0) & "0" when norm_c2='1' else
                         sigProd_c2(103 downto 0) & "00";
   expSig_c2 <= expPostNorm_c2 & sigProdExt_c2(105 downto 54);
   sticky_c2 <= sigProdExt_c2(53);
   guard_c2 <= '0' when sigProdExt_c2(52 downto 0)="00000000000000000000000000000000000000000000000000000" else '1';
   round_c2 <= sticky_c2 and ( (guard_c2 and not(sigProdExt_c2(54))) or (sigProdExt_c2(54) ))  ;
   RoundingAdder: IntAdder_65_Freq300_uid975
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 Cin => round_c2,
                 X => expSig_c2,
                 Y => "00000000000000000000000000000000000000000000000000000000000000000",
                 R => expSigPostRound_c3);
   with expSigPostRound_c3(64 downto 63)  select 
   excPostNorm_c3 <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_c3  select  
   finalExc_c3 <= exc_c3 when  "11"|"10"|"00",
                       excPostNorm_c3 when others; 
   R <= finalExc_c3 & sign_c3 & expSigPostRound_c3(62 downto 0);
end architecture;



