--------------------------------------------------------------------------------
--                  FixRealKCM_Freq300_uid8_T0_Freq300_uid11
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid8_T0_Freq300_uid11 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid8_T0_Freq300_uid11 is
signal Y0 :  std_logic_vector(14 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(14 downto 0);
begin
   with X  select  Y0 <= 
      "000000000001000" when "00000",
      "000001011101011" when "00001",
      "000010111001101" when "00010",
      "000100010110000" when "00011",
      "000101110010011" when "00100",
      "000111001110101" when "00101",
      "001000101011000" when "00110",
      "001010000111011" when "00111",
      "001011100011101" when "01000",
      "001101000000000" when "01001",
      "001110011100011" when "01010",
      "001111111000101" when "01011",
      "010001010101000" when "01100",
      "010010110001011" when "01101",
      "010100001101101" when "01110",
      "010101101010000" when "01111",
      "010111000110011" when "10000",
      "011000100010101" when "10001",
      "011001111111000" when "10010",
      "011011011011011" when "10011",
      "011100110111101" when "10100",
      "011110010100000" when "10101",
      "011111110000011" when "10110",
      "100001001100101" when "10111",
      "100010101001000" when "11000",
      "100100000101010" when "11001",
      "100101100001101" when "11010",
      "100110111110000" when "11011",
      "101000011010010" when "11100",
      "101001110110101" when "11101",
      "101011010011000" when "11110",
      "101100101111010" when "11111",
      "---------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                  FixRealKCM_Freq300_uid8_T1_Freq300_uid14
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid8_T1_Freq300_uid14 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid8_T1_Freq300_uid14 is
signal Y0 :  std_logic_vector(9 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(9 downto 0);
begin
   with X  select  Y0 <= 
      "0000000000" when "00000",
      "0000010111" when "00001",
      "0000101110" when "00010",
      "0001000101" when "00011",
      "0001011100" when "00100",
      "0001110011" when "00101",
      "0010001010" when "00110",
      "0010100010" when "00111",
      "0010111001" when "01000",
      "0011010000" when "01001",
      "0011100111" when "01010",
      "0011111110" when "01011",
      "0100010101" when "01100",
      "0100101100" when "01101",
      "0101000011" when "01110",
      "0101011010" when "01111",
      "0101110001" when "10000",
      "0110001000" when "10001",
      "0110011111" when "10010",
      "0110110111" when "10011",
      "0111001110" when "10100",
      "0111100101" when "10101",
      "0111111100" when "10110",
      "1000010011" when "10111",
      "1000101010" when "11000",
      "1001000001" when "11001",
      "1001011000" when "11010",
      "1001101111" when "11011",
      "1010000110" when "11100",
      "1010011101" when "11101",
      "1010110100" when "11110",
      "1011001100" when "11111",
      "----------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                  FixRealKCM_Freq300_uid8_T2_Freq300_uid17
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid8_T2_Freq300_uid17 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid8_T2_Freq300_uid17 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "000",
      "00011" when "001",
      "00110" when "010",
      "01001" when "011",
      "01100" when "100",
      "01110" when "101",
      "10001" when "110",
      "10100" when "111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq300_uid21
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid21 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid21 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq300_uid35_T0_Freq300_uid38
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid35_T0_Freq300_uid38 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(66 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid35_T0_Freq300_uid38 is
signal Y0 :  std_logic_vector(66 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(66 downto 0);
begin
   with X  select  Y0 <= 
      "0000000000000000000000000000000000000000000000000000000000000000000" when "00000",
      "0000010110001011100100001011111110111110100011100111101111001101011" when "00001",
      "0000101100010111001000010111111101111101000111001111011110011010110" when "00010",
      "0001000010100010101100100011111100111011101010110111001101101000001" when "00011",
      "0001011000101110010000101111111011111010001110011110111100110101100" when "00100",
      "0001101110111001110100111011111010111000110010000110101100000010111" when "00101",
      "0010000101000101011001000111111001110111010101101110011011010000010" when "00110",
      "0010011011010000111101010011111000110101111001010110001010011101101" when "00111",
      "0010110001011100100001011111110111110100011100111101111001101011000" when "01000",
      "0011000111101000000101101011110110110011000000100101101000111000011" when "01001",
      "0011011101110011101001110111110101110001100100001101011000000101101" when "01010",
      "0011110011111111001110000011110100110000000111110101000111010011000" when "01011",
      "0100001010001010110010001111110011101110101011011100110110100000011" when "01100",
      "0100100000010110010110011011110010101101001111000100100101101101110" when "01101",
      "0100110110100001111010100111110001101011110010101100010100111011001" when "01110",
      "0101001100101101011110110011110000101010010110010100000100001000100" when "01111",
      "0101100010111001000010111111101111101000111001111011110011010101111" when "10000",
      "0101111001000100100111001011101110100111011101100011100010100011010" when "10001",
      "0110001111010000001011010111101101100110000001001011010001110000101" when "10010",
      "0110100101011011101111100011101100100100100100110011000000111110000" when "10011",
      "0110111011100111010011101111101011100011001000011010110000001011011" when "10100",
      "0111010001110010110111111011101010100001101100000010011111011000110" when "10101",
      "0111100111111110011100000111101001100000001111101010001110100110001" when "10110",
      "0111111110001010000000010011101000011110110011010001111101110011100" when "10111",
      "1000010100010101100100011111100111011101010110111001101101000000111" when "11000",
      "1000101010100001001000101011100110011011111010100001011100001110010" when "11001",
      "1001000000101100101100110111100101011010011110001001001011011011101" when "11010",
      "1001010110111000010001000011100100011001000001110000111010101001000" when "11011",
      "1001101101000011110101001111100011010111100101011000101001110110011" when "11100",
      "1010000011001111011001011011100010010110001001000000011001000011101" when "11101",
      "1010011001011010111101100111100001010100101100101000001000010001000" when "11110",
      "1010101111100110100001110011100000010011010000001111110111011110011" when "11111",
      "-------------------------------------------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq300_uid35_T1_Freq300_uid41
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid35_T1_Freq300_uid41 is
    port (X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(61 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid35_T1_Freq300_uid41 is
signal Y0 :  std_logic_vector(61 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(61 downto 0);
begin
   with X  select  Y0 <= 
      "00000000000000000000000000000000000000000000000000000000000000" when "000000",
      "00000010110001011100100001011111110111110100011100111101111010" when "000001",
      "00000101100010111001000010111111101111101000111001111011110011" when "000010",
      "00001000010100010101100100011111100111011101010110111001101101" when "000011",
      "00001011000101110010000101111111011111010001110011110111100111" when "000100",
      "00001101110111001110100111011111010111000110010000110101100000" when "000101",
      "00010000101000101011001000111111001110111010101101110011011010" when "000110",
      "00010011011010000111101010011111000110101111001010110001010100" when "000111",
      "00010110001011100100001011111110111110100011100111101111001101" when "001000",
      "00011000111101000000101101011110110110011000000100101101000111" when "001001",
      "00011011101110011101001110111110101110001100100001101011000001" when "001010",
      "00011110011111111001110000011110100110000000111110101000111010" when "001011",
      "00100001010001010110010001111110011101110101011011100110110100" when "001100",
      "00100100000010110010110011011110010101101001111000100100101110" when "001101",
      "00100110110100001111010100111110001101011110010101100010100111" when "001110",
      "00101001100101101011110110011110000101010010110010100000100001" when "001111",
      "00101100010111001000010111111101111101000111001111011110011011" when "010000",
      "00101111001000100100111001011101110100111011101100011100010100" when "010001",
      "00110001111010000001011010111101101100110000001001011010001110" when "010010",
      "00110100101011011101111100011101100100100100100110011000001000" when "010011",
      "00110111011100111010011101111101011100011001000011010110000001" when "010100",
      "00111010001110010110111111011101010100001101100000010011111011" when "010101",
      "00111100111111110011100000111101001100000001111101010001110101" when "010110",
      "00111111110001010000000010011101000011110110011010001111101110" when "010111",
      "01000010100010101100100011111100111011101010110111001101101000" when "011000",
      "01000101010100001001000101011100110011011111010100001011100010" when "011001",
      "01001000000101100101100110111100101011010011110001001001011011" when "011010",
      "01001010110111000010001000011100100011001000001110000111010101" when "011011",
      "01001101101000011110101001111100011010111100101011000101001111" when "011100",
      "01010000011001111011001011011100010010110001001000000011001000" when "011101",
      "01010011001011010111101100111100001010100101100101000001000010" when "011110",
      "01010101111100110100001110011100000010011010000001111110111100" when "011111",
      "01011000101110010000101111111011111010001110011110111100110101" when "100000",
      "01011011011111101101010001011011110010000010111011111010101111" when "100001",
      "01011110010001001001110010111011101001110111011000111000101001" when "100010",
      "01100001000010100110010100011011100001101011110101110110100010" when "100011",
      "01100011110100000010110101111011011001100000010010110100011100" when "100100",
      "01100110100101011111010111011011010001010100101111110010010110" when "100101",
      "01101001010110111011111000111011001001001001001100110000001111" when "100110",
      "01101100001000011000011010011011000000111101101001101110001001" when "100111",
      "01101110111001110100111011111010111000110010000110101100000011" when "101000",
      "01110001101011010001011101011010110000100110100011101001111101" when "101001",
      "01110100011100101101111110111010101000011011000000100111110110" when "101010",
      "01110111001110001010100000011010100000001111011101100101110000" when "101011",
      "01111001111111100111000001111010011000000011111010100011101010" when "101100",
      "01111100110001000011100011011010001111111000010111100001100011" when "101101",
      "01111111100010100000000100111010000111101100110100011111011101" when "101110",
      "10000010010011111100100110011001111111100001010001011101010111" when "101111",
      "10000101000101011001000111111001110111010101101110011011010000" when "110000",
      "10000111110110110101101001011001101111001010001011011001001010" when "110001",
      "10001010101000010010001010111001100110111110101000010111000100" when "110010",
      "10001101011001101110101100011001011110110011000101010100111101" when "110011",
      "10010000001011001011001101111001010110100111100010010010110111" when "110100",
      "10010010111100100111101111011001001110011011111111010000110001" when "110101",
      "10010101101110000100010000111001000110010000011100001110101010" when "110110",
      "10011000011111100000110010011000111110000100111001001100100100" when "110111",
      "10011011010000111101010011111000110101111001010110001010011110" when "111000",
      "10011110000010011001110101011000101101101101110011001000010111" when "111001",
      "10100000110011110110010110111000100101100010010000000110010001" when "111010",
      "10100011100101010010111000011000011101010110101101000100001011" when "111011",
      "10100110010110101111011001111000010101001011001010000010000100" when "111100",
      "10101001001000001011111011011000001100111111100110111111111110" when "111101",
      "10101011111001101000011100111000000100110100000011111101111000" when "111110",
      "10101110101011000100111110010111111100101000100000111011110001" when "111111",
      "--------------------------------------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--          compressedTable_Freq300_uid52_subsampling_Freq300_uid54
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity compressedTable_Freq300_uid52_subsampling_Freq300_uid54 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of compressedTable_Freq300_uid52_subsampling_Freq300_uid54 is
signal Y0 :  std_logic_vector(8 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(8 downto 0);
begin
   with X  select  Y0 <= 
      "100000000" when "0000000",
      "100000010" when "0000001",
      "100000100" when "0000010",
      "100000110" when "0000011",
      "100001000" when "0000100",
      "100001010" when "0000101",
      "100001100" when "0000110",
      "100001110" when "0000111",
      "100010000" when "0001000",
      "100010010" when "0001001",
      "100010100" when "0001010",
      "100010110" when "0001011",
      "100011001" when "0001100",
      "100011011" when "0001101",
      "100011101" when "0001110",
      "100011111" when "0001111",
      "100100010" when "0010000",
      "100100100" when "0010001",
      "100100110" when "0010010",
      "100101000" when "0010011",
      "100101011" when "0010100",
      "100101101" when "0010101",
      "100110000" when "0010110",
      "100110010" when "0010111",
      "100110100" when "0011000",
      "100110111" when "0011001",
      "100111001" when "0011010",
      "100111100" when "0011011",
      "100111110" when "0011100",
      "101000001" when "0011101",
      "101000011" when "0011110",
      "101000110" when "0011111",
      "101001000" when "0100000",
      "101001011" when "0100001",
      "101001101" when "0100010",
      "101010000" when "0100011",
      "101010011" when "0100100",
      "101010101" when "0100101",
      "101011000" when "0100110",
      "101011011" when "0100111",
      "101011101" when "0101000",
      "101100000" when "0101001",
      "101100011" when "0101010",
      "101100110" when "0101011",
      "101101001" when "0101100",
      "101101011" when "0101101",
      "101101110" when "0101110",
      "101110001" when "0101111",
      "101110100" when "0110000",
      "101110111" when "0110001",
      "101111010" when "0110010",
      "101111101" when "0110011",
      "110000000" when "0110100",
      "110000011" when "0110101",
      "110000110" when "0110110",
      "110001001" when "0110111",
      "110001100" when "0111000",
      "110001111" when "0111001",
      "110010010" when "0111010",
      "110010101" when "0111011",
      "110011001" when "0111100",
      "110011100" when "0111101",
      "110011111" when "0111110",
      "110100010" when "0111111",
      "010011011" when "1000000",
      "010011100" when "1000001",
      "010011101" when "1000010",
      "010011110" when "1000011",
      "010100000" when "1000100",
      "010100001" when "1000101",
      "010100010" when "1000110",
      "010100011" when "1000111",
      "010100101" when "1001000",
      "010100110" when "1001001",
      "010100111" when "1001010",
      "010101001" when "1001011",
      "010101010" when "1001100",
      "010101011" when "1001101",
      "010101101" when "1001110",
      "010101110" when "1001111",
      "010101111" when "1010000",
      "010110001" when "1010001",
      "010110010" when "1010010",
      "010110100" when "1010011",
      "010110101" when "1010100",
      "010110110" when "1010101",
      "010111000" when "1010110",
      "010111001" when "1010111",
      "010111011" when "1011000",
      "010111100" when "1011001",
      "010111110" when "1011010",
      "010111111" when "1011011",
      "011000001" when "1011100",
      "011000010" when "1011101",
      "011000100" when "1011110",
      "011000101" when "1011111",
      "011000111" when "1100000",
      "011001000" when "1100001",
      "011001010" when "1100010",
      "011001100" when "1100011",
      "011001101" when "1100100",
      "011001111" when "1100101",
      "011010000" when "1100110",
      "011010010" when "1100111",
      "011010100" when "1101000",
      "011010101" when "1101001",
      "011010111" when "1101010",
      "011011001" when "1101011",
      "011011010" when "1101100",
      "011011100" when "1101101",
      "011011110" when "1101110",
      "011100000" when "1101111",
      "011100001" when "1110000",
      "011100011" when "1110001",
      "011100101" when "1110010",
      "011100111" when "1110011",
      "011101001" when "1110100",
      "011101010" when "1110101",
      "011101100" when "1110110",
      "011101110" when "1110111",
      "011110000" when "1111000",
      "011110010" when "1111001",
      "011110100" when "1111010",
      "011110110" when "1111011",
      "011111000" when "1111100",
      "011111010" when "1111101",
      "011111100" when "1111110",
      "011111110" when "1111111",
      "---------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          coeffTable_Freq300_uid61
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity coeffTable_Freq300_uid61 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(94 downto 0)   );
end entity;

architecture arch of coeffTable_Freq300_uid61 is
signal Y0 :  std_logic_vector(94 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(94 downto 0);
begin
   with X  select  Y0 <= 
      "00000000000000010000000000000000001001100000001000000000000000000101000100000000000000000100000" when "0000000",
      "00000000000010010000000000000010010100000000011000000000000000100101000100000000000000001100000" when "0000001",
      "00000000000110010000000000001010011110100000101000000000000001100101000100000000000000010100000" when "0000010",
      "00000000001100010000000000011100101001100000111000000000000011000101000100000000000000011100000" when "0000011",
      "00000000010100010000000000111100110100000001001000000000000101000101000100000000000000100100000" when "0000100",
      "00000000011110010000000001101110111110100001011000000000000111100101000100000000000000101100001" when "0000101",
      "00000000101010010000000010110111001001100001101000000000001010100101000100000000000000110100000" when "0000110",
      "00000000111000010000000100011001010100100001111000000000001110000101000100000000000000111011111" when "0000111",
      "00000001001000010000000110011001011111000010001000000000010010000101000100000000000001000100000" when "0001000",
      "00000001011010010000001000111011101010000010011000000000010110100101000100000000000001001100000" when "0001001",
      "00000001101110010000001100000011110101000010101000000000011011100101000100000000000001010100000" when "0001010",
      "00000010000100010000001111110110000000000010111000000000100001000101000100000000000001011100000" when "0001011",
      "00000010011100010000010100010110001011100011001000000000100111000101001100000000000001100100000" when "0001100",
      "00000010110110010000011001101000010110100011011000000000101101100101001100000000000001101100001" when "0001101",
      "00000011010010010000011111110000100010100011101000000000110100100101001100000000000001110011111" when "0001110",
      "00000011110000010000100110110010101110000011111000000000111100000101001100000000000001111100000" when "0001111",
      "00000100010000010000101110110010111010000100001000000001000100000101001100000000000010000100000" when "0010000",
      "00000100110010010000110111110101000110100100011000000001001100100101010100000000000010001100000" when "0010001",
      "00000101010110010001000001111101010011000100101000000001010101100101010100000000000010010100000" when "0010010",
      "00000101111100010001001101001111100000000100111000000001011111000101010100000000000010011011111" when "0010011",
      "00000110100100010001011001101111101101000101001000000001101001000101011100000000000010100100000" when "0010100",
      "00000111001110010001100111100001111010100101011000000001110011100101011100000000000010101100001" when "0010101",
      "00000111111010010001110110101010001001000101101000000001111110100101100100000000000010110100000" when "0010110",
      "00001000101000010010000111001100010111100101111000000010001010000101100100000000000010111100000" when "0010111",
      "00001001011000010010011001001100100110100110001000000010010110000101101100000000000011000100001" when "0011000",
      "00001010001010010010101100101110110110100110011000000010100010100101101100000000000011001100000" when "0011001",
      "00001010111110010011000001110111000111000110101000000010101111100101110100000000000011010100000" when "0011010",
      "00001011110100010011011000101001011000000110111000000010111101000101111100000000000011011100000" when "0011011",
      "00001100101100010011110001001001101001100111001000000011001011000110000100000000000011100100001" when "0011100",
      "00001101100110010100001011011011111100100111011000000011011001100110000100000000000011101100000" when "0011101",
      "00001110100010010100100111100100010000000111101000000011101000100110001100000000000011110100000" when "0011110",
      "00001111100000010101000101100110100100000111111000000011111000000110010100000000000011111100001" when "0011111",
      "00010000100000010101100101100110111001101000001000000100001000000110011100000000000100000100000" when "0100000",
      "00010001100010010110000111101001010000001000011000000100011000100110100100000000000100001100000" when "0100001",
      "00010010100110010110101011110001100111101000101000000100101001100110101100000000000100010100000" when "0100010",
      "00010011101100010111010010000100000000001000111000000100111011000110111100000000000100011100000" when "0100011",
      "00010100110100010111111010100100011010001001001000000101001101000111000100000000000100100100000" when "0100100",
      "00010101111110011000100101010110110101001001011000000101011111100111001100000000000100101100000" when "0100101",
      "00010111001010011001010010011111010001101001101000000101110010100111011100000000000100110100000" when "0100110",
      "00011000011000011010000010000001101111101001111000000110000110000111100100000000000100111100000" when "0100111",
      "00011001101000011010110100000010001111001010001000000110011010000111110100000000000101000100000" when "0101000",
      "00011010111010011011101000100100110000001010011000000110101110100111111100000000000101001100001" when "0101001",
      "00011100001110011100011111101101010011001010101000000111000011101000001100000000000101010100000" when "0101010",
      "00011101100100011101011001011111110111101010111000000111011001001000011100000000000101011100000" when "0101011",
      "00011110111100011110010110000000011110001011001000000111101111001000101100000000000101100100000" when "0101100",
      "00100000010110011111010101010011000110001011011000001000000101101000111100000000000101101100001" when "0101101",
      "00100001110010100000010111011011110000101011101000001000011100101001001100000000000101110100001" when "0101110",
      "00100011010000100001011100011110011101001011111000001000110100001001011100000000000101111100000" when "0101111",
      "00100100110000100010100100011111001011101100001000001001001100001001101100000000000110000100001" when "0110000",
      "00100110010010100011101111100001111100101100011000001001100100101001111100000000000110001100001" when "0110001",
      "00100111110110100100111101101010110000001100101000001001111101101010010100000000000110010100001" when "0110010",
      "00101001011100100110001110111101100110001100111000001010010111001010100100000000000110011100000" when "0110011",
      "00101011000100100111100011011110011110101101001000001010110001001010111100000000000110100100000" when "0110100",
      "00101100101110101000111011010001011001101101011000001011001011101011010100000000000110101100001" when "0110101",
      "00101110011010101010010110011010010111101101101000001011100110101011101100000000000110110100000" when "0110110",
      "00110000001000101011110100111101011000001101111000001100000010001100000100000000000110111100001" when "0110111",
      "00110001111000101101010110111110011100001110001000001100011110001100011100000000000111000100001" when "0111000",
      "00110011101010101110111100100001100011001110011000001100111010101100110100000000000111001100001" when "0111001",
      "00110101011110110000100101101010101101001110101000001101010111101101001100000000000111010100001" when "0111010",
      "00110111010100110010010010011101111010101110111000001101110101001101101100000000000111011100001" when "0111011",
      "00111001001100110100000010111111001011101111001000001110010011001110000100000000000111100100001" when "0111100",
      "00111011000110110101110111010010100000101111011000001110110001101110100100000000000111101100000" when "0111101",
      "00111101000010110111101111011011111000101111101000001111010000101110111100000000000111110100001" when "0111110",
      "00111111000000111001101011011111010100101111111000001111110000001111011100000000000111111100001" when "0111111",
      "01000001000000111011101011100000110100110000001000010000010000001111111100000000001000000100001" when "1000000",
      "01000011000010111101101111100100011000110000011000010000110000110000011100000000001000001100010" when "1000001",
      "01000101000110111111110111101110000001010000101000010001010001110001000100000000001000010100001" when "1000010",
      "01000111001101000010000100000001101101110000111000010001110011010001100100000000001000011100001" when "1000011",
      "01001001010101000100010100100011011110110001001000010010010101010010001100000000001000100100001" when "1000100",
      "01001011011111000110101001010111010100010001011000010010110111110010101100000000001000101100010" when "1000101",
      "01001101101011001001000010100001001110110001101000010011011010110011010100000000001000110100001" when "1000110",
      "01001111111001001011100000000101001110010001111000010011111110010011111100000000001000111100001" when "1000111",
      "01010010001001001110000010000111010010010010001000010100100010010100100100000000001001000100001" when "1001000",
      "01010100011011010000101000101011011011110010011000010101000110110101001100000000001001001100001" when "1001001",
      "01010110101111010011010011110101101010010010101000010101101011110101111100000000001001010100001" when "1001010",
      "01011001000101010110000011101001111110010010111000010110010001010110100100000000001001011100001" when "1001011",
      "01011011011101011000111000001100010111110011001000010110110111010111010100000000001001100100001" when "1001100",
      "01011101110111011011110001100000110111010011011000010111011101111000000100000000001001101100001" when "1001101",
      "01100000010011011110101111101011011100010011101000011000000100111000101100000000001001110100001" when "1001110",
      "01100010110001100001110010110000000111010011111000011000101100011001100100000000001001111100010" when "1001111",
      "01100101010001100100111010110010111000110100001000011001010100011010010100000000001010000100010" when "1010000",
      "01100111110011101000000111110111110000010100011000011001111100111011000100000000001010001100010" when "1010001",
      "01101010010111101011011010000010101110110100101000011010100101111011111100000000001010010100001" when "1010010",
      "01101100111101101110110001010111110011010100111000011011001111011100110100000000001010011100010" when "1010011",
      "01101111100101110010001101111010111111010101001000011011111001011101100100000000001010100100001" when "1010100",
      "01110010001111110101101111110000010001110101011000011100100011111110011100000000001010101100010" when "1010101",
      "01110100111011111001010110111011101011110101101000011101001110111111011100000000001010110100001" when "1010110",
      "01110111101001111101000011100001001100110101111000011101111010100000010100000000001010111100001" when "1010111",
      "01111010011010000000110101100100110101010110001000011110100110100001010100000000001011000100010" when "1011000",
      "01111101001100000100101101001010100101010110011000011111010011000010001100000000001011001100010" when "1011001",
      "10000000000000001000101010010110011101010110101000100000000000000011001100000000001011010100010" when "1011010",
      "10000010110110001100101101001100011101010110111000100000101101100100001100000000001011011100010" when "1011011",
      "10000101101110010000110101110000100101110111001000100001011011100101010100000000001011100100010" when "1011100",
      "10001000101000010101000100000110110110010111011000100010001010000110010100000000001011101100010" when "1011101",
      "10001011100100011001011000010011001111010111101000100010111001000111011100000000001011110100010" when "1011110",
      "10001110100010011101110010011001110001010111111000100011101000101000100100000000001011111100010" when "1011111",
      "10010001100010100010010010011110011011111000001000100100011000101001101100000000001100000100010" when "1100000",
      "10010100100100100110111000100101001111111000011000100101001001001010110100000000001100001100010" when "1100001",
      "10010111101000101011100100110010001100111000101000100101111010001011111100000000001100010100010" when "1100010",
      "10011010101110110000010111001001010011011000111000100110101011101101001100000000001100011100010" when "1100011",
      "10011101110110110101001111101110100011111001001000100111011101101110010100000000001100100100010" when "1100100",
      "10100001000000111010001110100101111101111001011000101000010000001111100100000000001100101100010" when "1100101",
      "10100100001100111111010011110011100001111001101000101001000011010000111100000000001100110100011" when "1100110",
      "10100111011011000100011111011011010000011001111000101001110110110010001100000000001100111100011" when "1100111",
      "10101010101011001001110001100001001001011010001000101010101010110011100100000000001101000100011" when "1101000",
      "10101101111101001111001010001001001100111010011000101011011111010100110100000000001101001100011" when "1101001",
      "10110001010001010100101001010111011011011010101000101100010100010110001100000000001101010100011" when "1101010",
      "10110100100111011010001111001111110100111010111000101101001001110111100100000000001101011100011" when "1101011",
      "10110111111111011111111011110110011001111011001000101101111111111001000100000000001101100100010" when "1101100",
      "10111011011001100101101111001111001001111011011000101110110110011010011100000000001101101100011" when "1101101",
      "10111110110101101011101001011110000101111011101000101111101101011011111100000000001101110100100" when "1101110",
      "11000010010011110001101010100111001101111011111000110000100100111101011100000000001101111100011" when "1101111",
      "11000101110011110111110010101110100010011100001000110001011100111111000100000000001110000100010" when "1110000",
      "11001001010101111110000001111000000010011100011000110010010101100000100100000000001110001100100" when "1110001",
      "11001100111010000100011000000111101111111100101000110011001110100010001100000000001110010100011" when "1110010",
      "11010000100000001010110101100001101001011100111000110100001000000011110100000000001110011100100" when "1110011",
      "11010100001000010001011010001001110000011101001000110101000010000101011100000000001110100100011" when "1110100",
      "11010111110010011000000110000100000100011101011000110101111100100111000100000000001110101100100" when "1110101",
      "11011011011110011110111001010100100110011101101000110110110111101000110100000000001110110100011" when "1110110",
      "11011111001100100101110011111111010101011101111000110111110011001010100100000000001110111100100" when "1110111",
      "11100010111100101100110110001000010010111110001000111000101111001100010100000000001111000100100" when "1111000",
      "11100110101110110011111111110011011110011110011000111001101011101110000100000000001111001100100" when "1111001",
      "11101010100010111011010001000100111000011110101000111010101000101111111100000000001111010100011" when "1111010",
      "11101110011001000010101010000000100000111110111000111011100110010001101100000000001111011100100" when "1111011",
      "11110010010001001010001010101010011000011111001000111100100100010011100100000000001111100100100" when "1111100",
      "11110110001011010001110011000110011110111111011000111101100010110101100100000000001111101100100" when "1111101",
      "11111010000111011001100011011000110100111111101000111110100001110111011100000000001111110100100" when "1111110",
      "11111110000101100001011011100101011010011111111000111111100001011001011100000000001111111100100" when "1111111",
      "-----------------------------------------------------------------------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid73
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid73 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid73 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid78
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid78 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid78 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid83
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid83 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid83 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid88
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid88 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid88 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid93
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid93 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid93 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid98
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid98 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid98 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid103
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid103 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid103 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid108
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid108 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid108 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid113
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid113 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid113 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid118
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid118 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid118 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid123
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid128
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid128 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid128 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid133
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid133 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid133 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid138
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid138 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid138 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid143
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid143 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid143 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid148
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid148 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid148 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid153
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid153 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid153 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid158
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid158 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid158 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid163
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid163 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid163 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid168
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid168 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid168 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid173
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid173 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid173 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid178
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid178 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid178 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid183
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid183 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid183 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid188
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid188 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid188 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid193
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid193 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid193 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid198
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid198 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid198 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid203
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid203 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid203 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid208
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid208 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid208 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid213
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid213 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid213 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid218
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid218 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid218 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid223
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid223 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid223 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid228
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid228 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid228 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid233
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid233 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid233 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid238
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid238 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid238 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "1110" when "0110",
      "1111" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "1100" when "1010",
      "1110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "1010" when "1110",
      "1101" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid243
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid243 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid243 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid248
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid248 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid248 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid255
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid255 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid255 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid260
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid260 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid260 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid265
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid265 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid265 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid270
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid270 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid270 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid275
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid275 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid275 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "01000" when "11000",
      "00111" when "11001",
      "00110" when "11010",
      "00101" when "11011",
      "00100" when "11100",
      "00011" when "11101",
      "00010" when "11110",
      "00001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid280
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid280 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid280 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq300_uid284
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid284 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid284 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid288
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid288 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid288 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq300_uid292
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid292 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid292 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid300
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid300 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid300 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq300_uid334
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq300_uid334 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq300_uid334 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid547
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid547 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid547 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid552
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid552 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid552 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid557
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid557 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid557 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid562
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid562 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid562 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid567
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid567 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid567 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid572
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid572 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid572 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid577
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid577 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid577 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid582
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid582 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid582 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid587
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid587 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid587 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid592
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid592 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid592 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid597
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid597 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid597 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid602
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid602 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid602 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid607
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid607 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid607 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid612
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid612 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid612 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid617
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid617 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid617 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid622
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid622 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid622 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid627
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid627 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid627 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid632
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid632 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid632 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid637
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid637 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid637 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid642
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid642 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid642 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid647
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid647 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid647 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid652
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid652 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid652 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid657
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid657 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid657 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid662
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid662 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid662 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid667
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid667 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid667 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid672
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid672 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid672 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid677
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid677 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid677 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid682
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid682 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid682 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid687
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid687 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid687 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "01000" when "11000",
      "00111" when "11001",
      "00110" when "11010",
      "00101" when "11011",
      "00100" when "11100",
      "00011" when "11101",
      "00010" when "11110",
      "00001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid692
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid692 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid692 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid697
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid697 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid697 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00000" when "01001",
      "00000" when "01010",
      "00000" when "01011",
      "00000" when "01100",
      "00000" when "01101",
      "00000" when "01110",
      "00000" when "01111",
      "00000" when "10000",
      "11111" when "10001",
      "11110" when "10010",
      "11101" when "10011",
      "11100" when "10100",
      "11011" when "10101",
      "11010" when "10110",
      "11001" when "10111",
      "11000" when "11000",
      "10111" when "11001",
      "10110" when "11010",
      "10101" when "11011",
      "10100" when "11100",
      "10011" when "11101",
      "10010" when "11110",
      "10001" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid702
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid702 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid702 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "11100" when "01100",
      "11101" when "01101",
      "11110" when "01110",
      "11111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "11000" when "10100",
      "11010" when "10101",
      "11100" when "10110",
      "11110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "10100" when "11100",
      "10111" when "11101",
      "11010" when "11110",
      "11101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid707
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid707 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid707 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid712
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid712 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid712 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid717
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid717 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid717 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid722
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid722 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid722 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "11100" when "01100",
      "11101" when "01101",
      "11110" when "01110",
      "11111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "11000" when "10100",
      "11010" when "10101",
      "11100" when "10110",
      "11110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "10100" when "11100",
      "10111" when "11101",
      "11010" when "11110",
      "11101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid727
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid727 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid727 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid732
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid732 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid732 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid737
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid737 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid737 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid742
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid742 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid742 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "11100" when "01100",
      "11101" when "01101",
      "11110" when "01110",
      "11111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "11000" when "10100",
      "11010" when "10101",
      "11100" when "10110",
      "11110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "10100" when "11100",
      "10111" when "11101",
      "11010" when "11110",
      "11101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid747
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid747 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid747 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid752
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid752 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid752 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid757
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid757 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid757 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid762
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid762 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid762 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "11100" when "01100",
      "11101" when "01101",
      "11110" when "01110",
      "11111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "11000" when "10100",
      "11010" when "10101",
      "11100" when "10110",
      "11110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "10100" when "11100",
      "10111" when "11101",
      "11010" when "11110",
      "11101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid767
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid767 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid767 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid772
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid772 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid772 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid777
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid777 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid777 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq300_uid781
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid781 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid781 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid789
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid789 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid789 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid797
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid797 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid797 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq300_uid813
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid813 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid813 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq300_uid839
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq300_uid839 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq300_uid839 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1122
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1122 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1122 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1131
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1131 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1131 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1138
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1138 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1138 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1143
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1143 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1143 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1150
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1150 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1150 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1155
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1155 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1155 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1160
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1160 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1160 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1169
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1169 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1169 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1174
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1174 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1174 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1179
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1179 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1179 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1186
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1186 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1186 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1191
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1191 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1191 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1196
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1196 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1196 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1201
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1201 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1201 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1214
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1214 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1214 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1223
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1223 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1223 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1230
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1230 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1230 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1235
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1235 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1235 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1242
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1242 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1242 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1247
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1247 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1247 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1252
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1252 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1252 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1261
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1261 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1261 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1266
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1266 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1266 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1271
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1271 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1271 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1276
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1276 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1276 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1281
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1281 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1281 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1286
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1286 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1286 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1291
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1291 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1291 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1296
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1296 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1296 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1301
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1301 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1301 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1306
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1306 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1306 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1311
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1311 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1311 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1316
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1316 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1316 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1321
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1321 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1321 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1326
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1326 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1326 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1331
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1331 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1331 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1336
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1336 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1336 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1341
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1341 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1341 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1346
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1346 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1346 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         MultTable_Freq300_uid1351
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid1351 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid1351 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                      Compressor_23_3_Freq300_uid1355
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid1355 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid1355 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid1359
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid1359 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid1359 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid1363
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid1363 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid1363 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                      Compressor_14_3_Freq300_uid1373
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid1373 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid1373 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq300_uid1557
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq300_uid1557 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq300_uid1557 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                    LeftShifter53_by_max_65_Freq300_uid4
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X S
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter53_by_max_65_Freq300_uid4 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          S : in  std_logic_vector(6 downto 0);
          R : out  std_logic_vector(117 downto 0)   );
end entity;

architecture arch of LeftShifter53_by_max_65_Freq300_uid4 is
signal ps_c0, ps_c1, ps_c2 :  std_logic_vector(6 downto 0);
signal level0_c0 :  std_logic_vector(52 downto 0);
signal level1_c0 :  std_logic_vector(53 downto 0);
signal level2_c0 :  std_logic_vector(55 downto 0);
signal level3_c0, level3_c1 :  std_logic_vector(59 downto 0);
signal level4_c1 :  std_logic_vector(67 downto 0);
signal level5_c1, level5_c2 :  std_logic_vector(83 downto 0);
signal level6_c2 :  std_logic_vector(115 downto 0);
signal level7_c2 :  std_logic_vector(179 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               ps_c1 <= ps_c0;
               level3_c1 <= level3_c0;
            end if;
            if ce_2 = '1' then
               ps_c2 <= ps_c1;
               level5_c2 <= level5_c1;
            end if;
         end if;
      end process;
   ps_c0<= S;
   level0_c0<= X;
   level1_c0<= level0_c0 & (0 downto 0 => '0') when ps_c0(0)= '1' else     (0 downto 0 => '0') & level0_c0;
   level2_c0<= level1_c0 & (1 downto 0 => '0') when ps_c0(1)= '1' else     (1 downto 0 => '0') & level1_c0;
   level3_c0<= level2_c0 & (3 downto 0 => '0') when ps_c0(2)= '1' else     (3 downto 0 => '0') & level2_c0;
   level4_c1<= level3_c1 & (7 downto 0 => '0') when ps_c1(3)= '1' else     (7 downto 0 => '0') & level3_c1;
   level5_c1<= level4_c1 & (15 downto 0 => '0') when ps_c1(4)= '1' else     (15 downto 0 => '0') & level4_c1;
   level6_c2<= level5_c2 & (31 downto 0 => '0') when ps_c2(5)= '1' else     (31 downto 0 => '0') & level5_c2;
   level7_c2<= level6_c2 & (63 downto 0 => '0') when ps_c2(6)= '1' else     (63 downto 0 => '0') & level6_c2;
   R <= level7_c2(117 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_15_Freq300_uid33
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_15_Freq300_uid33 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(14 downto 0);
          Y : in  std_logic_vector(14 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of IntAdder_15_Freq300_uid33 is
signal Rtmp_c2 :  std_logic_vector(14 downto 0);
signal Cin_c1, Cin_c2 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
         end if;
      end process;
   Rtmp_c2 <= X + Y + Cin_c2;
   R <= Rtmp_c2;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq300_uid8
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid8 is
    port (clk : in std_logic;
          X : in  std_logic_vector(12 downto 0);
          R : out  std_logic_vector(10 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid8 is
   component FixRealKCM_Freq300_uid8_T0_Freq300_uid11 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(14 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid8_T1_Freq300_uid14 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(9 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid8_T2_Freq300_uid17 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid21 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_15_Freq300_uid33 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(14 downto 0);
             Y : in  std_logic_vector(14 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(14 downto 0)   );
   end component;

signal FixRealKCM_Freq300_uid8_A0_c2 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq300_uid8_T0_c2 :  std_logic_vector(14 downto 0);
signal FixRealKCM_Freq300_uid8_T0_copy12_c2 :  std_logic_vector(14 downto 0);
signal bh9_w0_0_c2 :  std_logic;
signal bh9_w1_0_c2 :  std_logic;
signal bh9_w2_0_c2 :  std_logic;
signal bh9_w3_0_c2 :  std_logic;
signal bh9_w4_0_c2 :  std_logic;
signal bh9_w5_0_c2 :  std_logic;
signal bh9_w6_0_c2 :  std_logic;
signal bh9_w7_0_c2 :  std_logic;
signal bh9_w8_0_c2 :  std_logic;
signal bh9_w9_0_c2 :  std_logic;
signal bh9_w10_0_c2 :  std_logic;
signal bh9_w11_0_c2 :  std_logic;
signal bh9_w12_0_c2 :  std_logic;
signal bh9_w13_0_c2 :  std_logic;
signal bh9_w14_0_c2 :  std_logic;
signal FixRealKCM_Freq300_uid8_A1_c2 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq300_uid8_T1_c2 :  std_logic_vector(9 downto 0);
signal FixRealKCM_Freq300_uid8_T1_copy15_c2 :  std_logic_vector(9 downto 0);
signal bh9_w0_1_c2 :  std_logic;
signal bh9_w1_1_c2 :  std_logic;
signal bh9_w2_1_c2 :  std_logic;
signal bh9_w3_1_c2 :  std_logic;
signal bh9_w4_1_c2 :  std_logic;
signal bh9_w5_1_c2 :  std_logic;
signal bh9_w6_1_c2 :  std_logic;
signal bh9_w7_1_c2 :  std_logic;
signal bh9_w8_1_c2 :  std_logic;
signal bh9_w9_1_c2 :  std_logic;
signal FixRealKCM_Freq300_uid8_A2_c2 :  std_logic_vector(2 downto 0);
signal FixRealKCM_Freq300_uid8_T2_c2 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq300_uid8_T2_copy18_c2 :  std_logic_vector(4 downto 0);
signal bh9_w0_2_c2 :  std_logic;
signal bh9_w1_2_c2 :  std_logic;
signal bh9_w2_2_c2 :  std_logic;
signal bh9_w3_2_c2 :  std_logic;
signal bh9_w4_2_c2 :  std_logic;
signal Compressor_23_3_Freq300_uid21_bh9_uid22_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid22_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid22_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh9_w0_3_c2 :  std_logic;
signal bh9_w1_3_c2 :  std_logic;
signal bh9_w2_3_c2 :  std_logic;
signal Compressor_23_3_Freq300_uid21_bh9_uid22_Out0_copy23_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid24_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid24_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid24_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh9_w2_4_c2 :  std_logic;
signal bh9_w3_3_c2 :  std_logic;
signal bh9_w4_3_c2 :  std_logic;
signal Compressor_23_3_Freq300_uid21_bh9_uid24_Out0_copy25_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid26_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid26_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid26_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh9_w4_4_c2 :  std_logic;
signal bh9_w5_2_c2 :  std_logic;
signal bh9_w6_2_c2 :  std_logic;
signal Compressor_23_3_Freq300_uid21_bh9_uid26_Out0_copy27_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid28_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid28_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid28_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh9_w6_3_c2 :  std_logic;
signal bh9_w7_2_c2 :  std_logic;
signal bh9_w8_2_c2 :  std_logic;
signal Compressor_23_3_Freq300_uid21_bh9_uid28_Out0_copy29_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid30_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid30_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid21_bh9_uid30_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh9_w8_3_c2 :  std_logic;
signal bh9_w9_2_c2 :  std_logic;
signal bh9_w10_1_c2 :  std_logic;
signal Compressor_23_3_Freq300_uid21_bh9_uid30_Out0_copy31_c2 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh9_0_c2 :  std_logic_vector(0 downto 0);
signal bitheapFinalAdd_bh9_In0_c2 :  std_logic_vector(14 downto 0);
signal bitheapFinalAdd_bh9_In1_c2 :  std_logic_vector(14 downto 0);
signal bitheapFinalAdd_bh9_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh9_Out_c2 :  std_logic_vector(14 downto 0);
signal bitheapResult_bh9_c2 :  std_logic_vector(14 downto 0);
signal OutRes_c2 :  std_logic_vector(14 downto 0);
begin
-- This operator multiplies by 1/log(2)
   FixRealKCM_Freq300_uid8_A0_c2 <= X(12 downto 8);-- input address  m=9  l=5
   FixRealKCM_Freq300_uid8_Table0: FixRealKCM_Freq300_uid8_T0_Freq300_uid11
      port map ( X => FixRealKCM_Freq300_uid8_A0_c2,
                 Y => FixRealKCM_Freq300_uid8_T0_copy12_c2);
   FixRealKCM_Freq300_uid8_T0_c2 <= FixRealKCM_Freq300_uid8_T0_copy12_c2; -- output copy to hold a pipeline register if needed
   bh9_w0_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(0);
   bh9_w1_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(1);
   bh9_w2_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(2);
   bh9_w3_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(3);
   bh9_w4_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(4);
   bh9_w5_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(5);
   bh9_w6_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(6);
   bh9_w7_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(7);
   bh9_w8_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(8);
   bh9_w9_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(9);
   bh9_w10_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(10);
   bh9_w11_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(11);
   bh9_w12_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(12);
   bh9_w13_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(13);
   bh9_w14_0_c2 <= FixRealKCM_Freq300_uid8_T0_c2(14);
   FixRealKCM_Freq300_uid8_A1_c2 <= X(7 downto 3);-- input address  m=4  l=0
   FixRealKCM_Freq300_uid8_Table1: FixRealKCM_Freq300_uid8_T1_Freq300_uid14
      port map ( X => FixRealKCM_Freq300_uid8_A1_c2,
                 Y => FixRealKCM_Freq300_uid8_T1_copy15_c2);
   FixRealKCM_Freq300_uid8_T1_c2 <= FixRealKCM_Freq300_uid8_T1_copy15_c2; -- output copy to hold a pipeline register if needed
   bh9_w0_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(0);
   bh9_w1_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(1);
   bh9_w2_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(2);
   bh9_w3_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(3);
   bh9_w4_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(4);
   bh9_w5_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(5);
   bh9_w6_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(6);
   bh9_w7_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(7);
   bh9_w8_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(8);
   bh9_w9_1_c2 <= FixRealKCM_Freq300_uid8_T1_c2(9);
   FixRealKCM_Freq300_uid8_A2_c2 <= X(2 downto 0);-- input address  m=-1  l=-3
   FixRealKCM_Freq300_uid8_Table2: FixRealKCM_Freq300_uid8_T2_Freq300_uid17
      port map ( X => FixRealKCM_Freq300_uid8_A2_c2,
                 Y => FixRealKCM_Freq300_uid8_T2_copy18_c2);
   FixRealKCM_Freq300_uid8_T2_c2 <= FixRealKCM_Freq300_uid8_T2_copy18_c2; -- output copy to hold a pipeline register if needed
   bh9_w0_2_c2 <= FixRealKCM_Freq300_uid8_T2_c2(0);
   bh9_w1_2_c2 <= FixRealKCM_Freq300_uid8_T2_c2(1);
   bh9_w2_2_c2 <= FixRealKCM_Freq300_uid8_T2_c2(2);
   bh9_w3_2_c2 <= FixRealKCM_Freq300_uid8_T2_c2(3);
   bh9_w4_2_c2 <= FixRealKCM_Freq300_uid8_T2_c2(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq300_uid21_bh9_uid22_In0_c2 <= "" & bh9_w0_2_c2 & bh9_w0_1_c2 & bh9_w0_0_c2;
   Compressor_23_3_Freq300_uid21_bh9_uid22_In1_c2 <= "" & bh9_w1_2_c2 & bh9_w1_1_c2;
   bh9_w0_3_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid22_Out0_c2(0);
   bh9_w1_3_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid22_Out0_c2(1);
   bh9_w2_3_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid22_Out0_c2(2);
   Compressor_23_3_Freq300_uid21_uid22: Compressor_23_3_Freq300_uid21
      port map ( X0 => Compressor_23_3_Freq300_uid21_bh9_uid22_In0_c2,
                 X1 => Compressor_23_3_Freq300_uid21_bh9_uid22_In1_c2,
                 R => Compressor_23_3_Freq300_uid21_bh9_uid22_Out0_copy23_c2);
   Compressor_23_3_Freq300_uid21_bh9_uid22_Out0_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid22_Out0_copy23_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid21_bh9_uid24_In0_c2 <= "" & bh9_w2_2_c2 & bh9_w2_1_c2 & bh9_w2_0_c2;
   Compressor_23_3_Freq300_uid21_bh9_uid24_In1_c2 <= "" & bh9_w3_2_c2 & bh9_w3_1_c2;
   bh9_w2_4_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid24_Out0_c2(0);
   bh9_w3_3_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid24_Out0_c2(1);
   bh9_w4_3_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid24_Out0_c2(2);
   Compressor_23_3_Freq300_uid21_uid24: Compressor_23_3_Freq300_uid21
      port map ( X0 => Compressor_23_3_Freq300_uid21_bh9_uid24_In0_c2,
                 X1 => Compressor_23_3_Freq300_uid21_bh9_uid24_In1_c2,
                 R => Compressor_23_3_Freq300_uid21_bh9_uid24_Out0_copy25_c2);
   Compressor_23_3_Freq300_uid21_bh9_uid24_Out0_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid24_Out0_copy25_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid21_bh9_uid26_In0_c2 <= "" & bh9_w4_2_c2 & bh9_w4_1_c2 & bh9_w4_0_c2;
   Compressor_23_3_Freq300_uid21_bh9_uid26_In1_c2 <= "" & bh9_w5_1_c2 & bh9_w5_0_c2;
   bh9_w4_4_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid26_Out0_c2(0);
   bh9_w5_2_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid26_Out0_c2(1);
   bh9_w6_2_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid26_Out0_c2(2);
   Compressor_23_3_Freq300_uid21_uid26: Compressor_23_3_Freq300_uid21
      port map ( X0 => Compressor_23_3_Freq300_uid21_bh9_uid26_In0_c2,
                 X1 => Compressor_23_3_Freq300_uid21_bh9_uid26_In1_c2,
                 R => Compressor_23_3_Freq300_uid21_bh9_uid26_Out0_copy27_c2);
   Compressor_23_3_Freq300_uid21_bh9_uid26_Out0_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid26_Out0_copy27_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid21_bh9_uid28_In0_c2 <= "" & bh9_w6_1_c2 & bh9_w6_0_c2 & "0";
   Compressor_23_3_Freq300_uid21_bh9_uid28_In1_c2 <= "" & bh9_w7_1_c2 & bh9_w7_0_c2;
   bh9_w6_3_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid28_Out0_c2(0);
   bh9_w7_2_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid28_Out0_c2(1);
   bh9_w8_2_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid28_Out0_c2(2);
   Compressor_23_3_Freq300_uid21_uid28: Compressor_23_3_Freq300_uid21
      port map ( X0 => Compressor_23_3_Freq300_uid21_bh9_uid28_In0_c2,
                 X1 => Compressor_23_3_Freq300_uid21_bh9_uid28_In1_c2,
                 R => Compressor_23_3_Freq300_uid21_bh9_uid28_Out0_copy29_c2);
   Compressor_23_3_Freq300_uid21_bh9_uid28_Out0_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid28_Out0_copy29_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid21_bh9_uid30_In0_c2 <= "" & bh9_w8_1_c2 & bh9_w8_0_c2 & "0";
   Compressor_23_3_Freq300_uid21_bh9_uid30_In1_c2 <= "" & bh9_w9_1_c2 & bh9_w9_0_c2;
   bh9_w8_3_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid30_Out0_c2(0);
   bh9_w9_2_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid30_Out0_c2(1);
   bh9_w10_1_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid30_Out0_c2(2);
   Compressor_23_3_Freq300_uid21_uid30: Compressor_23_3_Freq300_uid21
      port map ( X0 => Compressor_23_3_Freq300_uid21_bh9_uid30_In0_c2,
                 X1 => Compressor_23_3_Freq300_uid21_bh9_uid30_In1_c2,
                 R => Compressor_23_3_Freq300_uid21_bh9_uid30_Out0_copy31_c2);
   Compressor_23_3_Freq300_uid21_bh9_uid30_Out0_c2 <= Compressor_23_3_Freq300_uid21_bh9_uid30_Out0_copy31_c2; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh9_0_c2(0) <= bh9_w0_3_c2;

   bitheapFinalAdd_bh9_In0_c2 <= "0" & bh9_w14_0_c2 & bh9_w13_0_c2 & bh9_w12_0_c2 & bh9_w11_0_c2 & bh9_w10_0_c2 & bh9_w9_2_c2 & bh9_w8_3_c2 & bh9_w7_2_c2 & bh9_w6_3_c2 & bh9_w5_2_c2 & bh9_w4_4_c2 & bh9_w3_0_c2 & bh9_w2_4_c2 & bh9_w1_0_c2;
   bitheapFinalAdd_bh9_In1_c2 <= "0" & "0" & "0" & "0" & "0" & bh9_w10_1_c2 & "0" & bh9_w8_2_c2 & "0" & bh9_w6_2_c2 & "0" & bh9_w4_3_c2 & bh9_w3_3_c2 & bh9_w2_3_c2 & bh9_w1_3_c2;
   bitheapFinalAdd_bh9_Cin_c0 <= '0';

   bitheapFinalAdd_bh9: IntAdder_15_Freq300_uid33
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 Cin => bitheapFinalAdd_bh9_Cin_c0,
                 X => bitheapFinalAdd_bh9_In0_c2,
                 Y => bitheapFinalAdd_bh9_In1_c2,
                 R => bitheapFinalAdd_bh9_Out_c2);
   bitheapResult_bh9_c2 <= bitheapFinalAdd_bh9_Out_c2(13 downto 0) & tmp_bitheapResult_bh9_0_c2;
   OutRes_c2 <= bitheapResult_bh9_c2(14 downto 0);
   R <= OutRes_c2(14 downto 4);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_68_Freq300_uid45
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_68_Freq300_uid45 is
    port (clk, ce_1, ce_2, ce_3 : in std_logic;
          X : in  std_logic_vector(67 downto 0);
          Y : in  std_logic_vector(67 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(67 downto 0)   );
end entity;

architecture arch of IntAdder_68_Freq300_uid45 is
signal Rtmp_c3 :  std_logic_vector(67 downto 0);
signal X_c3 :  std_logic_vector(67 downto 0);
signal Y_c3 :  std_logic_vector(67 downto 0);
signal Cin_c1, Cin_c2, Cin_c3 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               X_c3 <= X;
               Y_c3 <= Y;
               Cin_c3 <= Cin_c2;
            end if;
         end if;
      end process;
   Rtmp_c3 <= X_c3 + Y_c3 + Cin_c3;
   R <= Rtmp_c3;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq300_uid35
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq300_uid35 is
    port (clk, ce_3 : in std_logic;
          X : in  std_logic_vector(10 downto 0);
          R : out  std_logic_vector(66 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq300_uid35 is
   component FixRealKCM_Freq300_uid35_T0_Freq300_uid38 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(66 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid35_T1_Freq300_uid41 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(61 downto 0)   );
   end component;

   component IntAdder_68_Freq300_uid45 is
      port ( clk, ce_1, ce_2, ce_3 : in std_logic;
             X : in  std_logic_vector(67 downto 0);
             Y : in  std_logic_vector(67 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(67 downto 0)   );
   end component;

signal FixRealKCM_Freq300_uid35_A0_c2 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq300_uid35_T0_c2 :  std_logic_vector(66 downto 0);
signal FixRealKCM_Freq300_uid35_T0_copy39_c2 :  std_logic_vector(66 downto 0);
signal bh36_w0_0_c2 :  std_logic;
signal bh36_w1_0_c2 :  std_logic;
signal bh36_w2_0_c2 :  std_logic;
signal bh36_w3_0_c2 :  std_logic;
signal bh36_w4_0_c2 :  std_logic;
signal bh36_w5_0_c2 :  std_logic;
signal bh36_w6_0_c2 :  std_logic;
signal bh36_w7_0_c2 :  std_logic;
signal bh36_w8_0_c2 :  std_logic;
signal bh36_w9_0_c2 :  std_logic;
signal bh36_w10_0_c2 :  std_logic;
signal bh36_w11_0_c2 :  std_logic;
signal bh36_w12_0_c2 :  std_logic;
signal bh36_w13_0_c2 :  std_logic;
signal bh36_w14_0_c2 :  std_logic;
signal bh36_w15_0_c2 :  std_logic;
signal bh36_w16_0_c2 :  std_logic;
signal bh36_w17_0_c2 :  std_logic;
signal bh36_w18_0_c2 :  std_logic;
signal bh36_w19_0_c2 :  std_logic;
signal bh36_w20_0_c2 :  std_logic;
signal bh36_w21_0_c2 :  std_logic;
signal bh36_w22_0_c2 :  std_logic;
signal bh36_w23_0_c2 :  std_logic;
signal bh36_w24_0_c2 :  std_logic;
signal bh36_w25_0_c2 :  std_logic;
signal bh36_w26_0_c2 :  std_logic;
signal bh36_w27_0_c2 :  std_logic;
signal bh36_w28_0_c2 :  std_logic;
signal bh36_w29_0_c2 :  std_logic;
signal bh36_w30_0_c2 :  std_logic;
signal bh36_w31_0_c2 :  std_logic;
signal bh36_w32_0_c2 :  std_logic;
signal bh36_w33_0_c2 :  std_logic;
signal bh36_w34_0_c2 :  std_logic;
signal bh36_w35_0_c2 :  std_logic;
signal bh36_w36_0_c2 :  std_logic;
signal bh36_w37_0_c2 :  std_logic;
signal bh36_w38_0_c2 :  std_logic;
signal bh36_w39_0_c2 :  std_logic;
signal bh36_w40_0_c2 :  std_logic;
signal bh36_w41_0_c2 :  std_logic;
signal bh36_w42_0_c2 :  std_logic;
signal bh36_w43_0_c2 :  std_logic;
signal bh36_w44_0_c2 :  std_logic;
signal bh36_w45_0_c2 :  std_logic;
signal bh36_w46_0_c2 :  std_logic;
signal bh36_w47_0_c2 :  std_logic;
signal bh36_w48_0_c2 :  std_logic;
signal bh36_w49_0_c2 :  std_logic;
signal bh36_w50_0_c2 :  std_logic;
signal bh36_w51_0_c2 :  std_logic;
signal bh36_w52_0_c2 :  std_logic;
signal bh36_w53_0_c2 :  std_logic;
signal bh36_w54_0_c2 :  std_logic;
signal bh36_w55_0_c2 :  std_logic;
signal bh36_w56_0_c2 :  std_logic;
signal bh36_w57_0_c2 :  std_logic;
signal bh36_w58_0_c2 :  std_logic;
signal bh36_w59_0_c2 :  std_logic;
signal bh36_w60_0_c2 :  std_logic;
signal bh36_w61_0_c2 :  std_logic;
signal bh36_w62_0_c2 :  std_logic;
signal bh36_w63_0_c2 :  std_logic;
signal bh36_w64_0_c2 :  std_logic;
signal bh36_w65_0_c2 :  std_logic;
signal bh36_w66_0_c2 :  std_logic;
signal FixRealKCM_Freq300_uid35_A1_c2 :  std_logic_vector(5 downto 0);
signal FixRealKCM_Freq300_uid35_T1_c2 :  std_logic_vector(61 downto 0);
signal FixRealKCM_Freq300_uid35_T1_copy42_c2 :  std_logic_vector(61 downto 0);
signal bh36_w0_1_c2 :  std_logic;
signal bh36_w1_1_c2 :  std_logic;
signal bh36_w2_1_c2 :  std_logic;
signal bh36_w3_1_c2 :  std_logic;
signal bh36_w4_1_c2 :  std_logic;
signal bh36_w5_1_c2 :  std_logic;
signal bh36_w6_1_c2 :  std_logic;
signal bh36_w7_1_c2 :  std_logic;
signal bh36_w8_1_c2 :  std_logic;
signal bh36_w9_1_c2 :  std_logic;
signal bh36_w10_1_c2 :  std_logic;
signal bh36_w11_1_c2 :  std_logic;
signal bh36_w12_1_c2 :  std_logic;
signal bh36_w13_1_c2 :  std_logic;
signal bh36_w14_1_c2 :  std_logic;
signal bh36_w15_1_c2 :  std_logic;
signal bh36_w16_1_c2 :  std_logic;
signal bh36_w17_1_c2 :  std_logic;
signal bh36_w18_1_c2 :  std_logic;
signal bh36_w19_1_c2 :  std_logic;
signal bh36_w20_1_c2 :  std_logic;
signal bh36_w21_1_c2 :  std_logic;
signal bh36_w22_1_c2 :  std_logic;
signal bh36_w23_1_c2 :  std_logic;
signal bh36_w24_1_c2 :  std_logic;
signal bh36_w25_1_c2 :  std_logic;
signal bh36_w26_1_c2 :  std_logic;
signal bh36_w27_1_c2 :  std_logic;
signal bh36_w28_1_c2 :  std_logic;
signal bh36_w29_1_c2 :  std_logic;
signal bh36_w30_1_c2 :  std_logic;
signal bh36_w31_1_c2 :  std_logic;
signal bh36_w32_1_c2 :  std_logic;
signal bh36_w33_1_c2 :  std_logic;
signal bh36_w34_1_c2 :  std_logic;
signal bh36_w35_1_c2 :  std_logic;
signal bh36_w36_1_c2 :  std_logic;
signal bh36_w37_1_c2 :  std_logic;
signal bh36_w38_1_c2 :  std_logic;
signal bh36_w39_1_c2 :  std_logic;
signal bh36_w40_1_c2 :  std_logic;
signal bh36_w41_1_c2 :  std_logic;
signal bh36_w42_1_c2 :  std_logic;
signal bh36_w43_1_c2 :  std_logic;
signal bh36_w44_1_c2 :  std_logic;
signal bh36_w45_1_c2 :  std_logic;
signal bh36_w46_1_c2 :  std_logic;
signal bh36_w47_1_c2 :  std_logic;
signal bh36_w48_1_c2 :  std_logic;
signal bh36_w49_1_c2 :  std_logic;
signal bh36_w50_1_c2 :  std_logic;
signal bh36_w51_1_c2 :  std_logic;
signal bh36_w52_1_c2 :  std_logic;
signal bh36_w53_1_c2 :  std_logic;
signal bh36_w54_1_c2 :  std_logic;
signal bh36_w55_1_c2 :  std_logic;
signal bh36_w56_1_c2 :  std_logic;
signal bh36_w57_1_c2 :  std_logic;
signal bh36_w58_1_c2 :  std_logic;
signal bh36_w59_1_c2 :  std_logic;
signal bh36_w60_1_c2 :  std_logic;
signal bh36_w61_1_c2 :  std_logic;
signal bitheapFinalAdd_bh36_In0_c2 :  std_logic_vector(67 downto 0);
signal bitheapFinalAdd_bh36_In1_c2 :  std_logic_vector(67 downto 0);
signal bitheapFinalAdd_bh36_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh36_Out_c3 :  std_logic_vector(67 downto 0);
signal bitheapResult_bh36_c3 :  std_logic_vector(66 downto 0);
signal OutRes_c3 :  std_logic_vector(66 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_3 = '1' then
            end if;
         end if;
      end process;
-- This operator multiplies by log(2)
   FixRealKCM_Freq300_uid35_A0_c2 <= X(10 downto 6);-- input address  m=10  l=6
   FixRealKCM_Freq300_uid35_Table0: FixRealKCM_Freq300_uid35_T0_Freq300_uid38
      port map ( X => FixRealKCM_Freq300_uid35_A0_c2,
                 Y => FixRealKCM_Freq300_uid35_T0_copy39_c2);
   FixRealKCM_Freq300_uid35_T0_c2 <= FixRealKCM_Freq300_uid35_T0_copy39_c2; -- output copy to hold a pipeline register if needed
   bh36_w0_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(0);
   bh36_w1_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(1);
   bh36_w2_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(2);
   bh36_w3_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(3);
   bh36_w4_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(4);
   bh36_w5_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(5);
   bh36_w6_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(6);
   bh36_w7_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(7);
   bh36_w8_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(8);
   bh36_w9_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(9);
   bh36_w10_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(10);
   bh36_w11_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(11);
   bh36_w12_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(12);
   bh36_w13_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(13);
   bh36_w14_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(14);
   bh36_w15_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(15);
   bh36_w16_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(16);
   bh36_w17_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(17);
   bh36_w18_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(18);
   bh36_w19_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(19);
   bh36_w20_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(20);
   bh36_w21_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(21);
   bh36_w22_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(22);
   bh36_w23_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(23);
   bh36_w24_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(24);
   bh36_w25_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(25);
   bh36_w26_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(26);
   bh36_w27_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(27);
   bh36_w28_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(28);
   bh36_w29_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(29);
   bh36_w30_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(30);
   bh36_w31_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(31);
   bh36_w32_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(32);
   bh36_w33_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(33);
   bh36_w34_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(34);
   bh36_w35_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(35);
   bh36_w36_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(36);
   bh36_w37_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(37);
   bh36_w38_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(38);
   bh36_w39_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(39);
   bh36_w40_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(40);
   bh36_w41_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(41);
   bh36_w42_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(42);
   bh36_w43_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(43);
   bh36_w44_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(44);
   bh36_w45_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(45);
   bh36_w46_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(46);
   bh36_w47_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(47);
   bh36_w48_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(48);
   bh36_w49_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(49);
   bh36_w50_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(50);
   bh36_w51_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(51);
   bh36_w52_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(52);
   bh36_w53_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(53);
   bh36_w54_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(54);
   bh36_w55_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(55);
   bh36_w56_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(56);
   bh36_w57_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(57);
   bh36_w58_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(58);
   bh36_w59_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(59);
   bh36_w60_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(60);
   bh36_w61_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(61);
   bh36_w62_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(62);
   bh36_w63_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(63);
   bh36_w64_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(64);
   bh36_w65_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(65);
   bh36_w66_0_c2 <= FixRealKCM_Freq300_uid35_T0_c2(66);
   FixRealKCM_Freq300_uid35_A1_c2 <= X(5 downto 0);-- input address  m=5  l=0
   FixRealKCM_Freq300_uid35_Table1: FixRealKCM_Freq300_uid35_T1_Freq300_uid41
      port map ( X => FixRealKCM_Freq300_uid35_A1_c2,
                 Y => FixRealKCM_Freq300_uid35_T1_copy42_c2);
   FixRealKCM_Freq300_uid35_T1_c2 <= FixRealKCM_Freq300_uid35_T1_copy42_c2; -- output copy to hold a pipeline register if needed
   bh36_w0_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(0);
   bh36_w1_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(1);
   bh36_w2_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(2);
   bh36_w3_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(3);
   bh36_w4_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(4);
   bh36_w5_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(5);
   bh36_w6_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(6);
   bh36_w7_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(7);
   bh36_w8_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(8);
   bh36_w9_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(9);
   bh36_w10_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(10);
   bh36_w11_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(11);
   bh36_w12_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(12);
   bh36_w13_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(13);
   bh36_w14_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(14);
   bh36_w15_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(15);
   bh36_w16_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(16);
   bh36_w17_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(17);
   bh36_w18_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(18);
   bh36_w19_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(19);
   bh36_w20_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(20);
   bh36_w21_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(21);
   bh36_w22_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(22);
   bh36_w23_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(23);
   bh36_w24_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(24);
   bh36_w25_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(25);
   bh36_w26_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(26);
   bh36_w27_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(27);
   bh36_w28_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(28);
   bh36_w29_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(29);
   bh36_w30_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(30);
   bh36_w31_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(31);
   bh36_w32_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(32);
   bh36_w33_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(33);
   bh36_w34_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(34);
   bh36_w35_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(35);
   bh36_w36_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(36);
   bh36_w37_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(37);
   bh36_w38_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(38);
   bh36_w39_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(39);
   bh36_w40_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(40);
   bh36_w41_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(41);
   bh36_w42_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(42);
   bh36_w43_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(43);
   bh36_w44_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(44);
   bh36_w45_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(45);
   bh36_w46_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(46);
   bh36_w47_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(47);
   bh36_w48_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(48);
   bh36_w49_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(49);
   bh36_w50_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(50);
   bh36_w51_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(51);
   bh36_w52_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(52);
   bh36_w53_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(53);
   bh36_w54_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(54);
   bh36_w55_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(55);
   bh36_w56_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(56);
   bh36_w57_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(57);
   bh36_w58_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(58);
   bh36_w59_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(59);
   bh36_w60_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(60);
   bh36_w61_1_c2 <= FixRealKCM_Freq300_uid35_T1_c2(61);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh36_In0_c2 <= "0" & bh36_w66_0_c2 & bh36_w65_0_c2 & bh36_w64_0_c2 & bh36_w63_0_c2 & bh36_w62_0_c2 & bh36_w61_0_c2 & bh36_w60_0_c2 & bh36_w59_0_c2 & bh36_w58_0_c2 & bh36_w57_0_c2 & bh36_w56_0_c2 & bh36_w55_0_c2 & bh36_w54_0_c2 & bh36_w53_0_c2 & bh36_w52_0_c2 & bh36_w51_0_c2 & bh36_w50_0_c2 & bh36_w49_0_c2 & bh36_w48_0_c2 & bh36_w47_0_c2 & bh36_w46_0_c2 & bh36_w45_0_c2 & bh36_w44_0_c2 & bh36_w43_0_c2 & bh36_w42_0_c2 & bh36_w41_0_c2 & bh36_w40_0_c2 & bh36_w39_0_c2 & bh36_w38_0_c2 & bh36_w37_0_c2 & bh36_w36_0_c2 & bh36_w35_0_c2 & bh36_w34_0_c2 & bh36_w33_0_c2 & bh36_w32_0_c2 & bh36_w31_0_c2 & bh36_w30_0_c2 & bh36_w29_0_c2 & bh36_w28_0_c2 & bh36_w27_0_c2 & bh36_w26_0_c2 & bh36_w25_0_c2 & bh36_w24_0_c2 & bh36_w23_0_c2 & bh36_w22_0_c2 & bh36_w21_0_c2 & bh36_w20_0_c2 & bh36_w19_0_c2 & bh36_w18_0_c2 & bh36_w17_0_c2 & bh36_w16_0_c2 & bh36_w15_0_c2 & bh36_w14_0_c2 & bh36_w13_0_c2 & bh36_w12_0_c2 & bh36_w11_0_c2 & bh36_w10_0_c2 & bh36_w9_0_c2 & bh36_w8_0_c2 & bh36_w7_0_c2 & bh36_w6_0_c2 & bh36_w5_0_c2 & bh36_w4_0_c2 & bh36_w3_0_c2 & bh36_w2_0_c2 & bh36_w1_0_c2 & bh36_w0_0_c2;
   bitheapFinalAdd_bh36_In1_c2 <= "0" & "0" & "0" & "0" & "0" & "0" & bh36_w61_1_c2 & bh36_w60_1_c2 & bh36_w59_1_c2 & bh36_w58_1_c2 & bh36_w57_1_c2 & bh36_w56_1_c2 & bh36_w55_1_c2 & bh36_w54_1_c2 & bh36_w53_1_c2 & bh36_w52_1_c2 & bh36_w51_1_c2 & bh36_w50_1_c2 & bh36_w49_1_c2 & bh36_w48_1_c2 & bh36_w47_1_c2 & bh36_w46_1_c2 & bh36_w45_1_c2 & bh36_w44_1_c2 & bh36_w43_1_c2 & bh36_w42_1_c2 & bh36_w41_1_c2 & bh36_w40_1_c2 & bh36_w39_1_c2 & bh36_w38_1_c2 & bh36_w37_1_c2 & bh36_w36_1_c2 & bh36_w35_1_c2 & bh36_w34_1_c2 & bh36_w33_1_c2 & bh36_w32_1_c2 & bh36_w31_1_c2 & bh36_w30_1_c2 & bh36_w29_1_c2 & bh36_w28_1_c2 & bh36_w27_1_c2 & bh36_w26_1_c2 & bh36_w25_1_c2 & bh36_w24_1_c2 & bh36_w23_1_c2 & bh36_w22_1_c2 & bh36_w21_1_c2 & bh36_w20_1_c2 & bh36_w19_1_c2 & bh36_w18_1_c2 & bh36_w17_1_c2 & bh36_w16_1_c2 & bh36_w15_1_c2 & bh36_w14_1_c2 & bh36_w13_1_c2 & bh36_w12_1_c2 & bh36_w11_1_c2 & bh36_w10_1_c2 & bh36_w9_1_c2 & bh36_w8_1_c2 & bh36_w7_1_c2 & bh36_w6_1_c2 & bh36_w5_1_c2 & bh36_w4_1_c2 & bh36_w3_1_c2 & bh36_w2_1_c2 & bh36_w1_1_c2 & bh36_w0_1_c2;
   bitheapFinalAdd_bh36_Cin_c0 <= '0';

   bitheapFinalAdd_bh36: IntAdder_68_Freq300_uid45
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 Cin => bitheapFinalAdd_bh36_Cin_c0,
                 X => bitheapFinalAdd_bh36_In0_c2,
                 Y => bitheapFinalAdd_bh36_In1_c2,
                 R => bitheapFinalAdd_bh36_Out_c3);
   bitheapResult_bh36_c3 <= bitheapFinalAdd_bh36_Out_c3(66 downto 0);
   OutRes_c3 <= bitheapResult_bh36_c3(66 downto 0);
   R <= OutRes_c3(66 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_56_Freq300_uid48
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_56_Freq300_uid48 is
    port (clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntAdder_56_Freq300_uid48 is
signal Rtmp_c4 :  std_logic_vector(55 downto 0);
signal X_c3, X_c4 :  std_logic_vector(55 downto 0);
signal Y_c4 :  std_logic_vector(55 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               X_c3 <= X;
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               X_c4 <= X_c3;
               Y_c4 <= Y;
               Cin_c4 <= Cin_c3;
            end if;
         end if;
      end process;
   Rtmp_c4 <= X_c4 + Y_c4 + Cin_c4;
   R <= Rtmp_c4;
end architecture;

--------------------------------------------------------------------------------
--              compressedTable_Freq300_uid52_diff_Freq300_uid57
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity compressedTable_Freq300_uid52_diff_Freq300_uid57 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(49 downto 0)   );
end entity;

architecture arch of compressedTable_Freq300_uid52_diff_Freq300_uid57 is
signal Y0_c4 :  std_logic_vector(49 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "block";
signal Y1_c4 :  std_logic_vector(49 downto 0);
begin
   with X  select  Y0_c4 <= 
      "00000000000000000000000000000000000000000000000000" when "0000000000",
      "00010000000000100000000000101010101011010101010110" when "0000000001",
      "00100000000010000000000101010101100000000000010001" when "0000000010",
      "00110000000100100000010010000000110110000010000010" when "0000000011",
      "01000000001000000000101010101101010101011101111000" when "0000000100",
      "01010000001100100001010011011011110110011010000100" when "0000000101",
      "01100000010010000010010000001101100001000000110111" when "0000000110",
      "01110000011000100011100101000011101101100001100011" when "0000000111",
      "00000000100000000101010110000000000100010001011011" when "0000001000",
      "00010000101000100111100111000100011101101100110011" when "0000001001",
      "00100000110010001010011100010011000010011000000010" when "0000001010",
      "00110000111100101101111001101110001011000000100000" when "0000001011",
      "01000001001000010010000011011000100000011101101010" when "0000001100",
      "01010001010100110110111101010100111011110010000000" when "0000001101",
      "01100001100010011100101011100110100110001100000110" when "0000001110",
      "01110001110001000011010010010000111001000111100111" when "0000001111",
      "00000010000000101010110101010111011110001110010001" when "0000010000",
      "00010010010001010011011000111110001111011000111101" when "0000010001",
      "00100010100010111101000001001001010110110000101001" when "0000010010",
      "00110010110101100111110001111101001110101111011110" when "0000010011",
      "01000011001001010011101111011110100010000001101110" when "0000010100",
      "01010011011110000000111101110010001011100110110110" when "0000010101",
      "01100011110011101111100000111101010110110010100001" when "0000010110",
      "01110100001010011111011101000101011111001101101000" when "0000010111",
      "00000100100010010000110110010000010000110111010001" when "0000011000",
      "00010100111011000011110000100011101000000101110110" when "0000011001",
      "00100101010100111000010000000101110001100111111111" when "0000011010",
      "00110101101111101110011000111101001010100101101100" when "0000011011",
      "01000110001011100110001111010000100000100001001111" when "0000011100",
      "01010110101000011111110111000110110001011000010011" when "0000011101",
      "01100111000110011011010100100111001011100100111011" when "0000011110",
      "01110111100101011000101011111001001101111110100101" when "0000011111",
      "00001000000101011000000001000100100111111011001010" when "0000100000",
      "00011000100110011001011000010001011001010000000010" when "0000100001",
      "00101001001000011100110101100111110010010011001000" when "0000100010",
      "00111001101011100010011101010000010011111011110101" when "0000100011",
      "01001010001111101010010011010011101111100100001001" when "0000100100",
      "01011010110100110100011011111011000111001001101011" when "0000100101",
      "01101011011011000000111011001111101101001110101010" when "0000100110",
      "01111100000010001111110101011011000100111011000001" when "0000100111",
      "00001100101010100001001110100111000001111101011000" when "0000101000",
      "00011101010011110101001010111101101000101100001000" when "0000101001",
      "00101101111110001011101110101001001110000110011011" when "0000101010",
      "00111110101001100100111101110100010111110101010011" when "0000101011",
      "01001111010110000000111100101001111100001100100111" when "0000101100",
      "01100000000011011111101111010101000010001100001011" when "0000101101",
      "01110000110010000001011010000001000001100000101111" when "0000101110",
      "10000001100001100110000000111001100010100101000100" when "0000101111",
      "00010010010010001101101000001010011110100010111100" when "0000110000",
      "00100011000011111000010011111111111111010100010011" when "0000110001",
      "00110011110110100110001000100110011111100100001011" when "0000110010",
      "01000100101010010111001010001010101010101111110011" when "0000110011",
      "01010101011111001011011100111001011101000111101001" when "0000110100",
      "01100110010101000011000101000000000011110000100000" when "0000110101",
      "01110111001011111110000110101011111100100100011111" when "0000110110",
      "10001000000011111100100110001010110110010100000101" when "0000110111",
      "00011000111100111110100111101010110000100111010001" when "0000111000",
      "00101001110111000100001111011001111011111110100000" when "0000111001",
      "00111010110010001101100001100110111001110011110100" when "0000111010",
      "01001011101110011010100010100000011100011011110101" when "0000111011",
      "01011100101011101011010110010101100111000110110111" when "0000111100",
      "01101101101010000000000001010101101110000001111101" when "0000111101",
      "01111110101001011000100111110000010110010111111101" when "0000111110",
      "10001111101001110101001101110101010110010010100100" when "0000111111",
      "00100000101011010101110111110100110100111011011000" when "0001000000",
      "00110001101101111010101001111111001010011100111110" when "0001000001",
      "01000010110001100011101000100101000000000100000000" when "0001000010",
      "01010011110110010000110111110111010000000000001100" when "0001000011",
      "01100100111100000010011100000111000101100101011100" when "0001000100",
      "01110110000010111000011001100101111101001100111011" when "0001000101",
      "10000111001010110010110100100101100100010110000100" when "0001000110",
      "10011000010011110001110001010111111001100111101111" when "0001000111",
      "00101001011101110101010100001111001100110001001110" when "0001001000",
      "00111010101000111101100001011101111110101011010011" when "0001001001",
      "01001011110101001010011101010111000001011001011001" when "0001001010",
      "01011101000010011100001100001101011000001010100011" when "0001001011",
      "01101110010000110010110010010100010111011010100101" when "0001001100",
      "01111111100000001110010011111111100100110011000110" when "0001001101",
      "10010000110000101110110101100010110111001100100110" when "0001001110",
      "10100010000010010100011011010010010110101111100101" when "0001001111",
      "00110011010100111111001001100010011100110101100100" when "0001010000",
      "01000100101000101111000100100111110100001010001101" when "0001010001",
      "01010101111101100100010000110111011000101100010110" when "0001010010",
      "01100111010011011110110010100110010111101111001010" when "0001010011",
      "01111000101010011110101110001010001111111011001010" when "0001010100",
      "10001010000010100100000111111000110001001111010101" when "0001010101",
      "10011011011011101111000100000111111101000010001100" when "0001010110",
      "10101100110101111111100111001110000110000010111001" when "0001010111",
      "00111110010001010101110101100001110000011010010011" when "0001011000",
      "01001111101101110001110011011001110001101100000101" when "0001011001",
      "01100001001011010011100101001101010000110111110010" when "0001011010",
      "01110010101001111011001111010011100110011001111110" when "0001011011",
      "10000100001001101000110110000100011100001101010000" when "0001011100",
      "10010101101010011100011101110111101101101011011001" when "0001011101",
      "10100111001100010110001011000101100111101110011101" when "0001011110",
      "10111000101111010110000010000110101000110001110101" when "0001011111",
      "00001010010011011100000111010011100000110011010111" when "0001100000",
      "00011011111000101000011111000101010001010100011011" when "0001100001",
      "00101101011110111011001101110101001101011011000101" when "0001100010",
      "00111111000110010100010111111100111001110011000110" when "0001100011",
      "01010000101110110100000001110110001100101111000110" when "0001100100",
      "01100010011000011010001111111011001110001001101001" when "0001100101",
      "01110100000011000111000110100110010111100110010111" when "0001100110",
      "10000101101110111010101010010010010100010010111111" when "0001100111",
      "00010111011011110100111111011010000001001000100011" when "0001101000",
      "00101001001001110110001010011000101100101100011011" when "0001101001",
      "00111010111000111110001111101001110111010001011100" when "0001101010",
      "01001100101001001101010011101001010010111001000000" when "0001101011",
      "01011110011010100011011010110011000011010100001110" when "0001101100",
      "01110000001101000000101001100011011110000100111101" when "0001101101",
      "10000010000000100101000100010111001010011111000000" when "0001101110",
      "10010011110101010000101111101011000001101001001001" when "0001101111",
      "00100101101011000011101111111100001110011110010100" when "0001110000",
      "00110111100001111110001001101000001101101110101010" when "0001110001",
      "01001001011010000000000001001100101110000000101101" when "0001110010",
      "01011011010011001001011011000111101111110010011011" when "0001110011",
      "01101101001101011010011011110111100101011010011010" when "0001110100",
      "01111111001000110011000111111010110011001000111011" when "0001110101",
      "10010001000101010011100011110000001111001001000110" when "0001110110",
      "10100011000010111011110011110111000001100001111100" when "0001110111",
      "00110101000001101011111100101110100100010111100111" when "0001111000",
      "01000111000001100100000010110110100011101100011010" when "0001111001",
      "01011001000010100100001010101110111101100001111100" when "0001111010",
      "01101011000100101100011000111000000001111010010011" when "0001111011",
      "01111101000111111100110001110010010010111001000110" when "0001111100",
      "10001111001100010101011001111110100100100100101010" when "0001111101",
      "10100001010001110110010101111101111101000111001001" when "0001111110",
      "10110011011000011111101010010001110100101111100111" when "0001111111",
      "00000101100000010001011011011011110101110011010000" when "0010000000",
      "00010111101001001011101101111101111100101110011100" when "0010000001",
      "00101001110011001110100110011010011000000101111011" when "0010000010",
      "00111011111110011010001001010011101000100111111000" when "0010000011",
      "01001110001010101110011011001100100001001101001001" when "0010000100",
      "01100000011000001011100000101000000110111010010011" when "0010000101",
      "01110010100110110001011110001001110001000000110000" when "0010000110",
      "10000100110110100000011000010101001001000000000010" when "0010000111",
      "00010111000111011000010011101110001010100110101111" when "0010001000",
      "00101001011001011001010100111001000011110011110101" when "0010001001",
      "00111011101100100011100000011010010100110111101101" when "0010001010",
      "01001110000000110110111010110110110000010101010100" when "0010001011",
      "01100000010110010011101000110011011011000011011000" when "0010001100",
      "01110010101100111001101110110101101100001101011111" when "0010001101",
      "10000101000100101001010001100011001101010101001110" when "0010001110",
      "10010111011101100010010101100001111010010011011000" when "0010001111",
      "00101001110111100100111111011000000001011001000011" when "0010010000",
      "00111100010010110001010011101100000011010000110001" when "0010010001",
      "01001110101111000111010111000100110010111111101110" when "0010010010",
      "01100001001100100111001110001001010110000110110111" when "0010010011",
      "01110011101011010000111101100001000100100100000011" when "0010010100",
      "10000110001011000100101001110011101000110011001101" when "0010010101",
      "10011000101100000010010111101000111111101111100001" when "0010010110",
      "10101011001110001010001011101001011000110100100011" when "0010010111",
      "00111101110001011100001010011101010101111111010111" when "0010011000",
      "01010000010101111000011000101101101011101111110011" when "0010011001",
      "01100010111011011110111011000011100001001001011111" when "0010011010",
      "01110101100010001111110110001000001111110101000111" when "0010011011",
      "10001000001010001011001110100101100100000001100100" when "0010011100",
      "10011010110011010001001001000101011100100101000010" when "0010011101",
      "10101101011101100001101010010010001010111110001111" when "0010011110",
      "11000000001000111100110110110110010011010101100110" when "0010011111",
      "00010010110101100010110011011100101100011110010101" when "0010100000",
      "00100101100011010011100100110000011111110111101100" when "0010100001",
      "00111000010010001111001111011101001001101110000110" when "0010100010",
      "01001011000010010101111000001110011000111100010101" when "0010100011",
      "01011101110011100111100011110000001111001100101100" when "0010100100",
      "01110000100110000100010110101111000000111010001000" when "0010100101",
      "10000011011001101100010101110111010101010001100000" when "0010100110",
      "10010110001110011111100101110110000110010010101101" when "0010100111",
      "00101001000100011110001011011000100000110001110100" when "0010101000",
      "00111011111011101000001011001100000100011000010100" when "0010101001",
      "01001110110011111101101001111110100011100110010000" when "0010101010",
      "01100001101101011110101100011110000011110011011100" when "0010101011",
      "01110100101000001011010111011000111101010000100101" when "0010101100",
      "10000111100100000011101111011101111011001000100000" when "0010101101",
      "10011010100001000111111001011011111011100001010110" when "0010101110",
      "10101101011111010111111010000010001111011101101011" when "0010101111",
      "00000000011110110011110110000000011010111101110000" when "0010110000",
      "00010011011111011011110010000110010101000000101011" when "0010110001",
      "00100110100001001111110011000100000111100101100011" when "0010110010",
      "00111001100100001111111101101010001111101100101110" when "0010110011",
      "01001100101000011100010110101001011101011000111100" when "0010110100",
      "01011111101101110101000010110010110011110000100100" when "0010110101",
      "01110010110100011010000110110111101000111110101101" when "0010110110",
      "10000101111100001011100111101001100110010100100000" when "0010110111",
      "00011001000101001001101001111010101000001010010000" when "0010111000",
      "00101100001111010100010010011100111110000000100110" when "0010111001",
      "00111111011010101011100110000011001010100001110010" when "0010111010",
      "01010010100111001111101001100000000011100010110101" when "0010111011",
      "01100101110101000000100001100110110010000100101011" when "0010111100",
      "01111001000011111110010011001010110010010101011100" when "0010111101",
      "10001100010100001001000010111111110011110001101001" when "0010111110",
      "10011111100101100000110101111001111001000101010100" when "0010111111",
      "00110010111000000101110000101101011000001101010011" when "0011000000",
      "01000110001011110111111000001110111010011000011001" when "0011000001",
      "01011001100000110111010001010011011100001000100100" when "0011000010",
      "01101100110111000100000000110000001101010100001110" when "0011000011",
      "10000000001110011110001011011010110001000111010010" when "0011000100",
      "10010011100111000101110110001000111110000100100010" when "0011000101",
      "10100111000000111011000101110000111110000110110000" when "0011000110",
      "10111010011011111101111111001001001110100001111101" when "0011000111",
      "00001101111000001110100111001000100000000100100101" when "0011001000",
      "00100001010101101101000010100101110110111000101110" when "0011001001",
      "00110100110100011001010110011000101010100101010111" when "0011001010",
      "01001000010100010011100111011000100110001111100010" when "0011001011",
      "01011011110101011011111010011101101000011011100110" when "0011001100",
      "01101111010111110010010100100000000011001110011011" when "0011001101",
      "10000010111011010110111010011000011100001110100111" when "0011001110",
      "10010110100000001001110000111111101100100101110000" when "0011001111",
      "00101010000110001010111101001111000001000001100110" when "0011010000",
      "00111101101101011010100011111111111001110101010011" when "0011010001",
      "01010001010101111000101010001100001010111010101001" when "0011010010",
      "01100100111111100101010100101101111011110011010100" when "0011010011",
      "01111000101010100000101000011111100111101010000000" when "0011010100",
      "10001100010110101010101010011011111101010011110010" when "0011010101",
      "10100000000100000011011111011101111111010001010000" when "0011010110",
      "10110011110010101011001100100001000011101111101111" when "0011010111",
      "00000111100010100001110110100000110100101010101000" when "0011011000",
      "00011011010011100111100010011001001111101100100001" when "0011011001",
      "00101111000101111100010101000110100110010000011111" when "0011011010",
      "01000010111001100000010011100101011101100011010011" when "0011011011",
      "01010110101110010011100010110010101110100100101101" when "0011011100",
      "01101010100100010110000111101011100110001000100101" when "0011011101",
      "01111110011011101000000111001101100100111000010001" when "0011011110",
      "10010010010100001001100110010110011111010011110000" when "0011011111",
      "00100110001101111010101010000100011101110010111011" when "0011100000",
      "00111010001000111011010111010101111100100110110011" when "0011100001",
      "01001110000101001011110011001001101011111010110101" when "0011100010",
      "01100010000010101100000010011110101111110110000010" when "0011100011",
      "01110110000001011100001010010100100000011100011001" when "0011100100",
      "10001010000001011100001111101010101001101111111011" when "0011100101",
      "10011110000010101100010111100001001011110010000111" when "0011100110",
      "10110010000101001100100110111000011010100100111111" when "0011100111",
      "00000110001000111101000010110000111110001100100001" when "0011101000",
      "00011010001101111101110000001011110010101111110001" when "0011101001",
      "00101110010100001110110100001010001000011010001101" when "0011101010",
      "01000010011011110000010011101101100011011100111011" when "0011101011",
      "01010110100100100010010011110111111100001111111010" when "0011101100",
      "01101010101110100100111001101011011111010011010100" when "0011101101",
      "01111110111001111000001010001010101101010000101101" when "0011101110",
      "10010011000110011100001010011000011010111100010010" when "0011101111",
      "00100111010100010000111111010111110001010110001111" when "0011110000",
      "00111011100011010110101110001100001101101011111001" when "0011110001",
      "01001111110011101101011011111001100001011001000101" when "0011110010",
      "01100100000101010101001101100011110010001001010101" when "0011110011",
      "01111000011000001110001000001111011001111001001010" when "0011110100",
      "10001100101100011000010001000001000110110111010101" when "0011110101",
      "10100001000001110011101100111101111011100110001010" when "0011110110",
      "10110101011000100000100001001011001110111100101111" when "0011110111",
      "00001001110000011110110010101110101100001000001110" when "0011111000",
      "00011110001001101110100110101110010010101101000110" when "0011111001",
      "00110010100100010000000010010000010110101000011111" when "0011111010",
      "01000111000000000011001010011011100000010001010111" when "0011111011",
      "01011011011101001000000100010110101100011001111001" when "0011111100",
      "01101111111011011110110101001001001100010000101001" when "0011111101",
      "10000100011011000111100001111010100101100001111100" when "0011111110",
      "10011000111100000010001111110010110010011001000100" when "0011111111",
      "00101101011110001111000011111010000001100001100110" when "0100000000",
      "01000010000001101110000011011000110110001000101100" when "0100000001",
      "01010110100110011111010011011000000111111110010011" when "0100000010",
      "01101011001100100010111001000001000011010110100010" when "0100000011",
      "01111111110011111000111001011101001001001010111011" when "0100000100",
      "10010100011100100001011001110110001110111011101011" when "0100000101",
      "10101001000110011100011111010110011110110000111111" when "0100000110",
      "10111101110001101010001111001000010111011100010110" when "0100000111",
      "00010010011110001010101110010110101100011001110100" when "0100001000",
      "00100111001011111110000010001100100101110001010100" when "0100001001",
      "00111011111011000100001111110101100000010111111001" when "0100001010",
      "01010000101011011101011100011101001101110001000100" when "0100001011",
      "01100101011101001001101101001111110100010000000111" when "0100001100",
      "01111010010000001001000111011001101110111001010101" when "0100001101",
      "10001111000100011011110000000111101101100011011000" when "0100001110",
      "10100011111010000001101100100110110100111000100010" when "0100001111",
      "00111000110000111011000010000100011110011000000001" when "0100010000",
      "01001101101001000111110101101110011000010111010101" when "0100010001",
      "01100010100010101000001100110010100110000011011101" when "0100010010",
      "01110111011101011100001100011111011111100010010100" when "0100010011",
      "10001100011001100011111010000011110001110011111010" when "0100010100",
      "10100001010110111111011010101110011110110011110000" when "0100010101",
      "10110110010101101110110011101110111101011010000111" when "0100010110",
      "11001011010101110010001010010100111001011101010111" when "0100010111",
      "00100000010111001001100011110000010011110011001111" when "0100011000",
      "00110101011001110101000101010001100010010010001111" when "0100011001",
      "01001010011101110100110100001001001111110010110101" when "0100011010",
      "01011111100011001000110101101000011100010000110110" when "0100011011",
      "01110100101001110001001111000000011100101100110001" when "0100011100",
      "10001001110001101110000101100010111011001101000010" when "0100011101",
      "10011110111010111111011110100001110110111111011011" when "0100011110",
      "10110100000101100101011111001111100100011010010001" when "0100011111",
      "00001001010001100000001100111110101100111101110111" when "0100100000",
      "00011110011110101111101101000010001111010101101111" when "0100100001",
      "00110011101101010100000100101101011111011010000011" when "0100100010",
      "01001000111101001101011001010100000110010000110011" when "0100100011",
      "01011110001110011011110000001010000010001111010000" when "0100100100",
      "01110011100000111111001110100011100110111011001111" when "0100100101",
      "10001000110100110111111001110101011101001100011110" when "0100100110",
      "10011110001010000101110111010100100011001101111000" when "0100100111",
      "00110011100000101001001100010110001100011110111011" when "0100101000",
      "01001000111000100001111110010000000001110101000000" when "0100101001",
      "01011110010001110000010010011000000001011100101100" when "0100101010",
      "01110011101100010100001110000100011110111011001000" when "0100101011",
      "10001001001000001101110110101100000011001111010110" when "0100101100",
      "10011110100101011101010001100101101100110011101000" when "0100101101",
      "10110100000100000010100100001000101111011110110010" when "0100101110",
      "11001001100011111101110011101100110100100101100110" when "0100101111",
      "00011111000101001111000101101001111010111100000010" when "0100110000",
      "00110100100111110110011111011000010110110110101111" when "0100110001",
      "01001010001011110100000110010000110010001100001101" when "0100110010",
      "01011111110001000111111111101100001100010110010011" when "0100110011",
      "01110101010111110010010001000011111010010011011110" when "0100110100",
      "10001010111111110010111111110001100110101000001101" when "0100110101",
      "10100000101001001010010001001111010001100000010001" when "0100110110",
      "10110110010011111000001010110111010000110000001000" when "0100110111",
      "00001011111111111100110010000100001111110110010101" when "0100111000",
      "00100001101101011000001100010001001111111100110010" when "0100111001",
      "00110111011100001010011110111001100111111010001001" when "0100111010",
      "01001101001100010011101111011001000100010011001100" when "0100111011",
      "01100010111101110100000011001011100111011100001001" when "0100111100",
      "01111000110000101011011111101101101001011010000101" when "0100111101",
      "10001110100100111010001010011011111000000100001111" when "0100111110",
      "10100100011010100000001000110011010111000101011010" when "0100111111",
      "00111010010001011101100000010001011111111101010100" when "0101000000",
      "01010000001001110010010110010100000010000001111010" when "0101000001",
      "01100110000011011110110000011001000010100000110110" when "0101000010",
      "01111011111110100010110011111110111100100000110000" when "0101000011",
      "10010001111010111110100110100100100001000010100111" when "0101000100",
      "10100111111000110010001101101000110111000011001110" when "0101000101",
      "10111101110111111101101110101011011011011100011101" when "0101000110",
      "11010011111000100001001111001100000001000110101010" when "0101000111",
      "00101001111010011100110100101010110000111010000111" when "0101001000",
      "00111111111101110000100100101000001001110000010010" when "0101001001",
      "01010110000010011100100100100101000000100101010010" when "0101001010",
      "01101100001000100000111010000010100000011001001100" when "0101001011",
      "10000010001111111101101010100010001010010001100001" when "0101001100",
      "10011000011000110010111011100101110101011010011111" when "0101001101",
      "10101110100011000000110010101111101111001000011111" when "0101001110",
      "11000100101110100111010101100010011010111001011010" when "0101001111",
      "00011010111011100110101001100000110010010110000101" when "0101010000",
      "00110001001001111110110100001110000101010011100110" when "0101010001",
      "01000111011001101111111011001101111001110100110000" when "0101010010",
      "01011101101010111010000100000100001100001011011011" when "0101010011",
      "01110011111101011101010100010101001110111001111100" when "0101010100",
      "10001010010001011001110001100101101010110100011110" when "0101010101",
      "10100000100110101111100001011010011111000010011101" when "0101010110",
      "10110110111101011110101001011001000000111111111101" when "0101010111",
      "00001101010101100111001111000110111100011111000110" when "0101011000",
      "00100011101111001001011000001010010011101001011010" when "0101011001",
      "00111010001010000101001010001001011111000001010010" when "0101011010",
      "01010000100110011010101010101011001101100011010101" when "0101011011",
      "01100111000100001001111111010110100100100111110100" when "0101011100",
      "01111101100011010011001101110011000000000011111111" when "0101011101",
      "10010100000011110110011011101000010010001011100111" when "0101011110",
      "10101010100101110011101110011110100011110010001111" when "0101011111",
      "00000001001001001011001011111110010100001100101101" when "0101100000",
      "00010111101101111100111001110000011001010010100000" when "0101100001",
      "00101110010100001000111101011101111111011111001101" when "0101100010",
      "01000100111011101111011100110000101001110011110110" when "0101100011",
      "01011011100100110000011101010010010001111000011000" when "0101100100",
      "01110010001111001100000100101101000111111101000001" when "0101100101",
      "10001000111011000010011000101011110010111011110010" when "0101100110",
      "10011111101000010011011110111001010000011001110001" when "0101100111",
      "00110110010110111111011101000000110100101000101000" when "0101101000",
      "01001101000111000110011000101110001010101000000010" when "0101101001",
      "01100011111000101000010111101101010100000111000001" when "0101101010",
      "01111010101011100101011111101010101001100101011100" when "0101101011",
      "10010001011111111101110110010010111010010101011011" when "0101101100",
      "10101000010101110001100001010011001100011100110000" when "0101101101",
      "10111111001101000000100110011000111100110110010001" when "0101101110",
      "11010110000101101011001011010001111111010011011000" when "0101101111",
      "00101100111111110001010101101100011110011101011011" when "0101110000",
      "01000011111011010011001011010110111011110111001001" when "0101110001",
      "01011010111000010000110010000000001111111110000010" when "0101110010",
      "01110001110110101010001111010111101010001011111010" when "0101110011",
      "10001000110110011111101001001100110000111000001110" when "0101110100",
      "10011111110111110001000101001111100001011001100010" when "0101110101",
      "10110110111010011110101001010000010000000111000000" when "0101110110",
      "11001101111110101000011010111111101000011001101111" when "0101110111",
      "00100101000100001110100000001110101100101110010011" when "0101111000",
      "00111100001011010000111110101110110110100110000110" when "0101111001",
      "01010011010011101111111100010001110110101000111001" when "0101111010",
      "01101010011101101011011110101001110100100110001101" when "0101111011",
      "10000001101001000011101011101001001111010110101110" when "0101111100",
      "10011000110101111000101001000010111100111101110101" when "0101111101",
      "10110000000100001010011100101010001010101010111111" when "0101111110",
      "11000111010011111001001100010010011100111011001111" when "0101111111",
      "00011110100101000100111101101111101111011010100110" when "0110000000",
      "00110101110111101101110110110110010101000101100011" when "0110000001",
      "01001101001011110011111101011010111000001010100000" when "0110000010",
      "01100100100001010111010111010010011010001011001101" when "0110000011",
      "01111011111000011000001010010010010011111110010000" when "0110000100",
      "10010011010000110110011100010000010101110000100001" when "0110000101",
      "10101010101010110010010011000010100111000110100111" when "0110000110",
      "11000010000110001011110100011111100110111110010111" when "0110000111",
      "00011001100011000011000110011110001011110000001111" when "0110001000",
      "00110001000001011000001110110101100011010000110111" when "0110001001",
      "01001000100001001011010011011101010010110010011101" when "0110001010",
      "01100000000010011100011010001101010111000110010011" when "0110001011",
      "01110111100101001011101000111110000100011110001100" when "0110001100",
      "10001111001001011001000101101000000110101101111100" when "0110001101",
      "10100110101111000100110110000100100001001100110110" when "0110001110",
      "10111110010110001111000000001100101110110111001001" when "0110001111",
      "00010101111110110111101001111010100010001111011110" when "0110010000",
      "00101101101000111110111001001000000101100000011010" when "0110010001",
      "01000101010100100100110011101111111010011101110110" when "0110010010",
      "01011101000001101001011111101100111010100110100110" when "0110010011",
      "01110100110000001101000010111010010111000101110000" when "0110010100",
      "10001100100000001111100011010011111000110100001111" when "0110010101",
      "10100100010001110001000110110101100000011010010010" when "0110010110",
      "10111100000100110001110011011011100110010000111010" when "0110010111",
      "00010011111001010001101111000010111010100011010111" when "0110011000",
      "00101011101111010000111111101000100101010000101011" when "0110011001",
      "01000011100110101111101011001010000110001101001000" when "0110011010",
      "01011011011111101101110111100101010101000011101110" when "0110011011",
      "01110011011010001011101010111000100001010111101100" when "0110011100",
      "10001011010110001001001011000010010010100101111111" when "0110011101",
      "10100011010011100110011110000001101000000110110000" when "0110011110",
      "10111011010010100011101001110101111001001110111000" when "0110011111",
      "00010011010011000000110100011110110101010001011101" when "0110100000",
      "00101011010100111110000011111100100011100001001111" when "0110100001",
      "01000011011000011011011110001111100011010010001111" when "0110100010",
      "01011011011101011001001001011000101011111011001010" when "0110100011",
      "01110011100011110111001011011001001100110110111001" when "0110100100",
      "10001011101011110101101010010010101101100110000100" when "0110100101",
      "10100011110101010100101100000111001101110000100011" when "0110100110",
      "10111100000000010100010110111001000101000110111011" when "0110100111",
      "00010100001100110100110000101011000011100011111111" when "0110101000",
      "00101100011010110101111111100000010001001110010101" when "0110101001",
      "01000100101010011000001001011100001110011001110010" when "0110101010",
      "01011100111011011011010100100010110011101000111101" when "0110101011",
      "01110101001101111111100110111000010001101110101111" when "0110101100",
      "10001101100010000101000110100001010001101111110111" when "0110101101",
      "10100101110111101011111001100010110101000100010110" when "0110101110",
      "10111110001110110100000110000010010101011001000101" when "0110101111",
      "00010110100111011101110010000101100100110001010100" when "0110110000",
      "00101111000001101001000011110010101101101000001100" when "0110110001",
      "01000111011101010110000001010000010010110010010000" when "0110110010",
      "01011111111010100100110000100101001111011111000001" when "0110110011",
      "01111000011001010101010111111000110111011010011010" when "0110110100",
      "10010000111001100111111101010010110110101110011010" when "0110110101",
      "10101001011011011100100110111011010010000100011111" when "0110110110",
      "11000001111110110011011010111010100110100111001011" when "0110110111",
      "00011010100011101100011111011001101010000011100111" when "0110111000",
      "00110011001010000111111010100001101010101011000001" when "0110111001",
      "01001011110010000101110010011100001111010100010110" when "0110111010",
      "01100100011011100110001101010011010111011101101010" when "0110111011",
      "01111101000110101001010001010001011011001101110101" when "0110111100",
      "10010101110011001111000100100001001011010101111110" when "0110111101",
      "10101110100001010111101101001101110001010011000001" when "0110111110",
      "11000111010001000011010001100010101111001111010010" when "0110111111",
      "00100000000010010001110111101100000000000011111110" when "0111000000",
      "00111000110101000011100101110101110111011010101111" when "0111000001",
      "01010001101001011000100010001101000001101111010001" when "0111000010",
      "01101010011111010000110010111110100100010000110010" when "0111000011",
      "10000011010110101100011110010111111101000011100101" when "0111000100",
      "10011100001111101011101010100111000011000010101011" when "0111000101",
      "10110101001010001110011101111010000110000001001110" when "0111000110",
      "11001110000110010100111110011111101110101100001100" when "0111000111",
      "00100111000011111111010010100110111110101011110111" when "0111001000",
      "01000000000011001101100000011111010000100101011000" when "0111001001",
      "01011001000011111111101110011000010111111100010111" when "0111001010",
      "01110010000110010110000010100010100001010100011001" when "0111001011",
      "10001011001010010000100011001110010010010010101010" when "0111001100",
      "10100100001111101111010110101100101001011111011110" when "0111001101",
      "10111101010110110010100011001110111110100111110010" when "0111001110",
      "11010110011111011010001111000111000010011110111010" when "0111001111",
      "00101111101001100110100000100110111110111111111011" when "0111010000",
      "01001000110101010111011110000001010111001111010110" when "0111010001",
      "01100010000010101101001101101001000111011100101010" when "0111010010",
      "01111011010001100111110101110001100101000011111000" when "0111010011",
      "10010100100010000111011100101110011110101111001100" when "0111010100",
      "10101101110100001100001000110011111100011000011101" when "0111010101",
      "11000111000111110110000000010110011111001010110100" when "0111010110",
      "11100000011101000101001001101011000001100100010100" when "0111010111",
      "00111001110011111001101011000110110111010111011010" when "0111011000",
      "01010011001100010011101010111111101101101100100100" when "0111011001",
      "01101100100110010011001111101011101011000011111010" when "0111011010",
      "10000110000001111000011111100001001111010110101111" when "0111011011",
      "10011111011111000011100000110111010011111001001010" when "0111011100",
      "10111000111101110100011010000101001011011011100111" when "0111011101",
      "11010010011110001011010001100010100010001100100011" when "0111011110",
      "11101100000000001000001101100111011101111001111110" when "0111011111",
      "00000101100011101011010100101100011101110011000001" when "0111100000",
      "00011111001000110100101101001010011010101001100111" when "0111100001",
      "00111000101111100100011101011010100110110011111111" when "0111100010",
      "01010010010111111010101011110110101110001110010110" when "0111100011",
      "01101100000001110111011110111000110110011100011011" when "0111100100",
      "10000101101101011010111100111011011110101011001000" when "0111100101",
      "10011111011010100101001100011001011111110010000110" when "0111100110",
      "10111001001001010110010011101110001100010101010101" when "0111100111",
      "00010010111001101110011001010101010000100110110010" when "0111101000",
      "00101100101011101101100011101010110010101000000000" when "0111101001",
      "01000110011111010011111001001011010010001011101101" when "0111101010",
      "01100000010100100001100000010011101000110111011010" when "0111101011",
      "01111010001011010110011111100001001010000101000001" when "0111101100",
      "10010100000011110010111101010001100011000100011110" when "0111101101",
      "10101101111101110111000000000010111010111101010111" when "0111101110",
      "11000111111001100010101110010011110010110000100000" when "0111101111",
      "00100001110110110110001110100011000101011001100101" when "0111110000",
      "00111011110101110001100111010000000111110000110100" when "0111110001",
      "01010101110110010100111110111010101000101100100000" when "0111110010",
      "01101111111000100000011100000010110001000010101101" when "0111110011",
      "10001001111100010100000101001001000011101010110101" when "0111110100",
      "10100100000001110000000000101110011101011111010011" when "0111110101",
      "10111110001000110100010101010100010101011111001000" when "0111110110",
      "11011000010001100001001001011100011100101111100111" when "0111110111",
      "00110010011011110110100011101000111110011101111011" when "0111111000",
      "01001100100111110100101010011100100000000000101111" when "0111111001",
      "01100110110101011011100100011010000000111001111001" when "0111111010",
      "10000001000100101011011000000100111010111000000001" when "0111111011",
      "10011011010101100100001100000001000001111000001011" when "0111111100",
      "10110101101000000110000110110010100100000111011110" when "0111111101",
      "11001111111100010001001110111110001010000100101111" when "0111111110",
      "11101010010010000101101011001000110110100010001011" when "0111111111",
      "00010001011001011111100011011111001011000001010000" when "1000000000",
      "00011011000110111000100100000010011101100011001011" when "1000000001",
      "00100100110100111000011011010111011111000001111011" when "1000000010",
      "00101110100011011111001011111001101111011011010111" when "1000000011",
      "00111000010010101100111000000100111000011011101100" when "1000000100",
      "01000010000010100001100010010100101101011101111111" when "1000000101",
      "01001011110010111101001101000101001011101100111001" when "1000000110",
      "01010101100011111111111010110010011010000011000111" when "1000000111",
      "00011111010101101001101101111000101001001100001010" when "1000001000",
      "00101001000111111010101000110100010011100100110101" when "1000001001",
      "00110010111010110010101110000001111101011011111010" when "1000001010",
      "00111100101110010001111111111110010100110010110010" when "1000001011",
      "01000110100010011000100001000110010001011101111101" when "1000001100",
      "01010000010111000110010011110110110101000101110001" when "1000001101",
      "01011010001100011011011010101101001011000110111110" when "1000001110",
      "01100100000010010111111000000110101000110011010100" when "1000001111",
      "00101101111000111011101110100000101101010010001101" when "1000010000",
      "00110111110000000111000000011001000001100001010010" when "1000010001",
      "01000001100111111001110000001101011000010101000110" when "1000010010",
      "01001011100000010100000000011011101110011001101001" when "1000010011",
      "01010101011001010101110011100010001010010011000001" when "1000010100",
      "01011111010010111111001011111110111100011110000011" when "1000010101",
      "01101001001101010000001100010000011111010000111010" when "1000010110",
      "01110011001000001000110110110101010110111011101110" when "1000010111",
      "00111101000011101001001110001100010001101001001011" when "1000011000",
      "01000110111111110001010100110100000111011111001010" when "1000011001",
      "01010000111100100001001101001011111010011111011000" when "1000011010",
      "01011010111001111000111001110010110110100111111111" when "1000011011",
      "01100100110111111000011101001000010001110100001011" when "1000011100",
      "01101110110110011111111001101011101011111100110110" when "1000011101",
      "01111000110101101111010001111100101110111001001011" when "1000011110",
      "10000010110101100110101000011011001110011111010011" when "1000011111",
      "00001100110110000101111111100111001000100100110111" when "1000100000",
      "00010110110111001101011010000000100100111111101111" when "1000100001",
      "00100000111000111100111010000111110101100110100101" when "1000100010",
      "00101010111011010100100010011101010110010001011100" when "1000100011",
      "00110100111110010100010101100001101100111010011110" when "1000100100",
      "00111111000001111100010101110101101001011110100000" when "1000100101",
      "01001001000110001100100101111010000101111101101010" when "1000100110",
      "01010011001011000101001000010000000110011011111111" when "1000100111",
      "00011101010000100101111111011000111001000010001010" when "1000101000",
      "00100111010110101111001101110101110101111110000000" when "1000101001",
      "00110001011101100000110110001000011111100011001010" when "1000101010",
      "00111011100100111010111010110010100010001011110010" when "1000101011",
      "01000101101100111101011110010101110100011001000101" when "1000101100",
      "01001111110101101000100011010100010110110100000000" when "1000101101",
      "01011001111110111100001100010000010100001101110101" when "1000101110",
      "01100100001000111000011011101100000001100000110110" when "1000101111",
      "00101110010011011101010100001001111101110000111111" when "1000110000",
      "00111000011110101010111000001100110010001100011010" when "1000110001",
      "01000010101010100001001010010111010010001100001010" when "1000110010",
      "01001100110111000000001101001100011011010100110111" when "1000110011",
      "01010111000100001000000011001111010101010111010000" when "1000110100",
      "01100001010001111000101111000011010010010000111010" when "1000110101",
      "01101011100000010010010011001011101110001100110110" when "1000110110",
      "01110101101111010100110010001100001111100100001000" when "1000110111",
      "00111111111111000000001110101000100110111110100101" when "1000111000",
      "01001010001111010100101011000100101111010011010110" when "1000111001",
      "01010100100000010010001010000100101101101001100111" when "1000111010",
      "01011110110001111000101110001100110001011001001010" when "1000111011",
      "01101001000100001000011010000001010100001011000101" when "1000111100",
      "01110011010111000001010000000110111001111010011010" when "1000111101",
      "01111101101010100011010011000010010000110100101011" when "1000111110",
      "10000111111110101110100101011000010001011010101101" when "1000111111",
      "00010010010011100011001001101101111110100001000111" when "1001000000",
      "00011100101001000001000010101000100101010001000010" when "1001000001",
      "00100110111111001000010010101101011101001000110010" when "1001000010",
      "00110001010101111000111100100010000111111100011010" when "1001000011",
      "00111011101101010011000010101100010001110110011010" when "1001000100",
      "01000110000101010110100111110001110001011000011010" when "1001000101",
      "01010000011110000011101110011000100111011011101110" when "1001000110",
      "01011010110111011010011001000110111111010010000010" when "1001000111",
      "00100101010001011010101010100011001110100110000111" when "1001001000",
      "00101111101100000100100101010011110101011100010110" when "1001001001",
      "00111010000111011000001011111111011110010011011111" when "1001001010",
      "01000100100011010101100001001100111110000101010001" when "1001001011",
      "01001110111111111100100111100011010100000111000010" when "1001001100",
      "01011001011101001101100001101001101010001010011100" when "1001001101",
      "01100011111011001000010010000111010100011110000100" when "1001001110",
      "01101110011001101100111011100011110001101110000011" when "1001001111",
      "00111000111000111011100000100110101011000100110110" when "1001010000",
      "01000011011000110100000011110111110100001011110001" when "1001010001",
      "01001101111001010110100111111111001011001011101010" when "1001010010",
      "01011000011010100011001111100100111000101101101000" when "1001010011",
      "01100010111100011001111101010001001111111011100111" when "1001010100",
      "01101101011110111010110011101100101110100001000110" when "1001010101",
      "01111000000010000101110101011111111100101011101111" when "1001010110",
      "10000010100101111011000101010011101101001100000011" when "1001010111",
      "00001101001010011010100101110000111101010110000010" when "1001011000",
      "00010111101111100100011001100000110101000001111000" when "1001011001",
      "00100010010101011000100011001100100110101100100010" when "1001011010",
      "00101100111011110111000101011101101111011000100001" when "1001011011",
      "00110111100011000000000010111101110110101110011011" when "1001011100",
      "01000010001010110011011110010110101110111101101100" when "1001011101",
      "01001100110011010001011010010010010100111101001111" when "1001011110",
      "01010111011100011001111001011010110000001100000101" when "1001011111",
      "00100010000110001100111110011010010010110010000101" when "1001100000",
      "00101100110000101010101011111011011001100000100001" when "1001100001",
      "00110111011011110011000100101000101011110010110101" when "1001100010",
      "01000010000111100110001011001100111011101111010001" when "1001100011",
      "01001100110100000100000010010011000110000111100000" when "1001100100",
      "01010111100001001100101100100110010010011001011001" when "1001100101",
      "01100010001111000000001100110001110010101111100011" when "1001100110",
      "01101100111101011110100101100001000100000010000101" when "1001100111",
      "00110111101100100111111001011111101101110111001110" when "1001101000",
      "01000010011100011100001011011001100010100100000010" when "1001101001",
      "01001101001100111011011101111010011111001101000010" when "1001101010",
      "01010111111110000101110011101110101011100110111011" when "1001101011",
      "01100010101111111011001111100010011010010111001100" when "1001101100",
      "01101101100010011011110100000010001000110100111000" when "1001101101",
      "01111000010101100111100011111010011111001001001000" when "1001101110",
      "10000011001001011110100001111000010000001111111111" when "1001101111",
      "00001101111110000000110000101000011001111000111111" when "1001110000",
      "00011000110011001110010010111000000100100111111001" when "1001110001",
      "00100011101001000111001011010100100011110101010100" when "1001110010",
      "00101110011111101011011100101011010101101111011011" when "1001110011",
      "00111001010110111011001001101010000011011010100111" when "1001110100",
      "01000100001110110110010100111110100000110010001011" when "1001110101",
      "01001111000111011101000001010110101100101001000000" when "1001110110",
      "01011010000000101111010001100000110000101010010000" when "1001110111",
      "00100100111010101101001000001011000001011010000000" when "1001111000",
      "00101111110101010110101000000011111110010110000000" when "1001111001",
      "00111010110000101011110011111010010001110110010001" when "1001111010",
      "01000101101100101100101110011100110001001101110100" when "1001111011",
      "01010000101001011001011010011010011100101011010101" when "1001111100",
      "01011011100110110001111010100010011111011001111000" when "1001111101",
      "01100110100100110110010001100100001111100001100001" when "1001111110",
      "01110001100011100110100010001111001110001000000111" when "1001111111",
      "00111100100011000010101111010011000111010001110101" when "1010000000",
      "01000111100011001010111011011111110010000010000010" when "1010000001",
      "01010010100011111111001001100101010000011011110101" when "1010000010",
      "01011101100101011111011100010011101111100010110001" when "1010000011",
      "01101000100111101011110110011011100111011011100111" when "1010000100",
      "01110011101010100100011010101101011011001100111100" when "1010000101",
      "01111110101110001001001011111001111000111111111000" when "1010000110",
      "10001001110010011010001100110001111010000000110010" when "1010000111",
      "00010100110111010111100000000110100010011111111100" when "1010001000",
      "00011111111101000001001000101001000001110010001111" when "1010001001",
      "00101011000011010111001001001010110010010001110110" when "1010001010",
      "00110110001010011001100100011101011001011110111111" when "1010001011",
      "01000001010010001000011101010010101000000000100001" when "1010001100",
      "01001100011010100011110110011100011001100100101101" when "1010001101",
      "01010111100011101011110010101100110101000001111010" when "1010001110",
      "01100010101101100000010100110110001100010111001111" when "1010001111",
      "00101101111000000001011111101010111100101101010011" when "1010010000",
      "00111001000011001111010101111101101110010110110110" when "1010010001",
      "01000100001111001001111010100001010100110001100001" when "1010010010",
      "01001111011011110001010000001000101110100110100001" when "1010010011",
      "01011010101001000101011001100111000101101011010010" when "1010010100",
      "01100101110111000110011001101111101111000010010000" when "1010010101",
      "01110001000101110100010011010110001010111011100010" when "1010010110",
      "01111100010101001111001001001110000100110101100101" when "1010010111",
      "00000111100101010110111110001011010011011101111010" when "1010011000",
      "00010010110110001011110101000001111000110001110100" when "1010011001",
      "00011110000111101101110000100110000001111111000100" when "1010011010",
      "00101001011001111100110011101100000111100100101001" when "1010011011",
      "00110100101100111001000001001000101101010011010110" when "1010011100",
      "01000000000000100010011011110000100010001110100111" when "1010011101",
      "01001011010100111001000110011000100000101101001001" when "1010011110",
      "01010110101001111101000011110101101110011001101011" when "1010011111",
      "00100001111111101110010110111101011100010011100111" when "1010100000",
      "00101101010110001101000010100101000110101111110011" when "1010100001",
      "00111000101101011001001001100010010101011001001101" when "1010100010",
      "01000100000101010010101110101010111011010001100111" when "1010100011",
      "01001111011101111001110100110100110110110010011001" when "1010100100",
      "01011010110111001110011110110110010001101101000111" when "1010100101",
      "01100110010001010000101111100101100001001100010111" when "1010100110",
      "01110001101100000000101001111001000101110100010111" when "1010100111",
      "00111101000111011110010000100111101011100011110001" when "1010101000",
      "01001000100011101001100110101000001001110100010100" when "1010101001",
      "01010100000000100010101110110001100011011011100011" when "1010101010",
      "01011111011110001001101011111011000110101011100110" when "1010101011",
      "01101010111100011110100000111100001101010011110010" when "1010101100",
      "01110110011011100001010000101100011100100001011011" when "1010101101",
      "10000001111011010001111110000011100101000000100010" when "1010101110",
      "10001101011011110000101011111001100010111100100000" when "1010101111",
      "00011000111100111101011101000110011110000000110101" when "1010110000",
      "00100100011110111000010100100010101001011001111010" when "1010110001",
      "00110000000001100001010101000110100011110101101001" when "1010110010",
      "00111011100100111000100001101010110111100100010000" when "1010110011",
      "01000111001000111101111101001000011010011000111010" when "1010110100",
      "01010010101101110001101010011000001101101010100011" when "1010110101",
      "01011110010011010011101100010011011110010100100011" when "1010110110",
      "01101001111001100100000101110011100100110111011101" when "1010110111",
      "00110101100000100010111001110010000101011001101100" when "1010111000",
      "01000001001000010000001011001000101111101000010100" when "1010111001",
      "01001100110000101011111100110001011110110111101111" when "1010111010",
      "01011000011001110110010001100110011010000100011011" when "1010111011",
      "01100100000011101111001100100001110011110011101000" when "1010111100",
      "01101111101110010110110000011110001010010100001010" when "1010111101",
      "01111011011001101101000000010110000111011111000011" when "1010111110",
      "10000111000101110001111111000100100000111000010101" when "1010111111",
      "00010010110010100101101111100100010111101111110001" when "1011000000",
      "00011110100000001000010100110000111001000001100001" when "1011000001",
      "00101010001110011001110001100101011101010110111100" when "1011000010",
      "00110101111101011010001000111101101001000111010101" when "1011000011",
      "01000001101101001001011101110101001100011000100100" when "1011000100",
      "01001101011101100111110011001000000010111111111100" when "1011000101",
      "01011001001110110101001011110010010100100010110101" when "1011000110",
      "01100101000000110001101010110000010100010111011101" when "1011000111",
      "00110000110011011101010010111110100001100101101001" when "1011001000",
      "00111100100110111000000111011001100111000111011111" when "1011001001",
      "01001000011011000010001010111110011011101010001011" when "1011001010",
      "01010100001111111011100000101010000001101110101001" when "1011001011",
      "01100000000101100100001011011001100111101010011000" when "1011001100",
      "01101011111011111100001110001010100111101000001000" when "1011001101",
      "01110111110011000011101011111010100111101000101010" when "1011001110",
      "10000011101010111010100111100111011001100011011101" when "1011001111",
      "00001111100011100001000100001110111011000111100000" when "1011010000",
      "00011011011100110111000100101111010101111100000001" when "1011010001",
      "00100111010110111100101100000110111111100001001101" when "1011010010",
      "00110011010001110001111101010100011001010000111101" when "1011010011",
      "00111111001101010110111011010110010000011111101001" when "1011010100",
      "01001011001001101011101001001011011110011100110100" when "1011010101",
      "01010111000110110000001001110011001000010100000001" when "1011010110",
      "01100011000100100100100000001100011111001101011101" when "1011010111",
      "00101111000011001000101111010111000000001110110010" when "1011011000",
      "00111011000010011100111010010010010100011011111000" when "1011011001",
      "01000111000010100001000011111110010000110111100000" when "1011011010",
      "01010011000011010101001111011010110110100100001011" when "1011011011",
      "01011111000100111001011111101000010010100100110010" when "1011011100",
      "01101011000111001101110111100110111101111101011110" when "1011011101",
      "01110111001010010010011010010111011101110100010010" when "1011011110",
      "10000011001110000111001010111010100011010001111110" when "1011011111",
      "00001111010010101100001100010001001011100010101111" when "1011100000",
      "00011011011000000001100001011100011111110110111111" when "1011100001",
      "00100111011110000111001101011101110101100100000101" when "1011100010",
      "00110011100100111101010011010110101110000101000100" when "1011100011",
      "00111111101100100011110110001000110110111011100000" when "1011100100",
      "01001011110100111010111000110110001001110000001001" when "1011100101",
      "01010111111110000010011110100000101100010011101101" when "1011100110",
      "01100100000111111010101010001010110000011111101101" when "1011100111",
      "00110000010010100011011110110110110100010111000101" when "1011101000",
      "00111100011101111100111111100111100010000111000111" when "1011101001",
      "01001000101010000111001111011111110000001000000001" when "1011101010",
      "01010100110111000010010001100010100000111101110110" when "1011101011",
      "01100001000100101110001000110011000011011001001010" when "1011101100",
      "01101101010011001010111000010100110010010111110110" when "1011101101",
      "01111001100010011000100011001011010101000101110111" when "1011101110",
      "10000101110010010111001100011010011110111101111101" when "1011101111",
      "00010010000011000110110111000110001111101010100010" when "1011110000",
      "00011110010100100111100110010010110011000110010011" when "1011110001",
      "00101010100110111001011101000100100001011101001001" when "1011110010",
      "00110110111001111100011110011111111111001100110011" when "1011110011",
      "01000011001101110000101101101001111101000101101101" when "1011110100",
      "01001111100010010110001101100111011000001011101101" when "1011110101",
      "01011011110111101101000001011101011001110110110110" when "1011110110",
      "01101000001101110101001100010001010111110100001011" when "1011110111",
      "00110100100100101110110001001000110100000110011101" when "1011111000",
      "01000000111100011001110011001001011101000110111100" when "1011111001",
      "01001101010100110110010101011001001101100110001111" when "1011111010",
      "01011001101110000100011010111110001100101100111100" when "1011111011",
      "01100110001000000100000110111110101101111100100010" when "1011111100",
      "01110010100010110101011100100001010001010000000011" when "1011111101",
      "01111110111110011000011110101100100010111100111110" when "1011111110",
      "10001011011010101101010000100111011011110011111001" when "1011111111",
      "00010111110111110011110101011001000001000001010111" when "1100000000",
      "00100100010101101100010000001000100100001110101001" when "1100000001",
      "00110000110100010110100011111101100011100010011110" when "1100000010",
      "00111101010011110010110011111111101001100001111000" when "1100000011",
      "01001001110100000001000011010110101101010000111100" when "1100000100",
      "01010110010101000001010101001010110010010011100011" when "1100000101",
      "01100010110110110011101100100100001000101110010000" when "1100000110",
      "01101111011001011000001100101011001101000110111011" when "1100000111",
      "00111011111100101110111000101000101000100101101100" when "1100001000",
      "01001000100000110111110011100101010000110101100110" when "1100001001",
      "01010101000101110011000000101010001000000101011100" when "1100001010",
      "01100001101011100000100011000000011101001000100011" when "1100001011",
      "01101110010010000000011101110001101011010111100110" when "1100001100",
      "01111010111001010010110100000111011010110001010100" when "1100001101",
      "10000111100001010111101001001011011111111011011000" when "1100001110",
      "10010100001010001111000000000111111100000011000111" when "1100001111",
      "00100000110011111000111100000110111100111110010100" when "1100010000",
      "00101101011110010101100000010010111101001100000011" when "1100010001",
      "00111010001001100100101111110110100011110101011011" when "1100010010",
      "01000110110101100110101101111100100100101110011001" when "1100010011",
      "01010011100010011011011101110000000000010110100100" when "1100010100",
      "01100000010000000011000010011100000011111001111011" when "1100010101",
      "01101100111110011101011111001100001001010001101111" when "1100010110",
      "01111001101101101010110111001011110111000101010000" when "1100010111",
      "00000110011101101011001101100111000000101010100010" when "1100011000",
      "00010011001110011110100101101001100110000111001111" when "1100011001",
      "00100000000000000101000010011111110100010001011110" when "1100011010",
      "00101100110010011110100111010110000100110000011111" when "1100011011",
      "00111001100101101011010111011000111101111101100100" when "1100011100",
      "01000110011001101011010101110101010011000100110011" when "1100011101",
      "01010011001110011110100101111000000100000101110111" when "1100011110",
      "01100000000100000101001010101110011101110100110100" when "1100011111",
      "00101100111010011111000111100101111001111010111101" when "1100100000",
      "00111001110001101100011111101011111110110111100100" when "1100100001",
      "01000110101001101101010110001110100000000000101111" when "1100100010",
      "01010011100010100001101110011011011101100100001010" when "1100100011",
      "01100000011100001001101011100001000100100111111101" when "1100100100",
      "01101101010110100101010000101101101111001011011101" when "1100100101",
      "01111010010001110100100001010000000100001000000011" when "1100100110",
      "10000111001101110111100000010110110111010001111011" when "1100100111",
      "00010100001010101110010001010001001001011000111100" when "1100101000",
      "00100001001000011000110111001110001000001001010111" when "1100101001",
      "00101110000110110111010101011101001110001100110001" when "1100101010",
      "00111011000110001001101111001110000011001010110001" when "1100101011",
      "01001000000110010000000111110000011011101001111001" when "1100101100",
      "01010101000111001010100010010100011001010000010101" when "1100101101",
      "01100010001000111001000010001010001010100100110010" when "1100101110",
      "01101111001011011011101010100010001011001111010010" when "1100101111",
      "00111100001110110010011110101101000011111010000000" when "1100110000",
      "01001001010010111101100001111011101010010010000011" when "1100110001",
      "01010110010111111100110111011111000001001000010011" when "1100110010",
      "01100011011101110000100010101000011000010010001100" when "1100110011",
      "01110000100100011000100110101001001100101010100110" when "1100110100",
      "01111101101011110101000110110011001000010010100101" when "1100110101",
      "10001010110100000110000110011000000010010010010000" when "1100110110",
      "10010111111101001011101000101001111110111001100101" when "1100110111",
      "00100101000111000101110000111011001111100001001100" when "1100111000",
      "00110010010001110100100010011110010010101011001111" when "1100111001",
      "00111111011101011000000000100101110100000100001001" when "1100111010",
      "01001100101001110000001110100100101100100011100011" when "1100111011",
      "01011001110110111101001111101110000010001100111111" when "1100111100",
      "01100111000100111111000111010101001000010000110100" when "1100111101",
      "01110100010011110101111000101101011111001101000010" when "1100111110",
      "10000001100011100001100111001010110100101110000001" when "1100111111",
      "00001110110100000010010110000001000011101111011110" when "1101000000",
      "00011100000101011000001000100100010100011101001011" when "1101000001",
      "00101001010111100011000010001000111100010011110101" when "1101000010",
      "00110110101010100011000110000011011110000001111010" when "1101000011",
      "01000011111110011000010111101000101001101000011101" when "1101000100",
      "01010001010011000010111010001101011100011011111011" when "1101000101",
      "01011110101000100010110001000111000001000101000010" when "1101000110",
      "01101011111110110111111111101010101111100001100101" when "1101000111",
      "00111001010110000010101001001110001101000101010010" when "1101001000",
      "01000110101110000010110001000111001100011010100101" when "1101001001",
      "01010100000110111000011010101011101101100011100010" when "1101001010",
      "01100001100000100011101001010001111101111010100101" when "1101001011",
      "01101110111011000100100000010000011000010011011110" when "1101001100",
      "01111100010110011011000010111101100100111011111111" when "1101001101",
      "10001001110010100111010100110000011001011100111010" when "1101001110",
      "10010111001111101001011000111111111000111010101110" when "1101001111",
      "00100100101101100001010011000011010011110110100101" when "1101010000",
      "00110010001100001111000110010010001000001111000100" when "1101010001",
      "00111111101011110010110110000100000001100001000010" when "1101010010",
      "01001101001100001100100101110000111000101000100010" when "1101010011",
      "01011010101101011100011000110000110100000001100010" when "1101010100",
      "01101000001111100010010010011100000111101000110111" when "1101010101",
      "01110101110010011110010110001011010100111101000001" when "1101010110",
      "10000011010110010000100111010111001010111110111111" when "1101010111",
      "00010000111010111001001001011000100110010011001010" when "1101011000",
      "00011110100000010111111111101000110001000010000101" when "1101011001",
      "00101100000110101101001101100001000010111001011011" when "1101011010",
      "00111001101101111000110110011011000001001100101100" when "1101011011",
      "01000111010101111010111101110000011110110110001110" when "1101011100",
      "01010100111110110011100110111011011100010111111000" when "1101011101",
      "01100010101000100010110101010110000111111100000011" when "1101011110",
      "01110000010011001000101100011010111101010110011001" when "1101011111",
      "00111101111110100101001111100100100110000100110001" when "1101100000",
      "01001011101010111000100010001101111001010000000010" when "1101100001",
      "01011001011000000010100111110001111011101100111010" when "1101100010",
      "01100111000110000011100011101011111111111100110111" when "1101100011",
      "01110100110100111011011001010111100110001110111011" when "1101100100",
      "10000010100100101010001100010000011100100000101000" when "1101100101",
      "10010000010101001111111111110010011110011110101110" when "1101100110",
      "10011110000110101100110111011001110101100110001101" when "1101100111",
      "00101011111001000000110110100010111001000101000000" when "1101101000",
      "00111001101100001100000000101010001101111011000001" when "1101101001",
      "01000111100000001110011001001100100110111010110101" when "1101101010",
      "01010101010101001000000011100111000100101010101001" when "1101101011",
      "01100011001010111001000011010110110101100101001000" when "1101101100",
      "01110001000001100001011011111001010101111010010100" when "1101101101",
      "01111110111001000001010000101100001111110000011001" when "1101101110",
      "10001100110001011000100101001101011011000100101001" when "1101101111",
      "00011010101010100111011100111010111101101100010000" when "1101110000",
      "00101000100100101101111011010011001011010101001111" when "1101110001",
      "00110110011111101100000011110100100101100111010000" when "1101110010",
      "01000100011011100001111001111101111100000100100001" when "1101110011",
      "01010010011000001111100001001110001100001010101000" when "1101110100",
      "01100000010101110100111101000100100001010011011110" when "1101110101",
      "01101110010100010010010001000000010100110110000101" when "1101110110",
      "01111100010011100111100000100001001110000111100001" when "1101110111",
      "00001010010011110100101111000111000010011011101110" when "1101111000",
      "00011000010100111010000000010001110101000110011100" when "1101111001",
      "00100110010110110111010111100001110111011100000001" when "1101111010",
      "00110100011001101100111000010111101000110010010110" when "1101111011",
      "01000010011101011010100110010011110110100001101100" when "1101111100",
      "01010000100010000000100100110111011100000101101001" when "1101111101",
      "01011110100111011110110111100011100010111101111001" when "1101111110",
      "01101100101101110101100001111001100010101111001100" when "1101111111",
      "00111010110101000100100111011011000001000100001100" when "1110000000",
      "01001000111101001100001011101001110001101110010111" when "1110000001",
      "01010111000110001100010010000111110110100110110100" when "1110000010",
      "01100101010000000100111110010111011111101111010001" when "1110000011",
      "01110011011010110110010011111011001011010010110101" when "1110000100",
      "10000001100110100000010110010101100101100110111110" when "1110000101",
      "10001111110011000011001001001001101001001100011000" when "1110000110",
      "10011110000000011110101111111010011110101111110100" when "1110000111",
      "00101100001110110011001110001011011101001011000100" when "1110001000",
      "00111010011110000000100111100000001001100101110000" when "1110001001",
      "01001000101110000110111111011100010111010110010010" when "1110001010",
      "01010110111111000110011001100100001000000010101110" when "1110001011",
      "01100101010000111110111001011011101011100001101011" when "1110001100",
      "01110011100011110000100010100111011111111011001011" when "1110001101",
      "10000001110111011011011000101100010001101001100110" when "1110001110",
      "10010000001011111111011111001110111011011010100010" when "1110001111",
      "00011110100001011100111001110100100110001111101101" when "1110010000",
      "00101100110111110011101100000010101001011111110100" when "1110010001",
      "00111011001111000011111001011110101010110111100000" when "1110010010",
      "01001001100111001101100101101110011110011010001101" when "1110010011",
      "01011000000000010000110100011000000110100011000100" when "1110010100",
      "01100110011010001101101001000001110100000101110011" when "1110010101",
      "01110100110101000100000111010010000110001111101010" when "1110010110",
      "10000011010000110100010010101111101010101000010010" when "1110010111",
      "00010001101101011110001111000001011101010010100111" when "1110011000",
      "00100000001011000001111111101110101000101101110010" when "1110011001",
      "00101110101001011111101000011110100101110110000011" when "1110011010",
      "00111101001000110111001100111000111100000101101100" when "1110011011",
      "01001011101001001000110000100101100001010101110111" when "1110011100",
      "01011010001010010100010111001100011001111111100101" when "1110011101",
      "01101000101100011010000100010101111000111100100100" when "1110011110",
      "01110111001111011001111011101010011111101000001100" when "1110011111",
      "00000101110011010100000000110010111110000000010110" when "1110100000",
      "00010100011000001000010111011000010010100110011001" when "1110100001",
      "00100010111101110111000011000011101010100000000011" when "1110100010",
      "00110001100100100000000111011110100001011000010101" when "1110100011",
      "01000000001100000011101000010010100001100000011010" when "1110100100",
      "01001110110100100001101001001001100011110000100100" when "1110100101",
      "01011101011101111010001101101101101111101001000100" when "1110100110",
      "01101100001000001101011001101001011011010011001011" when "1110100111",
      "00111010110011011011010000100111001011100001111010" when "1110101000",
      "01001001011111100011110110010001110011110011000110" when "1110101001",
      "01011000001100100111001110010100010110010000010000" when "1110101010",
      "01100110111010100101011100011010000011101111011100" when "1110101011",
      "01110101101001011110100100001110011011110100010000" when "1110101100",
      "10000100011001010010101001011101001100110000110000" when "1110101101",
      "10010011001010000001101111110010010011100110010011" when "1110101110",
      "10100001111011101011111010111001111100000110100100" when "1110101111",
      "00110000101110010001001110100000100000110100011001" when "1110110000",
      "00111111100001110001101110010010101011000100110001" when "1110110001",
      "01001110010110001101011101111101010010111111101110" when "1110110010",
      "01011101001011100100100001001101011111100001001110" when "1110110011",
      "01101100000001110110111011110000100110011010001100" when "1110110100",
      "01111010111001000100110001010100001100010001010101" when "1110110101",
      "10001001110001001110000101100110000100100100000110" when "1110110110",
      "10011000101010010010111100010100010001100111101010" when "1110110111",
      "00100111100100010011011001001101000100101001110000" when "1110111000",
      "00110110011111001111011111111110111101110001101100" when "1110111001",
      "01000101011011000111010100011000101100000001001111" when "1110111010",
      "01010100010111111010111010001001001101010101100101" when "1110111011",
      "01100011010101101010010100111111101110101000001110" when "1110111100",
      "01110010010100010101101000101011101011101111111110" when "1110111101",
      "10000001010011111100111000111100101111100001110100" when "1110111110",
      "10010000010100100000001001100010110011110001111010" when "1110111111",
      "00011111010101111111011110001110000001010100011110" when "1111000000",
      "00101110011000011010111010101110101111111110110000" when "1111000001",
      "00111101011011110010100010110101100110100111111110" when "1111000010",
      "01001100100000000110011010010011011011001010001101" when "1111000011",
      "01011011100101010110100100111001010010100011011010" when "1111000100",
      "01101010101011100011000110011000100000110110010100" when "1111000101",
      "01111001110010101100000010100010101001001011011000" when "1111000110",
      "10001000111010110001011101001001011101110001101101" when "1111000111",
      "00011000000011110011011001111111000000000000000011" when "1111001000",
      "00100111001101110001111100110101100000010101101010" when "1111001001",
      "00110110011000101101001001011111011110011011010111" when "1111001010",
      "01000101100100100101000011101111101001000100011000" when "1111001011",
      "01010100110001011001101111011000111110001111011000" when "1111001100",
      "01100011111111001011010000001110101011000111010100" when "1111001101",
      "01110011001101111001101010000100001100000100100000" when "1111001110",
      "10000010011101100101000000101101001100101101011110" when "1111001111",
      "00010001101110001101010111111101100111110111111110" when "1111010000",
      "00100000111111110010110011101001100111101001111000" when "1111010001",
      "00110000010010010101010111100101100101011010001101" when "1111010010",
      "00111111100101110101000111100110001001110010000001" when "1111010011",
      "01001110111010010010000111100000001100101101011000" when "1111010100",
      "01011110001111101100011011001000110101011100011000" when "1111010101",
      "01101101100110000100000110010101011010100011111110" when "1111010110",
      "01111100111101011001001100111011100001111111000100" when "1111010111",
      "00001100010101101011110010110001000000111111011000" when "1111011000",
      "00011011101110111011111011101011111100001110011100" when "1111011001",
      "00101011001001001001101011100010100111101110100100" when "1111011010",
      "00111010100100010101000110001011100110111011110011" when "1111011011",
      "01001010000000011110001111011101101100101100111001" when "1111011100",
      "01011001011101100101001011001111111011010100001110" when "1111011101",
      "01101000111011101001111101011001100100100000110110" when "1111011110",
      "01111000011010101100101001110010001001011111010111" when "1111011111",
      "00000111111010101101010100010001011010111010111101" when "1111100000",
      "00010111011011101100000000101111011000111110010100" when "1111100001",
      "00100110111101101000110011000100010011010100101001" when "1111100010",
      "00110110100000100011101111001000101001001010101000" when "1111100011",
      "01000110000100011100111000110101001001001111010101" when "1111100100",
      "01010101101001010100010100000010110001110101010010" when "1111100101",
      "01100101001111001010000100101010110000110011010110" when "1111100110",
      "01110100110101111110001110100110100011100101110010" when "1111100111",
      "00000100011101110000110101101111110111001111001001" when "1111101000",
      "00010100000110100001111110000000101000011001010010" when "1111101001",
      "00100011110000010001101011010011000011010110011000" when "1111101010",
      "00110011011011000000000001100001100100000001110100" when "1111101011",
      "01000011000110101101000100100110110110000001001111" when "1111101100",
      "01010010110011011000111000011101110100100101011111" when "1111101101",
      "01100010100001000011100001000001101010101011100111" when "1111101110",
      "01110010001111101101000010001101110010111101110111" when "1111101111",
      "00000001111111010101011111111101110111110100100101" when "1111110000",
      "00010001101111111100111110001101110011010111010011" when "1111110001",
      "00100001100001100011100000111001101111011101101010" when "1111110010",
      "00110001010100001001001011111110000101110000011011" when "1111110011",
      "01000001000111101110000011010111011111101010011100" when "1111110100",
      "01010000111100010010001011000010110110011001101001" when "1111110101",
      "01100000110001110101100110111101010011000000000001" when "1111110110",
      "01110000101000011000011011000100001110010100101001" when "1111110111",
      "00000000011111111010101011010101010001000100101000" when "1111111000",
      "00010000011000011100011011101110010011110100000110" when "1111111001",
      "00100000010001111101110000001101011110111111010001" when "1111111010",
      "00110000001100011110101100110001001010111011010100" when "1111111011",
      "01000000000111111111010101010111111111110111011110" when "1111111100",
      "01010000000100011111101110000000110101111101111110" when "1111111101",
      "01100000000001111111111010101010110101010101000100" when "1111111110",
      "01110000000000011111111111010101010101111111111111" when "1111111111",
      "--------------------------------------------------" when others;
   Y1_c4 <= Y0_c4; -- for the possible blockram register
   Y <= Y1_c4;
end architecture;

--------------------------------------------------------------------------------
--                       compressedTable_Freq300_uid52
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Luc Forget, Maxime Christ (2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity compressedTable_Freq300_uid52 is
    port (clk, ce_5 : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of compressedTable_Freq300_uid52 is
   component compressedTable_Freq300_uid52_subsampling_Freq300_uid54 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(8 downto 0)   );
   end component;

   component compressedTable_Freq300_uid52_diff_Freq300_uid57 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(49 downto 0)   );
   end component;

signal X_subsampling_c4 :  std_logic_vector(6 downto 0);
signal Y_subsampling_c4, Y_subsampling_c5 :  std_logic_vector(8 downto 0);
signal Y_subsampling_copy55_c4 :  std_logic_vector(8 downto 0);
signal Y_diff_c4, Y_diff_c5 :  std_logic_vector(49 downto 0);
signal fullOut_topbits_c5 :  std_logic_vector(8 downto 0);
signal fullOut_c5 :  std_logic_vector(56 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               Y_subsampling_c5 <= Y_subsampling_c4;
               Y_diff_c5 <= Y_diff_c4;
            end if;
         end if;
      end process;
   X_subsampling_c4 <= X(9 downto 3);
   compressedTable_Freq300_uid52_subsampling: compressedTable_Freq300_uid52_subsampling_Freq300_uid54
      port map ( X => X_subsampling_c4,
                 Y => Y_subsampling_copy55_c4);
   Y_subsampling_c4 <= Y_subsampling_copy55_c4; -- output copy to hold a pipeline register if needed
   compressedTable_Freq300_uid52_diff: compressedTable_Freq300_uid52_diff_Freq300_uid57
      port map ( clk  => clk,
                 X => X,
                 Y => Y_diff_c4);
   fullOut_topbits_c5 <= Y_subsampling_c5 + ("0000000"& (Y_diff_c5(49 downto 48)));
   fullOut_c5 <= fullOut_topbits_c5 & (Y_diff_c5(47 downto 0));
   Y <= fullOut_c5;
end architecture;

--------------------------------------------------------------------------------
--                      FixFunctionByTable_Freq300_uid50
-- Evaluator for exp(x*1b-1) on [-1,1) for lsbIn=-9 (wIn=10), msbout=0, lsbOut=-56 (wOut=57). Out interval: [0.606531; 1.64711]. Output is unsigned

-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq300_uid50 is
    port (clk, ce_5 : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq300_uid50 is
   component compressedTable_Freq300_uid52 is
      port ( clk, ce_5 : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(56 downto 0)   );
   end component;

begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
            end if;
         end if;
      end process;
   compressedTable: compressedTable_Freq300_uid52
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 X => X,
                 Y => Y);
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid69
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid69 is
    port (clk, ce_5 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid69 is
signal Mfull_c4, Mfull_c5 :  std_logic_vector(40 downto 0);
signal M_c5 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               Mfull_c5 <= Mfull_c4;
            end if;
         end if;
      end process;
   Mfull_c4 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c5 <= Mfull_c5(40 downto 0);
   R <= M_c5;
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid71
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid71 is
   component MultTable_Freq300_uid73 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy74_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid73
      port map ( X => Xtable_c4,
                 Y => Y1_copy74_c4);
   Y1_c4 <= Y1_copy74_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid76
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid76 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid76 is
   component MultTable_Freq300_uid78 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy79_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid78
      port map ( X => Xtable_c4,
                 Y => Y1_copy79_c4);
   Y1_c4 <= Y1_copy79_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid81
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid81 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid81 is
   component MultTable_Freq300_uid83 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy84_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid83
      port map ( X => Xtable_c4,
                 Y => Y1_copy84_c4);
   Y1_c4 <= Y1_copy84_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid86
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid86 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid86 is
   component MultTable_Freq300_uid88 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy89_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid88
      port map ( X => Xtable_c4,
                 Y => Y1_copy89_c4);
   Y1_c4 <= Y1_copy89_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid91
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid91 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid91 is
   component MultTable_Freq300_uid93 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy94_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid93
      port map ( X => Xtable_c4,
                 Y => Y1_copy94_c4);
   Y1_c4 <= Y1_copy94_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid96
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid96 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid96 is
   component MultTable_Freq300_uid98 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy99_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid98
      port map ( X => Xtable_c4,
                 Y => Y1_copy99_c4);
   Y1_c4 <= Y1_copy99_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid101
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid101 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid101 is
   component MultTable_Freq300_uid103 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy104_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid103
      port map ( X => Xtable_c4,
                 Y => Y1_copy104_c4);
   Y1_c4 <= Y1_copy104_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid106
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid106 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid106 is
   component MultTable_Freq300_uid108 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy109_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid108
      port map ( X => Xtable_c4,
                 Y => Y1_copy109_c4);
   Y1_c4 <= Y1_copy109_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid111
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid111 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid111 is
   component MultTable_Freq300_uid113 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy114_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid113
      port map ( X => Xtable_c4,
                 Y => Y1_copy114_c4);
   Y1_c4 <= Y1_copy114_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid116
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid116 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid116 is
   component MultTable_Freq300_uid118 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy119_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid118
      port map ( X => Xtable_c4,
                 Y => Y1_copy119_c4);
   Y1_c4 <= Y1_copy119_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid121
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid121 is
   component MultTable_Freq300_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy124_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid123
      port map ( X => Xtable_c4,
                 Y => Y1_copy124_c4);
   Y1_c4 <= Y1_copy124_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid126
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid126 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid126 is
   component MultTable_Freq300_uid128 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy129_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid128
      port map ( X => Xtable_c4,
                 Y => Y1_copy129_c4);
   Y1_c4 <= Y1_copy129_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid131
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid131 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid131 is
   component MultTable_Freq300_uid133 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy134_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid133
      port map ( X => Xtable_c4,
                 Y => Y1_copy134_c4);
   Y1_c4 <= Y1_copy134_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid136
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid136 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid136 is
   component MultTable_Freq300_uid138 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy139_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid138
      port map ( X => Xtable_c4,
                 Y => Y1_copy139_c4);
   Y1_c4 <= Y1_copy139_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid141
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid141 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid141 is
   component MultTable_Freq300_uid143 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy144_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid143
      port map ( X => Xtable_c4,
                 Y => Y1_copy144_c4);
   Y1_c4 <= Y1_copy144_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid146
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid146 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid146 is
   component MultTable_Freq300_uid148 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy149_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid148
      port map ( X => Xtable_c4,
                 Y => Y1_copy149_c4);
   Y1_c4 <= Y1_copy149_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid151
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid151 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid151 is
   component MultTable_Freq300_uid153 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy154_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid153
      port map ( X => Xtable_c4,
                 Y => Y1_copy154_c4);
   Y1_c4 <= Y1_copy154_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid156
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid156 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid156 is
   component MultTable_Freq300_uid158 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy159_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid158
      port map ( X => Xtable_c4,
                 Y => Y1_copy159_c4);
   Y1_c4 <= Y1_copy159_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid161
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid161 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid161 is
   component MultTable_Freq300_uid163 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy164_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid163
      port map ( X => Xtable_c4,
                 Y => Y1_copy164_c4);
   Y1_c4 <= Y1_copy164_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid166
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid166 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid166 is
   component MultTable_Freq300_uid168 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy169_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid168
      port map ( X => Xtable_c4,
                 Y => Y1_copy169_c4);
   Y1_c4 <= Y1_copy169_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid171
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid171 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid171 is
   component MultTable_Freq300_uid173 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy174_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid173
      port map ( X => Xtable_c4,
                 Y => Y1_copy174_c4);
   Y1_c4 <= Y1_copy174_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid176
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid176 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid176 is
   component MultTable_Freq300_uid178 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy179_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid178
      port map ( X => Xtable_c4,
                 Y => Y1_copy179_c4);
   Y1_c4 <= Y1_copy179_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid181
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid181 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid181 is
   component MultTable_Freq300_uid183 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy184_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid183
      port map ( X => Xtable_c4,
                 Y => Y1_copy184_c4);
   Y1_c4 <= Y1_copy184_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid186
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid186 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid186 is
   component MultTable_Freq300_uid188 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy189_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid188
      port map ( X => Xtable_c4,
                 Y => Y1_copy189_c4);
   Y1_c4 <= Y1_copy189_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid191
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid191 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid191 is
   component MultTable_Freq300_uid193 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy194_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid193
      port map ( X => Xtable_c4,
                 Y => Y1_copy194_c4);
   Y1_c4 <= Y1_copy194_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid196
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid196 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid196 is
   component MultTable_Freq300_uid198 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy199_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid198
      port map ( X => Xtable_c4,
                 Y => Y1_copy199_c4);
   Y1_c4 <= Y1_copy199_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid201
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid201 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid201 is
   component MultTable_Freq300_uid203 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy204_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid203
      port map ( X => Xtable_c4,
                 Y => Y1_copy204_c4);
   Y1_c4 <= Y1_copy204_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid206
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid206 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid206 is
   component MultTable_Freq300_uid208 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy209_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid208
      port map ( X => Xtable_c4,
                 Y => Y1_copy209_c4);
   Y1_c4 <= Y1_copy209_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid211
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid211 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid211 is
   component MultTable_Freq300_uid213 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy214_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid213
      port map ( X => Xtable_c4,
                 Y => Y1_copy214_c4);
   Y1_c4 <= Y1_copy214_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid216
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid216 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid216 is
   component MultTable_Freq300_uid218 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy219_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid218
      port map ( X => Xtable_c4,
                 Y => Y1_copy219_c4);
   Y1_c4 <= Y1_copy219_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid221
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid221 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid221 is
   component MultTable_Freq300_uid223 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy224_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid223
      port map ( X => Xtable_c4,
                 Y => Y1_copy224_c4);
   Y1_c4 <= Y1_copy224_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid226
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid226 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid226 is
   component MultTable_Freq300_uid228 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy229_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid228
      port map ( X => Xtable_c4,
                 Y => Y1_copy229_c4);
   Y1_c4 <= Y1_copy229_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid231
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid231 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid231 is
   component MultTable_Freq300_uid233 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy234_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid233
      port map ( X => Xtable_c4,
                 Y => Y1_copy234_c4);
   Y1_c4 <= Y1_copy234_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_2_signedx2_Freq300_uid236
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2_signedx2_Freq300_uid236 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2_signedx2_Freq300_uid236 is
   component MultTable_Freq300_uid238 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(3 downto 0);
signal Y1_c4 :  std_logic_vector(3 downto 0);
signal Y1_copy239_c4 :  std_logic_vector(3 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid238
      port map ( X => Xtable_c4,
                 Y => Y1_copy239_c4);
   Y1_c4 <= Y1_copy239_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid241
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid241 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid241 is
   component MultTable_Freq300_uid243 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy244_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid243
      port map ( X => Xtable_c4,
                 Y => Y1_copy244_c4);
   Y1_c4 <= Y1_copy244_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid246
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid246 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid246 is
   component MultTable_Freq300_uid248 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy249_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid248
      port map ( X => Xtable_c4,
                 Y => Y1_copy249_c4);
   Y1_c4 <= Y1_copy249_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_1x1_signed_Freq300_uid251
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_signed_Freq300_uid251 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_signed_Freq300_uid251 is
signal replicated_c4 :  std_logic_vector(0 downto 0);
signal prod_c4 :  std_logic_vector(0 downto 0);
begin
   replicated_c4 <= (0 downto 0 => X(0));
   prod_c4 <= Y and replicated_c4;
   R <= prod_c4;
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid253
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid253 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid253 is
   component MultTable_Freq300_uid255 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy256_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid255
      port map ( X => Xtable_c4,
                 Y => Y1_copy256_c4);
   Y1_c4 <= Y1_copy256_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid258
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid258 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid258 is
   component MultTable_Freq300_uid260 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy261_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid260
      port map ( X => Xtable_c4,
                 Y => Y1_copy261_c4);
   Y1_c4 <= Y1_copy261_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid263
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid263 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid263 is
   component MultTable_Freq300_uid265 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy266_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid265
      port map ( X => Xtable_c4,
                 Y => Y1_copy266_c4);
   Y1_c4 <= Y1_copy266_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid268
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid268 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid268 is
   component MultTable_Freq300_uid270 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy271_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid270
      port map ( X => Xtable_c4,
                 Y => Y1_copy271_c4);
   Y1_c4 <= Y1_copy271_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--             IntMultiplierLUT_4_signedx1_signed_Freq300_uid273
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4_signedx1_signed_Freq300_uid273 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4_signedx1_signed_Freq300_uid273 is
   component MultTable_Freq300_uid275 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy276_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid275
      port map ( X => Xtable_c4,
                 Y => Y1_copy276_c4);
   Y1_c4 <= Y1_copy276_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid278
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid278 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid278 is
   component MultTable_Freq300_uid280 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c4 :  std_logic_vector(4 downto 0);
signal Y1_c4 :  std_logic_vector(4 downto 0);
signal Y1_copy281_c4 :  std_logic_vector(4 downto 0);
begin
Xtable_c4 <= Y & X;
   R <= Y1_c4;
   TableMult: MultTable_Freq300_uid280
      port map ( X => Xtable_c4,
                 Y => Y1_copy281_c4);
   Y1_c4 <= Y1_copy281_c4; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_Freq300_uid534
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_Freq300_uid534 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(32 downto 0);
          Y : in  std_logic_vector(32 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_Freq300_uid534 is
signal Rtmp_c6 :  std_logic_vector(32 downto 0);
signal X_c6 :  std_logic_vector(32 downto 0);
signal Y_c6 :  std_logic_vector(32 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               X_c6 <= X;
               Y_c6 <= Y;
               Cin_c6 <= Cin_c5;
            end if;
         end if;
      end process;
   Rtmp_c6 <= X_c6 + Y_c6 + Cin_c6;
   R <= Rtmp_c6;
end architecture;

--------------------------------------------------------------------------------
--    FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid66
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Matei Istoan, 2012-2014, 2024
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y A
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid66 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(24 downto 0);
          Y : in  std_logic_vector(24 downto 0);
          A : in  std_logic_vector(32 downto 0);
          R : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid66 is
   component DSPBlock_17x24_Freq300_uid69 is
      port ( clk, ce_5 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid76 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid81 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid86 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid91 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid96 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid101 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid106 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid111 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid116 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid126 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid131 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid136 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid141 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid146 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid151 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid156 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid161 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid166 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid171 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid176 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid181 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid186 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid191 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid196 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid201 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid206 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid211 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid216 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid221 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid226 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid231 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2_signedx2_Freq300_uid236 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid241 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid246 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_signed_Freq300_uid251 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid253 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid258 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid263 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid268 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4_signedx1_signed_Freq300_uid273 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid278 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid284 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid288 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid292 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid300 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq300_uid334 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_33_Freq300_uid534 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(32 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(32 downto 0)   );
   end component;

signal XX_c4 :  signed(0+24 downto 0);
signal YY_c4 :  signed(-17+41 downto 0);
signal AA_c4 :  signed(-9+41 downto 0);
signal tile_0_X_c4 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c4 :  std_logic_vector(23 downto 0);
signal tile_0_output_c5 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c5 :  unsigned(40-0 downto 0);
signal bh67_wm65_0_c5 :  std_logic;
signal bh67_wm64_0_c5 :  std_logic;
signal bh67_wm63_0_c5 :  std_logic;
signal bh67_wm62_0_c5 :  std_logic;
signal bh67_wm61_0_c5 :  std_logic;
signal bh67_wm60_0_c5 :  std_logic;
signal bh67_wm59_0_c5 :  std_logic;
signal bh67_wm58_0_c5 :  std_logic;
signal bh67_wm57_0_c5 :  std_logic;
signal bh67_wm56_0_c5 :  std_logic;
signal bh67_wm55_0_c5 :  std_logic;
signal bh67_wm54_0_c5 :  std_logic;
signal bh67_wm53_0_c5 :  std_logic;
signal bh67_wm52_0_c5 :  std_logic;
signal bh67_wm51_0_c5 :  std_logic;
signal bh67_wm50_0_c5 :  std_logic;
signal bh67_wm49_0_c5 :  std_logic;
signal bh67_wm48_0_c5 :  std_logic;
signal bh67_wm47_0_c5 :  std_logic;
signal bh67_wm46_0_c5 :  std_logic;
signal bh67_wm45_0_c5 :  std_logic;
signal bh67_wm44_0_c5 :  std_logic;
signal bh67_wm43_0_c5 :  std_logic;
signal bh67_wm42_0_c5 :  std_logic;
signal bh67_wm41_0_c5 :  std_logic;
signal bh67_wm40_0_c5 :  std_logic;
signal bh67_wm39_0_c5 :  std_logic;
signal bh67_wm38_0_c5 :  std_logic;
signal bh67_wm37_0_c5 :  std_logic;
signal bh67_wm36_0_c5 :  std_logic;
signal bh67_wm35_0_c5 :  std_logic;
signal bh67_wm34_0_c5 :  std_logic;
signal bh67_wm33_0_c5 :  std_logic;
signal bh67_wm32_0_c5 :  std_logic;
signal bh67_wm31_0_c5 :  std_logic;
signal bh67_wm30_0_c5 :  std_logic;
signal bh67_wm29_0_c5 :  std_logic;
signal bh67_wm28_0_c5 :  std_logic;
signal bh67_wm27_0_c5 :  std_logic;
signal bh67_wm26_0_c5 :  std_logic;
signal bh67_wm25_0_c5 :  std_logic;
signal tile_1_X_c4 :  std_logic_vector(1 downto 0);
signal tile_1_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_1_output_c4 :  std_logic_vector(3 downto 0);
signal tile_1_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm20_0_c4 :  std_logic;
signal bh67_wm19_0_c4 :  std_logic;
signal bh67_wm18_0_c4 :  std_logic;
signal bh67_wm17_0_c4 :  std_logic;
signal tile_2_X_c4 :  std_logic_vector(2 downto 0);
signal tile_2_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_2_output_c4 :  std_logic_vector(4 downto 0);
signal tile_2_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm23_0_c4 :  std_logic;
signal bh67_wm22_0_c4 :  std_logic;
signal bh67_wm21_0_c4 :  std_logic;
signal bh67_wm20_1_c4 :  std_logic;
signal bh67_wm19_1_c4 :  std_logic;
signal tile_3_X_c4 :  std_logic_vector(2 downto 0);
signal tile_3_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_3_output_c4 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm26_1_c4, bh67_wm26_1_c5 :  std_logic;
signal bh67_wm25_1_c4 :  std_logic;
signal bh67_wm24_0_c4 :  std_logic;
signal bh67_wm23_1_c4 :  std_logic;
signal bh67_wm22_1_c4 :  std_logic;
signal tile_4_X_c4 :  std_logic_vector(1 downto 0);
signal tile_4_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_4_output_c4 :  std_logic_vector(3 downto 0);
signal tile_4_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm22_2_c4 :  std_logic;
signal bh67_wm21_1_c4 :  std_logic;
signal bh67_wm20_2_c4 :  std_logic;
signal bh67_wm19_2_c4 :  std_logic;
signal tile_5_X_c4 :  std_logic_vector(2 downto 0);
signal tile_5_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_5_output_c4 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm25_2_c4 :  std_logic;
signal bh67_wm24_1_c4 :  std_logic;
signal bh67_wm23_2_c4 :  std_logic;
signal bh67_wm22_3_c4 :  std_logic;
signal bh67_wm21_2_c4 :  std_logic;
signal tile_6_X_c4 :  std_logic_vector(2 downto 0);
signal tile_6_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_6_output_c4 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm28_1_c4, bh67_wm28_1_c5 :  std_logic;
signal bh67_wm27_1_c4 :  std_logic;
signal bh67_wm26_2_c4, bh67_wm26_2_c5 :  std_logic;
signal bh67_wm25_3_c4 :  std_logic;
signal bh67_wm24_2_c4 :  std_logic;
signal tile_7_X_c4 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_7_output_c4 :  std_logic_vector(3 downto 0);
signal tile_7_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm24_3_c4 :  std_logic;
signal bh67_wm23_3_c4 :  std_logic;
signal bh67_wm22_4_c4 :  std_logic;
signal bh67_wm21_3_c4 :  std_logic;
signal tile_8_X_c4 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_8_output_c4 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm27_2_c4 :  std_logic;
signal bh67_wm26_3_c4, bh67_wm26_3_c5 :  std_logic;
signal bh67_wm25_4_c4 :  std_logic;
signal bh67_wm24_4_c4 :  std_logic;
signal bh67_wm23_4_c4 :  std_logic;
signal tile_9_X_c4 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_9_output_c4 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm30_1_c4, bh67_wm30_1_c5 :  std_logic;
signal bh67_wm29_1_c4, bh67_wm29_1_c5 :  std_logic;
signal bh67_wm28_2_c4, bh67_wm28_2_c5 :  std_logic;
signal bh67_wm27_3_c4 :  std_logic;
signal bh67_wm26_4_c4, bh67_wm26_4_c5 :  std_logic;
signal tile_10_X_c4 :  std_logic_vector(1 downto 0);
signal tile_10_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_10_output_c4 :  std_logic_vector(3 downto 0);
signal tile_10_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm26_5_c4, bh67_wm26_5_c5 :  std_logic;
signal bh67_wm25_5_c4 :  std_logic;
signal bh67_wm24_5_c4 :  std_logic;
signal bh67_wm23_5_c4 :  std_logic;
signal tile_11_X_c4 :  std_logic_vector(2 downto 0);
signal tile_11_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_11_output_c4 :  std_logic_vector(4 downto 0);
signal tile_11_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm29_2_c4, bh67_wm29_2_c5 :  std_logic;
signal bh67_wm28_3_c4, bh67_wm28_3_c5 :  std_logic;
signal bh67_wm27_4_c4 :  std_logic;
signal bh67_wm26_6_c4 :  std_logic;
signal bh67_wm25_6_c4 :  std_logic;
signal tile_12_X_c4 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_12_output_c4 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm32_1_c4, bh67_wm32_1_c5 :  std_logic;
signal bh67_wm31_1_c4 :  std_logic;
signal bh67_wm30_2_c4, bh67_wm30_2_c5 :  std_logic;
signal bh67_wm29_3_c4, bh67_wm29_3_c5 :  std_logic;
signal bh67_wm28_4_c4, bh67_wm28_4_c5 :  std_logic;
signal tile_13_X_c4 :  std_logic_vector(1 downto 0);
signal tile_13_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_13_output_c4 :  std_logic_vector(3 downto 0);
signal tile_13_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm28_5_c4, bh67_wm28_5_c5 :  std_logic;
signal bh67_wm27_5_c4 :  std_logic;
signal bh67_wm26_7_c4 :  std_logic;
signal bh67_wm25_7_c4 :  std_logic;
signal tile_14_X_c4 :  std_logic_vector(2 downto 0);
signal tile_14_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_14_output_c4 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm31_2_c4 :  std_logic;
signal bh67_wm30_3_c4, bh67_wm30_3_c5 :  std_logic;
signal bh67_wm29_4_c4, bh67_wm29_4_c5 :  std_logic;
signal bh67_wm28_6_c4 :  std_logic;
signal bh67_wm27_6_c4 :  std_logic;
signal tile_15_X_c4 :  std_logic_vector(2 downto 0);
signal tile_15_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_15_output_c4 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm34_1_c4, bh67_wm34_1_c5 :  std_logic;
signal bh67_wm33_1_c4, bh67_wm33_1_c5 :  std_logic;
signal bh67_wm32_2_c4, bh67_wm32_2_c5 :  std_logic;
signal bh67_wm31_3_c4 :  std_logic;
signal bh67_wm30_4_c4, bh67_wm30_4_c5 :  std_logic;
signal tile_16_X_c4 :  std_logic_vector(1 downto 0);
signal tile_16_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_16_output_c4 :  std_logic_vector(3 downto 0);
signal tile_16_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm30_5_c4, bh67_wm30_5_c5 :  std_logic;
signal bh67_wm29_5_c4, bh67_wm29_5_c5 :  std_logic;
signal bh67_wm28_7_c4 :  std_logic;
signal bh67_wm27_7_c4 :  std_logic;
signal tile_17_X_c4 :  std_logic_vector(2 downto 0);
signal tile_17_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_17_output_c4 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm33_2_c4, bh67_wm33_2_c5 :  std_logic;
signal bh67_wm32_3_c4, bh67_wm32_3_c5 :  std_logic;
signal bh67_wm31_4_c4 :  std_logic;
signal bh67_wm30_6_c4 :  std_logic;
signal bh67_wm29_6_c4 :  std_logic;
signal tile_18_X_c4 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_18_output_c4 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm36_1_c4, bh67_wm36_1_c5 :  std_logic;
signal bh67_wm35_1_c4 :  std_logic;
signal bh67_wm34_2_c4, bh67_wm34_2_c5 :  std_logic;
signal bh67_wm33_3_c4, bh67_wm33_3_c5 :  std_logic;
signal bh67_wm32_4_c4, bh67_wm32_4_c5 :  std_logic;
signal tile_19_X_c4 :  std_logic_vector(1 downto 0);
signal tile_19_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_19_output_c4 :  std_logic_vector(3 downto 0);
signal tile_19_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm32_5_c4, bh67_wm32_5_c5 :  std_logic;
signal bh67_wm31_5_c4 :  std_logic;
signal bh67_wm30_7_c4 :  std_logic;
signal bh67_wm29_7_c4 :  std_logic;
signal tile_20_X_c4 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_20_output_c4 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm35_2_c4 :  std_logic;
signal bh67_wm34_3_c4, bh67_wm34_3_c5 :  std_logic;
signal bh67_wm33_4_c4, bh67_wm33_4_c5 :  std_logic;
signal bh67_wm32_6_c4 :  std_logic;
signal bh67_wm31_6_c4 :  std_logic;
signal tile_21_X_c4 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_21_output_c4 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm38_1_c4 :  std_logic;
signal bh67_wm37_1_c4, bh67_wm37_1_c5 :  std_logic;
signal bh67_wm36_2_c4, bh67_wm36_2_c5 :  std_logic;
signal bh67_wm35_3_c4 :  std_logic;
signal bh67_wm34_4_c4, bh67_wm34_4_c5 :  std_logic;
signal tile_22_X_c4 :  std_logic_vector(1 downto 0);
signal tile_22_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_22_output_c4 :  std_logic_vector(3 downto 0);
signal tile_22_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm34_5_c4, bh67_wm34_5_c5 :  std_logic;
signal bh67_wm33_5_c4, bh67_wm33_5_c5 :  std_logic;
signal bh67_wm32_7_c4 :  std_logic;
signal bh67_wm31_7_c4 :  std_logic;
signal tile_23_X_c4 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_23_output_c4 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm37_2_c4, bh67_wm37_2_c5 :  std_logic;
signal bh67_wm36_3_c4, bh67_wm36_3_c5 :  std_logic;
signal bh67_wm35_4_c4 :  std_logic;
signal bh67_wm34_6_c4 :  std_logic;
signal bh67_wm33_6_c4 :  std_logic;
signal tile_24_X_c4 :  std_logic_vector(2 downto 0);
signal tile_24_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_24_output_c4 :  std_logic_vector(4 downto 0);
signal tile_24_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm40_1_c4, bh67_wm40_1_c5 :  std_logic;
signal bh67_wm39_1_c4 :  std_logic;
signal bh67_wm38_2_c4 :  std_logic;
signal bh67_wm37_3_c4, bh67_wm37_3_c5 :  std_logic;
signal bh67_wm36_4_c4, bh67_wm36_4_c5 :  std_logic;
signal tile_25_X_c4 :  std_logic_vector(1 downto 0);
signal tile_25_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_25_output_c4 :  std_logic_vector(3 downto 0);
signal tile_25_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm36_5_c4, bh67_wm36_5_c5 :  std_logic;
signal bh67_wm35_5_c4 :  std_logic;
signal bh67_wm34_7_c4 :  std_logic;
signal bh67_wm33_7_c4 :  std_logic;
signal tile_26_X_c4 :  std_logic_vector(2 downto 0);
signal tile_26_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_26_output_c4 :  std_logic_vector(4 downto 0);
signal tile_26_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm39_2_c4 :  std_logic;
signal bh67_wm38_3_c4 :  std_logic;
signal bh67_wm37_4_c4, bh67_wm37_4_c5 :  std_logic;
signal bh67_wm36_6_c4 :  std_logic;
signal bh67_wm35_6_c4 :  std_logic;
signal tile_27_X_c4 :  std_logic_vector(2 downto 0);
signal tile_27_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_27_output_c4 :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm42_1_c4 :  std_logic;
signal bh67_wm41_1_c4, bh67_wm41_1_c5 :  std_logic;
signal bh67_wm40_2_c4, bh67_wm40_2_c5 :  std_logic;
signal bh67_wm39_3_c4 :  std_logic;
signal bh67_wm38_4_c4 :  std_logic;
signal tile_28_X_c4 :  std_logic_vector(1 downto 0);
signal tile_28_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_28_output_c4 :  std_logic_vector(3 downto 0);
signal tile_28_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm38_5_c4 :  std_logic;
signal bh67_wm37_5_c4, bh67_wm37_5_c5 :  std_logic;
signal bh67_wm36_7_c4 :  std_logic;
signal bh67_wm35_7_c4 :  std_logic;
signal tile_29_X_c4 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_29_output_c4 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm41_2_c4, bh67_wm41_2_c5 :  std_logic;
signal bh67_wm40_3_c4, bh67_wm40_3_c5 :  std_logic;
signal bh67_wm39_4_c4 :  std_logic;
signal bh67_wm38_6_c4 :  std_logic;
signal bh67_wm37_6_c4 :  std_logic;
signal tile_30_X_c4 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_30_output_c4 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm44_1_c4 :  std_logic;
signal bh67_wm43_1_c4 :  std_logic;
signal bh67_wm42_2_c4 :  std_logic;
signal bh67_wm41_3_c4, bh67_wm41_3_c5 :  std_logic;
signal bh67_wm40_4_c4, bh67_wm40_4_c5 :  std_logic;
signal tile_31_X_c4 :  std_logic_vector(1 downto 0);
signal tile_31_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_31_output_c4 :  std_logic_vector(3 downto 0);
signal tile_31_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm40_5_c4, bh67_wm40_5_c5 :  std_logic;
signal bh67_wm39_5_c4 :  std_logic;
signal bh67_wm38_7_c4 :  std_logic;
signal bh67_wm37_7_c4 :  std_logic;
signal tile_32_X_c4 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_32_output_c4 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm43_2_c4 :  std_logic;
signal bh67_wm42_3_c4 :  std_logic;
signal bh67_wm41_4_c4, bh67_wm41_4_c5 :  std_logic;
signal bh67_wm40_6_c4 :  std_logic;
signal bh67_wm39_6_c4 :  std_logic;
signal tile_33_X_c4 :  std_logic_vector(2 downto 0);
signal tile_33_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_33_output_c4 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm46_1_c4, bh67_wm46_1_c5 :  std_logic;
signal bh67_wm45_1_c4, bh67_wm45_1_c5 :  std_logic;
signal bh67_wm44_2_c4 :  std_logic;
signal bh67_wm43_3_c4 :  std_logic;
signal bh67_wm42_4_c4 :  std_logic;
signal tile_34_X_c4 :  std_logic_vector(1 downto 0);
signal tile_34_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_34_output_c4 :  std_logic_vector(3 downto 0);
signal tile_34_filtered_output_c4 :  signed(3-0 downto 0);
signal bh67_wm42_5_c4 :  std_logic;
signal bh67_wm41_5_c4, bh67_wm41_5_c5 :  std_logic;
signal bh67_wm40_7_c4 :  std_logic;
signal bh67_wm39_7_c4 :  std_logic;
signal tile_35_X_c4 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_35_output_c4 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm45_2_c4, bh67_wm45_2_c5 :  std_logic;
signal bh67_wm44_3_c4 :  std_logic;
signal bh67_wm43_4_c4 :  std_logic;
signal bh67_wm42_6_c4 :  std_logic;
signal bh67_wm41_6_c4 :  std_logic;
signal tile_36_X_c4 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c4 :  std_logic_vector(1 downto 0);
signal tile_36_output_c4 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c4 :  unsigned(4-0 downto 0);
signal bh67_wm48_1_c4, bh67_wm48_1_c5 :  std_logic;
signal bh67_wm47_1_c4, bh67_wm47_1_c5 :  std_logic;
signal bh67_wm46_2_c4, bh67_wm46_2_c5 :  std_logic;
signal bh67_wm45_3_c4, bh67_wm45_3_c5 :  std_logic;
signal bh67_wm44_4_c4 :  std_logic;
signal tile_37_X_c4 :  std_logic_vector(0 downto 0);
signal tile_37_Y_c4 :  std_logic_vector(0 downto 0);
signal tile_37_output_c4 :  std_logic_vector(0 downto 0);
signal tile_37_filtered_output_c4 :  signed(0-0 downto 0);
signal bh67_wm25_8_c4 :  std_logic;
signal tile_38_X_c4 :  std_logic_vector(3 downto 0);
signal tile_38_Y_c4 :  std_logic_vector(0 downto 0);
signal tile_38_output_c4 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c4 :  signed(4-0 downto 0);
signal bh67_wm29_8_c4 :  std_logic;
signal bh67_wm28_8_c4 :  std_logic;
signal bh67_wm27_8_c4 :  std_logic;
signal bh67_wm26_8_c4 :  std_logic;
signal bh67_wm25_9_c4 :  std_logic;
signal tile_39_X_c4 :  std_logic_vector(3 downto 0);
signal tile_39_Y_c4 :  std_logic_vector(0 downto 0);
signal tile_39_output_c4 :  std_logic_vector(4 downto 0);
signal tile_39_filtered_output_c4 :  signed(4-0 downto 0);
signal bh67_wm33_8_c4 :  std_logic;
signal bh67_wm32_8_c4 :  std_logic;
signal bh67_wm31_8_c4 :  std_logic;
signal bh67_wm30_8_c4 :  std_logic;
signal bh67_wm29_9_c4 :  std_logic;
signal tile_40_X_c4 :  std_logic_vector(3 downto 0);
signal tile_40_Y_c4 :  std_logic_vector(0 downto 0);
signal tile_40_output_c4 :  std_logic_vector(4 downto 0);
signal tile_40_filtered_output_c4 :  signed(4-0 downto 0);
signal bh67_wm37_8_c4 :  std_logic;
signal bh67_wm36_8_c4 :  std_logic;
signal bh67_wm35_8_c4 :  std_logic;
signal bh67_wm34_8_c4 :  std_logic;
signal bh67_wm33_9_c4 :  std_logic;
signal tile_41_X_c4 :  std_logic_vector(3 downto 0);
signal tile_41_Y_c4 :  std_logic_vector(0 downto 0);
signal tile_41_output_c4 :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output_c4 :  signed(4-0 downto 0);
signal bh67_wm41_7_c4 :  std_logic;
signal bh67_wm40_8_c4 :  std_logic;
signal bh67_wm39_8_c4 :  std_logic;
signal bh67_wm38_8_c4 :  std_logic;
signal bh67_wm37_9_c4 :  std_logic;
signal tile_42_X_c4 :  std_logic_vector(3 downto 0);
signal tile_42_Y_c4 :  std_logic_vector(0 downto 0);
signal tile_42_output_c4 :  std_logic_vector(4 downto 0);
signal tile_42_filtered_output_c4 :  signed(4-0 downto 0);
signal bh67_wm20_3_c4 :  std_logic;
signal bh67_wm19_3_c4 :  std_logic;
signal bh67_wm18_1_c4 :  std_logic;
signal bh67_wm17_1_c4 :  std_logic;
signal bh67_wm16_0_c4 :  std_logic;
signal tile_43_X_c4 :  std_logic_vector(3 downto 0);
signal tile_43_Y_c4 :  std_logic_vector(0 downto 0);
signal tile_43_output_c4 :  std_logic_vector(4 downto 0);
signal tile_43_filtered_output_c4 :  signed(4-0 downto 0);
signal bh67_wm24_6_c4 :  std_logic;
signal bh67_wm23_6_c4 :  std_logic;
signal bh67_wm22_5_c4 :  std_logic;
signal bh67_wm21_4_c4 :  std_logic;
signal bh67_wm20_4_c4 :  std_logic;
signal bh67_wm41_8_c4 :  std_logic;
signal bh67_wm40_9_c4 :  std_logic;
signal bh67_wm39_9_c4 :  std_logic;
signal bh67_wm38_9_c4 :  std_logic;
signal bh67_wm37_10_c4 :  std_logic;
signal bh67_wm36_9_c4 :  std_logic;
signal bh67_wm35_9_c4 :  std_logic;
signal bh67_wm34_9_c4 :  std_logic;
signal bh67_wm33_10_c4 :  std_logic;
signal bh67_wm32_9_c4 :  std_logic;
signal bh67_wm31_9_c4 :  std_logic;
signal bh67_wm30_9_c4 :  std_logic;
signal bh67_wm29_10_c4 :  std_logic;
signal bh67_wm28_9_c4 :  std_logic;
signal bh67_wm27_9_c4 :  std_logic;
signal bh67_wm26_9_c4 :  std_logic;
signal bh67_wm25_10_c4 :  std_logic;
signal bh67_wm24_7_c4, bh67_wm24_7_c5 :  std_logic;
signal bh67_wm23_7_c4 :  std_logic;
signal bh67_wm22_6_c4 :  std_logic;
signal bh67_wm21_5_c4 :  std_logic;
signal bh67_wm20_5_c4 :  std_logic;
signal bh67_wm19_4_c4 :  std_logic;
signal bh67_wm18_2_c4 :  std_logic;
signal bh67_wm17_2_c4 :  std_logic;
signal bh67_wm16_1_c4 :  std_logic;
signal bh67_wm15_0_c4 :  std_logic;
signal bh67_wm14_0_c4 :  std_logic;
signal bh67_wm13_0_c4 :  std_logic;
signal bh67_wm12_0_c4 :  std_logic;
signal bh67_wm11_0_c4 :  std_logic;
signal bh67_wm10_0_c4 :  std_logic;
signal bh67_wm9_0_c4 :  std_logic;
signal bh67_wm42_7_c0, bh67_wm42_7_c1, bh67_wm42_7_c2, bh67_wm42_7_c3, bh67_wm42_7_c4, bh67_wm42_7_c5 :  std_logic;
signal bh67_wm39_10_c0, bh67_wm39_10_c1, bh67_wm39_10_c2, bh67_wm39_10_c3, bh67_wm39_10_c4 :  std_logic;
signal bh67_wm38_10_c0, bh67_wm38_10_c1, bh67_wm38_10_c2, bh67_wm38_10_c3, bh67_wm38_10_c4, bh67_wm38_10_c5 :  std_logic;
signal bh67_wm37_11_c0, bh67_wm37_11_c1, bh67_wm37_11_c2, bh67_wm37_11_c3, bh67_wm37_11_c4 :  std_logic;
signal bh67_wm34_10_c0, bh67_wm34_10_c1, bh67_wm34_10_c2, bh67_wm34_10_c3, bh67_wm34_10_c4 :  std_logic;
signal bh67_wm33_11_c0, bh67_wm33_11_c1, bh67_wm33_11_c2, bh67_wm33_11_c3, bh67_wm33_11_c4 :  std_logic;
signal bh67_wm30_10_c0, bh67_wm30_10_c1, bh67_wm30_10_c2, bh67_wm30_10_c3, bh67_wm30_10_c4 :  std_logic;
signal bh67_wm29_11_c0, bh67_wm29_11_c1, bh67_wm29_11_c2, bh67_wm29_11_c3, bh67_wm29_11_c4 :  std_logic;
signal bh67_wm26_10_c0, bh67_wm26_10_c1, bh67_wm26_10_c2, bh67_wm26_10_c3, bh67_wm26_10_c4, bh67_wm26_10_c5 :  std_logic;
signal bh67_wm22_7_c0, bh67_wm22_7_c1, bh67_wm22_7_c2, bh67_wm22_7_c3, bh67_wm22_7_c4 :  std_logic;
signal bh67_wm18_3_c0, bh67_wm18_3_c1, bh67_wm18_3_c2, bh67_wm18_3_c3, bh67_wm18_3_c4 :  std_logic;
signal bh67_wm15_1_c0, bh67_wm15_1_c1, bh67_wm15_1_c2, bh67_wm15_1_c3, bh67_wm15_1_c4 :  std_logic;
signal bh67_wm14_1_c0, bh67_wm14_1_c1, bh67_wm14_1_c2, bh67_wm14_1_c3, bh67_wm14_1_c4 :  std_logic;
signal bh67_wm13_1_c0, bh67_wm13_1_c1, bh67_wm13_1_c2, bh67_wm13_1_c3, bh67_wm13_1_c4 :  std_logic;
signal bh67_wm12_1_c0, bh67_wm12_1_c1, bh67_wm12_1_c2, bh67_wm12_1_c3, bh67_wm12_1_c4 :  std_logic;
signal bh67_wm11_1_c0, bh67_wm11_1_c1, bh67_wm11_1_c2, bh67_wm11_1_c3, bh67_wm11_1_c4 :  std_logic;
signal bh67_wm10_1_c0, bh67_wm10_1_c1, bh67_wm10_1_c2, bh67_wm10_1_c3, bh67_wm10_1_c4 :  std_logic;
signal bh67_wm9_1_c0, bh67_wm9_1_c1, bh67_wm9_1_c2, bh67_wm9_1_c3, bh67_wm9_1_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid285_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid285_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid285_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm48_2_c5 :  std_logic;
signal bh67_wm47_2_c5 :  std_logic;
signal bh67_wm46_3_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid285_Out0_copy286_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid289_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid289_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm46_4_c5 :  std_logic;
signal bh67_wm45_4_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid289_Out0_copy290_c5 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid293_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid293_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid293_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm45_5_c5 :  std_logic;
signal bh67_wm44_5_c5 :  std_logic;
signal bh67_wm43_5_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid293_Out0_copy294_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid295_In0_c4, Compressor_14_3_Freq300_uid292_bh67_uid295_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid295_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid295_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm44_6_c5 :  std_logic;
signal bh67_wm43_6_c5 :  std_logic;
signal bh67_wm42_8_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid295_Out0_copy296_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid297_In0_c4, Compressor_14_3_Freq300_uid292_bh67_uid297_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid297_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid297_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm43_7_c5 :  std_logic;
signal bh67_wm42_9_c5 :  std_logic;
signal bh67_wm41_9_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid297_Out0_copy298_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid301_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid301_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm42_10_c4, bh67_wm42_10_c5 :  std_logic;
signal bh67_wm41_10_c4, bh67_wm41_10_c5 :  std_logic;
signal bh67_wm40_10_c4, bh67_wm40_10_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid301_Out0_copy302_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid303_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid303_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm41_11_c5 :  std_logic;
signal bh67_wm40_11_c5 :  std_logic;
signal bh67_wm39_11_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid303_Out0_copy304_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid305_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid305_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh67_wm41_12_c4, bh67_wm41_12_c5 :  std_logic;
signal bh67_wm40_12_c4, bh67_wm40_12_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid305_Out0_copy306_c4 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid307_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid307_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm40_13_c5 :  std_logic;
signal bh67_wm39_12_c5 :  std_logic;
signal bh67_wm38_11_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid307_Out0_copy308_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid309_In0_c4, Compressor_14_3_Freq300_uid292_bh67_uid309_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid309_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid309_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm40_14_c5 :  std_logic;
signal bh67_wm39_13_c5 :  std_logic;
signal bh67_wm38_12_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid309_Out0_copy310_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid311_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid311_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm39_14_c4, bh67_wm39_14_c5 :  std_logic;
signal bh67_wm38_13_c4, bh67_wm38_13_c5 :  std_logic;
signal bh67_wm37_12_c4, bh67_wm37_12_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid311_Out0_copy312_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid313_In0_c4, Compressor_14_3_Freq300_uid292_bh67_uid313_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid313_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid313_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm39_15_c5 :  std_logic;
signal bh67_wm38_14_c5 :  std_logic;
signal bh67_wm37_13_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid313_Out0_copy314_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid315_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid315_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm38_15_c4, bh67_wm38_15_c5 :  std_logic;
signal bh67_wm37_14_c4, bh67_wm37_14_c5 :  std_logic;
signal bh67_wm36_10_c4, bh67_wm36_10_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid315_Out0_copy316_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid317_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid317_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh67_wm38_16_c4 :  std_logic;
signal bh67_wm37_15_c4, bh67_wm37_15_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid317_Out0_copy318_c4 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid319_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid319_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm37_16_c5 :  std_logic;
signal bh67_wm36_11_c5 :  std_logic;
signal bh67_wm35_10_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid319_Out0_copy320_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid321_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid321_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm37_17_c4, bh67_wm37_17_c5 :  std_logic;
signal bh67_wm36_12_c4, bh67_wm36_12_c5 :  std_logic;
signal bh67_wm35_11_c4, bh67_wm35_11_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid321_Out0_copy322_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid323_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid323_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm36_13_c5 :  std_logic;
signal bh67_wm35_12_c5 :  std_logic;
signal bh67_wm34_11_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid323_Out0_copy324_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid325_In0_c4, Compressor_14_3_Freq300_uid292_bh67_uid325_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid325_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid325_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm36_14_c5 :  std_logic;
signal bh67_wm35_13_c5 :  std_logic;
signal bh67_wm34_12_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid325_Out0_copy326_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid327_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid327_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm35_14_c4, bh67_wm35_14_c5 :  std_logic;
signal bh67_wm34_13_c4, bh67_wm34_13_c5 :  std_logic;
signal bh67_wm33_12_c4, bh67_wm33_12_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid327_Out0_copy328_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid329_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid329_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh67_wm35_15_c4, bh67_wm35_15_c5 :  std_logic;
signal bh67_wm34_14_c4, bh67_wm34_14_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid329_Out0_copy330_c4 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid331_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid331_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm34_15_c5 :  std_logic;
signal bh67_wm33_13_c5 :  std_logic;
signal bh67_wm32_10_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid331_Out0_copy332_c5 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid335_In0_c4 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid335_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm34_16_c4, bh67_wm34_16_c5 :  std_logic;
signal bh67_wm33_14_c4, bh67_wm33_14_c5 :  std_logic;
signal bh67_wm32_11_c4, bh67_wm32_11_c5 :  std_logic;
signal Compressor_5_3_Freq300_uid334_bh67_uid335_Out0_copy336_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid337_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid337_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm33_15_c5 :  std_logic;
signal bh67_wm32_12_c5 :  std_logic;
signal bh67_wm31_10_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid337_Out0_copy338_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid339_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid339_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm33_16_c4, bh67_wm33_16_c5 :  std_logic;
signal bh67_wm32_13_c4, bh67_wm32_13_c5 :  std_logic;
signal bh67_wm31_11_c4, bh67_wm31_11_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid339_Out0_copy340_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid341_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid341_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm32_14_c5 :  std_logic;
signal bh67_wm31_12_c5 :  std_logic;
signal bh67_wm30_11_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid341_Out0_copy342_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid343_In0_c4, Compressor_14_3_Freq300_uid292_bh67_uid343_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid343_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid343_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm32_15_c5 :  std_logic;
signal bh67_wm31_13_c5 :  std_logic;
signal bh67_wm30_12_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid343_Out0_copy344_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid345_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid345_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm31_14_c4, bh67_wm31_14_c5 :  std_logic;
signal bh67_wm30_13_c4, bh67_wm30_13_c5 :  std_logic;
signal bh67_wm29_12_c4, bh67_wm29_12_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid345_Out0_copy346_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid347_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid347_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh67_wm31_15_c4, bh67_wm31_15_c5 :  std_logic;
signal bh67_wm30_14_c4, bh67_wm30_14_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid347_Out0_copy348_c4 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid349_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid349_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm30_15_c5 :  std_logic;
signal bh67_wm29_13_c5 :  std_logic;
signal bh67_wm28_10_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid349_Out0_copy350_c5 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid351_In0_c4 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid351_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm30_16_c4, bh67_wm30_16_c5 :  std_logic;
signal bh67_wm29_14_c4, bh67_wm29_14_c5 :  std_logic;
signal bh67_wm28_11_c4, bh67_wm28_11_c5 :  std_logic;
signal Compressor_5_3_Freq300_uid334_bh67_uid351_Out0_copy352_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid353_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid353_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm29_15_c5 :  std_logic;
signal bh67_wm28_12_c5 :  std_logic;
signal bh67_wm27_10_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid353_Out0_copy354_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid355_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid355_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm29_16_c4, bh67_wm29_16_c5 :  std_logic;
signal bh67_wm28_13_c4, bh67_wm28_13_c5 :  std_logic;
signal bh67_wm27_11_c4, bh67_wm27_11_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid355_Out0_copy356_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid357_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid357_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm28_14_c5 :  std_logic;
signal bh67_wm27_12_c5 :  std_logic;
signal bh67_wm26_11_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid357_Out0_copy358_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid359_In0_c4, Compressor_14_3_Freq300_uid292_bh67_uid359_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid359_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid359_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm28_15_c5 :  std_logic;
signal bh67_wm27_13_c5 :  std_logic;
signal bh67_wm26_12_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid359_Out0_copy360_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid361_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid361_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm27_14_c4, bh67_wm27_14_c5 :  std_logic;
signal bh67_wm26_13_c4, bh67_wm26_13_c5 :  std_logic;
signal bh67_wm25_11_c4, bh67_wm25_11_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid361_Out0_copy362_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid363_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid363_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh67_wm27_15_c4, bh67_wm27_15_c5 :  std_logic;
signal bh67_wm26_14_c4, bh67_wm26_14_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid363_Out0_copy364_c4 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid365_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid365_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm26_15_c5 :  std_logic;
signal bh67_wm25_12_c5 :  std_logic;
signal bh67_wm24_8_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid365_Out0_copy366_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid367_In0_c4, Compressor_14_3_Freq300_uid292_bh67_uid367_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid367_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid367_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm26_16_c5 :  std_logic;
signal bh67_wm25_13_c5 :  std_logic;
signal bh67_wm24_9_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid367_Out0_copy368_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid369_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid369_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm25_14_c4, bh67_wm25_14_c5 :  std_logic;
signal bh67_wm24_10_c4, bh67_wm24_10_c5 :  std_logic;
signal bh67_wm23_8_c4 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid369_Out0_copy370_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid371_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid371_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid371_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm25_15_c4, bh67_wm25_15_c5 :  std_logic;
signal bh67_wm24_11_c4, bh67_wm24_11_c5 :  std_logic;
signal bh67_wm23_9_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid371_Out0_copy372_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid373_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid373_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm24_12_c4, bh67_wm24_12_c5 :  std_logic;
signal bh67_wm23_10_c4 :  std_logic;
signal bh67_wm22_8_c4 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid373_Out0_copy374_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid375_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid375_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm23_11_c4 :  std_logic;
signal bh67_wm22_9_c4 :  std_logic;
signal bh67_wm21_6_c4 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid375_Out0_copy376_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid377_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid377_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid377_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm23_12_c4, bh67_wm23_12_c5 :  std_logic;
signal bh67_wm22_10_c4 :  std_logic;
signal bh67_wm21_7_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid377_Out0_copy378_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid379_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid379_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm22_11_c4 :  std_logic;
signal bh67_wm21_8_c4 :  std_logic;
signal bh67_wm20_6_c4 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid379_Out0_copy380_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid381_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid381_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm21_9_c4 :  std_logic;
signal bh67_wm20_7_c4 :  std_logic;
signal bh67_wm19_5_c4 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid381_Out0_copy382_c4 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid383_In0_c4 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid383_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm20_8_c4 :  std_logic;
signal bh67_wm19_6_c4 :  std_logic;
signal bh67_wm18_4_c4 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid383_Out0_copy384_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid385_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid385_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid385_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm19_7_c4 :  std_logic;
signal bh67_wm18_5_c4 :  std_logic;
signal bh67_wm17_3_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid385_Out0_copy386_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid387_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid387_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid387_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm18_6_c4 :  std_logic;
signal bh67_wm17_4_c4 :  std_logic;
signal bh67_wm16_2_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid387_Out0_copy388_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid389_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid389_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid389_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm16_3_c4 :  std_logic;
signal bh67_wm15_2_c4 :  std_logic;
signal bh67_wm14_2_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid389_Out0_copy390_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid391_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid391_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid391_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm14_3_c4 :  std_logic;
signal bh67_wm13_2_c4 :  std_logic;
signal bh67_wm12_2_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid391_Out0_copy392_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid393_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid393_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid393_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm12_3_c4 :  std_logic;
signal bh67_wm11_2_c4 :  std_logic;
signal bh67_wm10_2_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid393_Out0_copy394_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid395_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid395_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid395_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm10_3_c4 :  std_logic;
signal bh67_wm9_2_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid395_Out0_copy396_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid397_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid397_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid397_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm46_5_c5 :  std_logic;
signal bh67_wm45_6_c5 :  std_logic;
signal bh67_wm44_7_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid397_Out0_copy398_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid399_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid399_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm44_8_c5 :  std_logic;
signal bh67_wm43_8_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid399_Out0_copy400_c5 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid401_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid401_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm43_9_c5 :  std_logic;
signal bh67_wm42_11_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid401_Out0_copy402_c5 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid403_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid403_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid403_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm42_12_c5 :  std_logic;
signal bh67_wm41_13_c5 :  std_logic;
signal bh67_wm40_15_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid403_Out0_copy404_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid405_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid405_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm41_14_c5 :  std_logic;
signal bh67_wm40_16_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid405_Out0_copy406_c5 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid407_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid407_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid407_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm40_17_c5 :  std_logic;
signal bh67_wm39_16_c5 :  std_logic;
signal bh67_wm38_17_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid407_Out0_copy408_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid409_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid409_In1_c4, Compressor_14_3_Freq300_uid292_bh67_uid409_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid409_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm39_17_c5 :  std_logic;
signal bh67_wm38_18_c5 :  std_logic;
signal bh67_wm37_18_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid409_Out0_copy410_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid411_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid411_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm38_19_c5 :  std_logic;
signal bh67_wm37_19_c5 :  std_logic;
signal bh67_wm36_15_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid411_Out0_copy412_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid413_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid413_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm37_20_c5 :  std_logic;
signal bh67_wm36_16_c5 :  std_logic;
signal bh67_wm35_16_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid413_Out0_copy414_c5 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid415_In0_c5 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid415_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm36_17_c5 :  std_logic;
signal bh67_wm35_17_c5 :  std_logic;
signal bh67_wm34_17_c5 :  std_logic;
signal Compressor_5_3_Freq300_uid334_bh67_uid415_Out0_copy416_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid417_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid417_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm35_18_c5 :  std_logic;
signal bh67_wm34_18_c5 :  std_logic;
signal bh67_wm33_17_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid417_Out0_copy418_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid419_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid419_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm34_19_c5 :  std_logic;
signal bh67_wm33_18_c5 :  std_logic;
signal bh67_wm32_16_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid419_Out0_copy420_c5 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid421_In0_c5 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid421_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm33_19_c5 :  std_logic;
signal bh67_wm32_17_c5 :  std_logic;
signal bh67_wm31_16_c5 :  std_logic;
signal Compressor_5_3_Freq300_uid334_bh67_uid421_Out0_copy422_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid423_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid423_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm32_18_c5 :  std_logic;
signal bh67_wm31_17_c5 :  std_logic;
signal bh67_wm30_17_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid423_Out0_copy424_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid425_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid425_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm31_18_c5 :  std_logic;
signal bh67_wm30_18_c5 :  std_logic;
signal bh67_wm29_17_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid425_Out0_copy426_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid427_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid427_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm30_19_c5 :  std_logic;
signal bh67_wm29_18_c5 :  std_logic;
signal bh67_wm28_16_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid427_Out0_copy428_c5 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid429_In0_c5 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid429_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm29_19_c5 :  std_logic;
signal bh67_wm28_17_c5 :  std_logic;
signal bh67_wm27_16_c5 :  std_logic;
signal Compressor_5_3_Freq300_uid334_bh67_uid429_Out0_copy430_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid431_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid431_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm28_18_c5 :  std_logic;
signal bh67_wm27_17_c5 :  std_logic;
signal bh67_wm26_17_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid431_Out0_copy432_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid433_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid433_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm27_18_c5 :  std_logic;
signal bh67_wm26_18_c5 :  std_logic;
signal bh67_wm25_16_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid433_Out0_copy434_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid435_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid435_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm26_19_c5 :  std_logic;
signal bh67_wm25_17_c5 :  std_logic;
signal bh67_wm24_13_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid435_Out0_copy436_c5 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid437_In0_c5 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid334_bh67_uid437_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm25_18_c5 :  std_logic;
signal bh67_wm24_14_c5 :  std_logic;
signal bh67_wm23_13_c5 :  std_logic;
signal Compressor_5_3_Freq300_uid334_bh67_uid437_Out0_copy438_c5 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid439_In0_c5 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid300_bh67_uid439_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm24_15_c5 :  std_logic;
signal bh67_wm23_14_c5 :  std_logic;
signal bh67_wm22_12_c5 :  std_logic;
signal Compressor_6_3_Freq300_uid300_bh67_uid439_Out0_copy440_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid441_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid441_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid441_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm23_15_c4, bh67_wm23_15_c5 :  std_logic;
signal bh67_wm22_13_c4, bh67_wm22_13_c5 :  std_logic;
signal bh67_wm21_10_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid441_Out0_copy442_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid443_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid443_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh67_wm22_14_c4, bh67_wm22_14_c5 :  std_logic;
signal bh67_wm21_11_c4 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid443_Out0_copy444_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid445_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid445_In1_c0, Compressor_14_3_Freq300_uid292_bh67_uid445_In1_c1, Compressor_14_3_Freq300_uid292_bh67_uid445_In1_c2, Compressor_14_3_Freq300_uid292_bh67_uid445_In1_c3, Compressor_14_3_Freq300_uid292_bh67_uid445_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid445_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm21_12_c4 :  std_logic;
signal bh67_wm20_9_c4 :  std_logic;
signal bh67_wm19_8_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid445_Out0_copy446_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid447_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid447_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh67_wm20_10_c4 :  std_logic;
signal bh67_wm19_9_c4 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid447_Out0_copy448_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid449_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid449_In1_c0, Compressor_14_3_Freq300_uid292_bh67_uid449_In1_c1, Compressor_14_3_Freq300_uid292_bh67_uid449_In1_c2, Compressor_14_3_Freq300_uid292_bh67_uid449_In1_c3, Compressor_14_3_Freq300_uid292_bh67_uid449_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid449_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm19_10_c4 :  std_logic;
signal bh67_wm18_7_c4 :  std_logic;
signal bh67_wm17_5_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid449_Out0_copy450_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid451_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid451_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh67_wm18_8_c4 :  std_logic;
signal bh67_wm17_6_c4 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid451_Out0_copy452_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid453_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid453_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid453_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm17_7_c4 :  std_logic;
signal bh67_wm16_4_c4, bh67_wm16_4_c5 :  std_logic;
signal bh67_wm15_3_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid453_Out0_copy454_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid455_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid455_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid455_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm14_4_c4 :  std_logic;
signal bh67_wm13_3_c4 :  std_logic;
signal bh67_wm12_4_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid455_Out0_copy456_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid457_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid457_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid457_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm12_5_c4 :  std_logic;
signal bh67_wm11_3_c4 :  std_logic;
signal bh67_wm10_4_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid457_Out0_copy458_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid459_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid459_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid459_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm10_5_c4 :  std_logic;
signal bh67_wm9_3_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid459_Out0_copy460_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid461_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid461_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid461_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm44_9_c5 :  std_logic;
signal bh67_wm43_10_c5 :  std_logic;
signal bh67_wm42_13_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid461_Out0_copy462_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid463_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid463_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid463_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm42_14_c5 :  std_logic;
signal bh67_wm41_15_c5 :  std_logic;
signal bh67_wm40_18_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid463_Out0_copy464_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid465_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid465_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid465_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm40_19_c5 :  std_logic;
signal bh67_wm39_18_c5 :  std_logic;
signal bh67_wm38_20_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid465_Out0_copy466_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid467_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid467_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid467_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm38_21_c5 :  std_logic;
signal bh67_wm37_21_c5 :  std_logic;
signal bh67_wm36_18_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid467_Out0_copy468_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid469_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid469_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid469_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm36_19_c5 :  std_logic;
signal bh67_wm35_19_c5 :  std_logic;
signal bh67_wm34_20_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid469_Out0_copy470_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid471_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid471_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid471_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm34_21_c5 :  std_logic;
signal bh67_wm33_20_c5 :  std_logic;
signal bh67_wm32_19_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid471_Out0_copy472_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid473_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid473_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid473_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm32_20_c5 :  std_logic;
signal bh67_wm31_19_c5 :  std_logic;
signal bh67_wm30_20_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid473_Out0_copy474_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid475_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid475_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid475_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm30_21_c5 :  std_logic;
signal bh67_wm29_20_c5 :  std_logic;
signal bh67_wm28_19_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid475_Out0_copy476_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid477_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid477_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid477_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm28_20_c5 :  std_logic;
signal bh67_wm27_19_c5 :  std_logic;
signal bh67_wm26_20_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid477_Out0_copy478_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid479_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c0, Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c1, Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c2, Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c3, Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c4, Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid479_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm26_21_c5 :  std_logic;
signal bh67_wm25_19_c5 :  std_logic;
signal bh67_wm24_16_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid479_Out0_copy480_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid481_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid481_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm25_20_c5 :  std_logic;
signal bh67_wm24_17_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid481_Out0_copy482_c5 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid483_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid483_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm24_18_c5 :  std_logic;
signal bh67_wm23_16_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid483_Out0_copy484_c5 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid485_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c0, Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c1, Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c2, Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c3, Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c4, Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid485_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm23_17_c5 :  std_logic;
signal bh67_wm22_15_c5 :  std_logic;
signal bh67_wm21_13_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid485_Out0_copy486_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid487_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid487_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm22_16_c5 :  std_logic;
signal bh67_wm21_14_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid487_Out0_copy488_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid489_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid489_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm21_15_c5 :  std_logic;
signal bh67_wm20_11_c5 :  std_logic;
signal bh67_wm19_11_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_copy490_c4, Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_copy490_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid491_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid491_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm19_12_c5 :  std_logic;
signal bh67_wm18_9_c5 :  std_logic;
signal bh67_wm17_8_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_copy492_c4, Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_copy492_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid493_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm17_9_c5 :  std_logic;
signal bh67_wm16_5_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_copy494_c4, Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_copy494_c5 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid495_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid495_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid495_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm15_4_c4, bh67_wm15_4_c5 :  std_logic;
signal bh67_wm14_5_c4, bh67_wm14_5_c5 :  std_logic;
signal bh67_wm13_4_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid495_Out0_copy496_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid497_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid497_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid497_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm12_6_c4 :  std_logic;
signal bh67_wm11_4_c4, bh67_wm11_4_c5 :  std_logic;
signal bh67_wm10_6_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid497_Out0_copy498_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid499_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid499_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid499_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh67_wm10_7_c4 :  std_logic;
signal bh67_wm9_4_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid499_Out0_copy500_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid501_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid501_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid501_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm42_15_c5 :  std_logic;
signal bh67_wm41_16_c5 :  std_logic;
signal bh67_wm40_20_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid501_Out0_copy502_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid503_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid503_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid503_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm40_21_c5 :  std_logic;
signal bh67_wm39_19_c5 :  std_logic;
signal bh67_wm38_22_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid503_Out0_copy504_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid505_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid505_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid505_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm38_23_c5 :  std_logic;
signal bh67_wm37_22_c5 :  std_logic;
signal bh67_wm36_20_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid505_Out0_copy506_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid507_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid507_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid507_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm36_21_c5 :  std_logic;
signal bh67_wm35_20_c5 :  std_logic;
signal bh67_wm34_22_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid507_Out0_copy508_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid509_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid509_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid509_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm34_23_c5 :  std_logic;
signal bh67_wm33_21_c5 :  std_logic;
signal bh67_wm32_21_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid509_Out0_copy510_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid511_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid511_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid511_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm32_22_c5 :  std_logic;
signal bh67_wm31_20_c5 :  std_logic;
signal bh67_wm30_22_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid511_Out0_copy512_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid513_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid513_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid513_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm30_23_c5 :  std_logic;
signal bh67_wm29_21_c5 :  std_logic;
signal bh67_wm28_21_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid513_Out0_copy514_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid515_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid515_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid515_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm28_22_c5 :  std_logic;
signal bh67_wm27_20_c5 :  std_logic;
signal bh67_wm26_22_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid515_Out0_copy516_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid517_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid517_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid517_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm26_23_c5 :  std_logic;
signal bh67_wm25_21_c5 :  std_logic;
signal bh67_wm24_19_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid517_Out0_copy518_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid519_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid519_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid519_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm24_20_c5 :  std_logic;
signal bh67_wm23_18_c5 :  std_logic;
signal bh67_wm22_17_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid519_Out0_copy520_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid521_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid521_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm22_18_c5 :  std_logic;
signal bh67_wm21_16_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid521_Out0_copy522_c5 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid523_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid288_bh67_uid523_Out0_c5 :  std_logic_vector(1 downto 0);
signal bh67_wm21_17_c5 :  std_logic;
signal bh67_wm20_12_c5 :  std_logic;
signal Compressor_3_2_Freq300_uid288_bh67_uid523_Out0_copy524_c5 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid525_In0_c5 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid525_In1_c5 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid525_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm19_13_c5 :  std_logic;
signal bh67_wm18_10_c5 :  std_logic;
signal bh67_wm17_10_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid525_Out0_copy526_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid527_In0_c5 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid527_In1_c5 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid284_bh67_uid527_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm17_11_c5 :  std_logic;
signal bh67_wm16_6_c5 :  std_logic;
signal bh67_wm15_5_c5 :  std_logic;
signal Compressor_23_3_Freq300_uid284_bh67_uid527_Out0_copy528_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid529_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid529_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm13_5_c5 :  std_logic;
signal bh67_wm12_7_c5 :  std_logic;
signal bh67_wm11_5_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_copy530_c4, Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_copy530_c5 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid531_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid531_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_c5 :  std_logic_vector(2 downto 0);
signal bh67_wm10_8_c5 :  std_logic;
signal bh67_wm9_5_c5 :  std_logic;
signal Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_copy532_c4, Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_copy532_c5 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh67_24_c5, tmp_bitheapResult_bh67_24_c6 :  std_logic_vector(24 downto 0);
signal bitheapFinalAdd_bh67_In0_c5 :  std_logic_vector(32 downto 0);
signal bitheapFinalAdd_bh67_In1_c5 :  std_logic_vector(32 downto 0);
signal bitheapFinalAdd_bh67_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh67_Out_c6 :  std_logic_vector(32 downto 0);
signal bitheapResult_bh67_c6 :  std_logic_vector(56 downto 0);
signal RR_c6 :  signed(-9+41 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               bh67_wm26_1_c5 <= bh67_wm26_1_c4;
               bh67_wm28_1_c5 <= bh67_wm28_1_c4;
               bh67_wm26_2_c5 <= bh67_wm26_2_c4;
               bh67_wm26_3_c5 <= bh67_wm26_3_c4;
               bh67_wm30_1_c5 <= bh67_wm30_1_c4;
               bh67_wm29_1_c5 <= bh67_wm29_1_c4;
               bh67_wm28_2_c5 <= bh67_wm28_2_c4;
               bh67_wm26_4_c5 <= bh67_wm26_4_c4;
               bh67_wm26_5_c5 <= bh67_wm26_5_c4;
               bh67_wm29_2_c5 <= bh67_wm29_2_c4;
               bh67_wm28_3_c5 <= bh67_wm28_3_c4;
               bh67_wm32_1_c5 <= bh67_wm32_1_c4;
               bh67_wm30_2_c5 <= bh67_wm30_2_c4;
               bh67_wm29_3_c5 <= bh67_wm29_3_c4;
               bh67_wm28_4_c5 <= bh67_wm28_4_c4;
               bh67_wm28_5_c5 <= bh67_wm28_5_c4;
               bh67_wm30_3_c5 <= bh67_wm30_3_c4;
               bh67_wm29_4_c5 <= bh67_wm29_4_c4;
               bh67_wm34_1_c5 <= bh67_wm34_1_c4;
               bh67_wm33_1_c5 <= bh67_wm33_1_c4;
               bh67_wm32_2_c5 <= bh67_wm32_2_c4;
               bh67_wm30_4_c5 <= bh67_wm30_4_c4;
               bh67_wm30_5_c5 <= bh67_wm30_5_c4;
               bh67_wm29_5_c5 <= bh67_wm29_5_c4;
               bh67_wm33_2_c5 <= bh67_wm33_2_c4;
               bh67_wm32_3_c5 <= bh67_wm32_3_c4;
               bh67_wm36_1_c5 <= bh67_wm36_1_c4;
               bh67_wm34_2_c5 <= bh67_wm34_2_c4;
               bh67_wm33_3_c5 <= bh67_wm33_3_c4;
               bh67_wm32_4_c5 <= bh67_wm32_4_c4;
               bh67_wm32_5_c5 <= bh67_wm32_5_c4;
               bh67_wm34_3_c5 <= bh67_wm34_3_c4;
               bh67_wm33_4_c5 <= bh67_wm33_4_c4;
               bh67_wm37_1_c5 <= bh67_wm37_1_c4;
               bh67_wm36_2_c5 <= bh67_wm36_2_c4;
               bh67_wm34_4_c5 <= bh67_wm34_4_c4;
               bh67_wm34_5_c5 <= bh67_wm34_5_c4;
               bh67_wm33_5_c5 <= bh67_wm33_5_c4;
               bh67_wm37_2_c5 <= bh67_wm37_2_c4;
               bh67_wm36_3_c5 <= bh67_wm36_3_c4;
               bh67_wm40_1_c5 <= bh67_wm40_1_c4;
               bh67_wm37_3_c5 <= bh67_wm37_3_c4;
               bh67_wm36_4_c5 <= bh67_wm36_4_c4;
               bh67_wm36_5_c5 <= bh67_wm36_5_c4;
               bh67_wm37_4_c5 <= bh67_wm37_4_c4;
               bh67_wm41_1_c5 <= bh67_wm41_1_c4;
               bh67_wm40_2_c5 <= bh67_wm40_2_c4;
               bh67_wm37_5_c5 <= bh67_wm37_5_c4;
               bh67_wm41_2_c5 <= bh67_wm41_2_c4;
               bh67_wm40_3_c5 <= bh67_wm40_3_c4;
               bh67_wm41_3_c5 <= bh67_wm41_3_c4;
               bh67_wm40_4_c5 <= bh67_wm40_4_c4;
               bh67_wm40_5_c5 <= bh67_wm40_5_c4;
               bh67_wm41_4_c5 <= bh67_wm41_4_c4;
               bh67_wm46_1_c5 <= bh67_wm46_1_c4;
               bh67_wm45_1_c5 <= bh67_wm45_1_c4;
               bh67_wm41_5_c5 <= bh67_wm41_5_c4;
               bh67_wm45_2_c5 <= bh67_wm45_2_c4;
               bh67_wm48_1_c5 <= bh67_wm48_1_c4;
               bh67_wm47_1_c5 <= bh67_wm47_1_c4;
               bh67_wm46_2_c5 <= bh67_wm46_2_c4;
               bh67_wm45_3_c5 <= bh67_wm45_3_c4;
               bh67_wm24_7_c5 <= bh67_wm24_7_c4;
               bh67_wm42_7_c5 <= bh67_wm42_7_c4;
               bh67_wm38_10_c5 <= bh67_wm38_10_c4;
               bh67_wm26_10_c5 <= bh67_wm26_10_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid295_In0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid295_In0_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid297_In0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid297_In0_c4;
               bh67_wm42_10_c5 <= bh67_wm42_10_c4;
               bh67_wm41_10_c5 <= bh67_wm41_10_c4;
               bh67_wm40_10_c5 <= bh67_wm40_10_c4;
               bh67_wm41_12_c5 <= bh67_wm41_12_c4;
               bh67_wm40_12_c5 <= bh67_wm40_12_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid309_In0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid309_In0_c4;
               bh67_wm39_14_c5 <= bh67_wm39_14_c4;
               bh67_wm38_13_c5 <= bh67_wm38_13_c4;
               bh67_wm37_12_c5 <= bh67_wm37_12_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid313_In0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid313_In0_c4;
               bh67_wm38_15_c5 <= bh67_wm38_15_c4;
               bh67_wm37_14_c5 <= bh67_wm37_14_c4;
               bh67_wm36_10_c5 <= bh67_wm36_10_c4;
               bh67_wm37_15_c5 <= bh67_wm37_15_c4;
               bh67_wm37_17_c5 <= bh67_wm37_17_c4;
               bh67_wm36_12_c5 <= bh67_wm36_12_c4;
               bh67_wm35_11_c5 <= bh67_wm35_11_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid325_In0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid325_In0_c4;
               bh67_wm35_14_c5 <= bh67_wm35_14_c4;
               bh67_wm34_13_c5 <= bh67_wm34_13_c4;
               bh67_wm33_12_c5 <= bh67_wm33_12_c4;
               bh67_wm35_15_c5 <= bh67_wm35_15_c4;
               bh67_wm34_14_c5 <= bh67_wm34_14_c4;
               bh67_wm34_16_c5 <= bh67_wm34_16_c4;
               bh67_wm33_14_c5 <= bh67_wm33_14_c4;
               bh67_wm32_11_c5 <= bh67_wm32_11_c4;
               bh67_wm33_16_c5 <= bh67_wm33_16_c4;
               bh67_wm32_13_c5 <= bh67_wm32_13_c4;
               bh67_wm31_11_c5 <= bh67_wm31_11_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid343_In0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid343_In0_c4;
               bh67_wm31_14_c5 <= bh67_wm31_14_c4;
               bh67_wm30_13_c5 <= bh67_wm30_13_c4;
               bh67_wm29_12_c5 <= bh67_wm29_12_c4;
               bh67_wm31_15_c5 <= bh67_wm31_15_c4;
               bh67_wm30_14_c5 <= bh67_wm30_14_c4;
               bh67_wm30_16_c5 <= bh67_wm30_16_c4;
               bh67_wm29_14_c5 <= bh67_wm29_14_c4;
               bh67_wm28_11_c5 <= bh67_wm28_11_c4;
               bh67_wm29_16_c5 <= bh67_wm29_16_c4;
               bh67_wm28_13_c5 <= bh67_wm28_13_c4;
               bh67_wm27_11_c5 <= bh67_wm27_11_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid359_In0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid359_In0_c4;
               bh67_wm27_14_c5 <= bh67_wm27_14_c4;
               bh67_wm26_13_c5 <= bh67_wm26_13_c4;
               bh67_wm25_11_c5 <= bh67_wm25_11_c4;
               bh67_wm27_15_c5 <= bh67_wm27_15_c4;
               bh67_wm26_14_c5 <= bh67_wm26_14_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid367_In0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid367_In0_c4;
               bh67_wm25_14_c5 <= bh67_wm25_14_c4;
               bh67_wm24_10_c5 <= bh67_wm24_10_c4;
               bh67_wm25_15_c5 <= bh67_wm25_15_c4;
               bh67_wm24_11_c5 <= bh67_wm24_11_c4;
               bh67_wm24_12_c5 <= bh67_wm24_12_c4;
               bh67_wm23_12_c5 <= bh67_wm23_12_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid409_In1_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid409_In1_c4;
               bh67_wm23_15_c5 <= bh67_wm23_15_c4;
               bh67_wm22_13_c5 <= bh67_wm22_13_c4;
               bh67_wm22_14_c5 <= bh67_wm22_14_c4;
               bh67_wm16_4_c5 <= bh67_wm16_4_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c4;
               Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_copy490_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_copy490_c4;
               Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_copy492_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_copy492_c4;
               Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_copy494_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_copy494_c4;
               bh67_wm15_4_c5 <= bh67_wm15_4_c4;
               bh67_wm14_5_c5 <= bh67_wm14_5_c4;
               bh67_wm11_4_c5 <= bh67_wm11_4_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_copy530_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_copy530_c4;
               Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_copy532_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_copy532_c4;
            end if;
            if ce_6 = '1' then
               tmp_bitheapResult_bh67_24_c6 <= tmp_bitheapResult_bh67_24_c5;
            end if;
         end if;
      end process;
XX_c4 <= signed(X);
YY_c4 <= signed(Y);
AA_c4 <= signed(A);
   tile_0_X_c4 <= X(16 downto 0);
   tile_0_Y_c4 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid69
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 X => tile_0_X_c4,
                 Y => tile_0_Y_c4,
                 R => tile_0_output_c5);

   tile_0_filtered_output_c5 <= unsigned(tile_0_output_c5(40 downto 0));
   bh67_wm65_0_c5 <= tile_0_filtered_output_c5(0);
   bh67_wm64_0_c5 <= tile_0_filtered_output_c5(1);
   bh67_wm63_0_c5 <= tile_0_filtered_output_c5(2);
   bh67_wm62_0_c5 <= tile_0_filtered_output_c5(3);
   bh67_wm61_0_c5 <= tile_0_filtered_output_c5(4);
   bh67_wm60_0_c5 <= tile_0_filtered_output_c5(5);
   bh67_wm59_0_c5 <= tile_0_filtered_output_c5(6);
   bh67_wm58_0_c5 <= tile_0_filtered_output_c5(7);
   bh67_wm57_0_c5 <= tile_0_filtered_output_c5(8);
   bh67_wm56_0_c5 <= tile_0_filtered_output_c5(9);
   bh67_wm55_0_c5 <= tile_0_filtered_output_c5(10);
   bh67_wm54_0_c5 <= tile_0_filtered_output_c5(11);
   bh67_wm53_0_c5 <= tile_0_filtered_output_c5(12);
   bh67_wm52_0_c5 <= tile_0_filtered_output_c5(13);
   bh67_wm51_0_c5 <= tile_0_filtered_output_c5(14);
   bh67_wm50_0_c5 <= tile_0_filtered_output_c5(15);
   bh67_wm49_0_c5 <= tile_0_filtered_output_c5(16);
   bh67_wm48_0_c5 <= tile_0_filtered_output_c5(17);
   bh67_wm47_0_c5 <= tile_0_filtered_output_c5(18);
   bh67_wm46_0_c5 <= tile_0_filtered_output_c5(19);
   bh67_wm45_0_c5 <= tile_0_filtered_output_c5(20);
   bh67_wm44_0_c5 <= tile_0_filtered_output_c5(21);
   bh67_wm43_0_c5 <= tile_0_filtered_output_c5(22);
   bh67_wm42_0_c5 <= tile_0_filtered_output_c5(23);
   bh67_wm41_0_c5 <= tile_0_filtered_output_c5(24);
   bh67_wm40_0_c5 <= tile_0_filtered_output_c5(25);
   bh67_wm39_0_c5 <= tile_0_filtered_output_c5(26);
   bh67_wm38_0_c5 <= tile_0_filtered_output_c5(27);
   bh67_wm37_0_c5 <= tile_0_filtered_output_c5(28);
   bh67_wm36_0_c5 <= tile_0_filtered_output_c5(29);
   bh67_wm35_0_c5 <= tile_0_filtered_output_c5(30);
   bh67_wm34_0_c5 <= tile_0_filtered_output_c5(31);
   bh67_wm33_0_c5 <= tile_0_filtered_output_c5(32);
   bh67_wm32_0_c5 <= tile_0_filtered_output_c5(33);
   bh67_wm31_0_c5 <= tile_0_filtered_output_c5(34);
   bh67_wm30_0_c5 <= tile_0_filtered_output_c5(35);
   bh67_wm29_0_c5 <= tile_0_filtered_output_c5(36);
   bh67_wm28_0_c5 <= tile_0_filtered_output_c5(37);
   bh67_wm27_0_c5 <= tile_0_filtered_output_c5(38);
   bh67_wm26_0_c5 <= tile_0_filtered_output_c5(39);
   bh67_wm25_0_c5 <= tile_0_filtered_output_c5(40);
   tile_1_X_c4 <= X(24 downto 23);
   tile_1_Y_c4 <= Y(23 downto 22);
   tile_1_mult: IntMultiplierLUT_2_signedx2_Freq300_uid71
      port map ( clk  => clk,
                 X => tile_1_X_c4,
                 Y => tile_1_Y_c4,
                 R => tile_1_output_c4);

   tile_1_filtered_output_c4 <= signed(tile_1_output_c4(3 downto 0));
   bh67_wm20_0_c4 <= tile_1_filtered_output_c4(0);
   bh67_wm19_0_c4 <= tile_1_filtered_output_c4(1);
   bh67_wm18_0_c4 <= tile_1_filtered_output_c4(2);
   bh67_wm17_0_c4 <= not tile_1_filtered_output_c4(3);
   tile_2_X_c4 <= X(22 downto 20);
   tile_2_Y_c4 <= Y(23 downto 22);
   tile_2_mult: IntMultiplierLUT_3x2_Freq300_uid76
      port map ( clk  => clk,
                 X => tile_2_X_c4,
                 Y => tile_2_Y_c4,
                 R => tile_2_output_c4);

   tile_2_filtered_output_c4 <= unsigned(tile_2_output_c4(4 downto 0));
   bh67_wm23_0_c4 <= tile_2_filtered_output_c4(0);
   bh67_wm22_0_c4 <= tile_2_filtered_output_c4(1);
   bh67_wm21_0_c4 <= tile_2_filtered_output_c4(2);
   bh67_wm20_1_c4 <= tile_2_filtered_output_c4(3);
   bh67_wm19_1_c4 <= tile_2_filtered_output_c4(4);
   tile_3_X_c4 <= X(19 downto 17);
   tile_3_Y_c4 <= Y(23 downto 22);
   tile_3_mult: IntMultiplierLUT_3x2_Freq300_uid81
      port map ( clk  => clk,
                 X => tile_3_X_c4,
                 Y => tile_3_Y_c4,
                 R => tile_3_output_c4);

   tile_3_filtered_output_c4 <= unsigned(tile_3_output_c4(4 downto 0));
   bh67_wm26_1_c4 <= tile_3_filtered_output_c4(0);
   bh67_wm25_1_c4 <= tile_3_filtered_output_c4(1);
   bh67_wm24_0_c4 <= tile_3_filtered_output_c4(2);
   bh67_wm23_1_c4 <= tile_3_filtered_output_c4(3);
   bh67_wm22_1_c4 <= tile_3_filtered_output_c4(4);
   tile_4_X_c4 <= X(24 downto 23);
   tile_4_Y_c4 <= Y(21 downto 20);
   tile_4_mult: IntMultiplierLUT_2_signedx2_Freq300_uid86
      port map ( clk  => clk,
                 X => tile_4_X_c4,
                 Y => tile_4_Y_c4,
                 R => tile_4_output_c4);

   tile_4_filtered_output_c4 <= signed(tile_4_output_c4(3 downto 0));
   bh67_wm22_2_c4 <= tile_4_filtered_output_c4(0);
   bh67_wm21_1_c4 <= tile_4_filtered_output_c4(1);
   bh67_wm20_2_c4 <= tile_4_filtered_output_c4(2);
   bh67_wm19_2_c4 <= not tile_4_filtered_output_c4(3);
   tile_5_X_c4 <= X(22 downto 20);
   tile_5_Y_c4 <= Y(21 downto 20);
   tile_5_mult: IntMultiplierLUT_3x2_Freq300_uid91
      port map ( clk  => clk,
                 X => tile_5_X_c4,
                 Y => tile_5_Y_c4,
                 R => tile_5_output_c4);

   tile_5_filtered_output_c4 <= unsigned(tile_5_output_c4(4 downto 0));
   bh67_wm25_2_c4 <= tile_5_filtered_output_c4(0);
   bh67_wm24_1_c4 <= tile_5_filtered_output_c4(1);
   bh67_wm23_2_c4 <= tile_5_filtered_output_c4(2);
   bh67_wm22_3_c4 <= tile_5_filtered_output_c4(3);
   bh67_wm21_2_c4 <= tile_5_filtered_output_c4(4);
   tile_6_X_c4 <= X(19 downto 17);
   tile_6_Y_c4 <= Y(21 downto 20);
   tile_6_mult: IntMultiplierLUT_3x2_Freq300_uid96
      port map ( clk  => clk,
                 X => tile_6_X_c4,
                 Y => tile_6_Y_c4,
                 R => tile_6_output_c4);

   tile_6_filtered_output_c4 <= unsigned(tile_6_output_c4(4 downto 0));
   bh67_wm28_1_c4 <= tile_6_filtered_output_c4(0);
   bh67_wm27_1_c4 <= tile_6_filtered_output_c4(1);
   bh67_wm26_2_c4 <= tile_6_filtered_output_c4(2);
   bh67_wm25_3_c4 <= tile_6_filtered_output_c4(3);
   bh67_wm24_2_c4 <= tile_6_filtered_output_c4(4);
   tile_7_X_c4 <= X(24 downto 23);
   tile_7_Y_c4 <= Y(19 downto 18);
   tile_7_mult: IntMultiplierLUT_2_signedx2_Freq300_uid101
      port map ( clk  => clk,
                 X => tile_7_X_c4,
                 Y => tile_7_Y_c4,
                 R => tile_7_output_c4);

   tile_7_filtered_output_c4 <= signed(tile_7_output_c4(3 downto 0));
   bh67_wm24_3_c4 <= tile_7_filtered_output_c4(0);
   bh67_wm23_3_c4 <= tile_7_filtered_output_c4(1);
   bh67_wm22_4_c4 <= tile_7_filtered_output_c4(2);
   bh67_wm21_3_c4 <= not tile_7_filtered_output_c4(3);
   tile_8_X_c4 <= X(22 downto 20);
   tile_8_Y_c4 <= Y(19 downto 18);
   tile_8_mult: IntMultiplierLUT_3x2_Freq300_uid106
      port map ( clk  => clk,
                 X => tile_8_X_c4,
                 Y => tile_8_Y_c4,
                 R => tile_8_output_c4);

   tile_8_filtered_output_c4 <= unsigned(tile_8_output_c4(4 downto 0));
   bh67_wm27_2_c4 <= tile_8_filtered_output_c4(0);
   bh67_wm26_3_c4 <= tile_8_filtered_output_c4(1);
   bh67_wm25_4_c4 <= tile_8_filtered_output_c4(2);
   bh67_wm24_4_c4 <= tile_8_filtered_output_c4(3);
   bh67_wm23_4_c4 <= tile_8_filtered_output_c4(4);
   tile_9_X_c4 <= X(19 downto 17);
   tile_9_Y_c4 <= Y(19 downto 18);
   tile_9_mult: IntMultiplierLUT_3x2_Freq300_uid111
      port map ( clk  => clk,
                 X => tile_9_X_c4,
                 Y => tile_9_Y_c4,
                 R => tile_9_output_c4);

   tile_9_filtered_output_c4 <= unsigned(tile_9_output_c4(4 downto 0));
   bh67_wm30_1_c4 <= tile_9_filtered_output_c4(0);
   bh67_wm29_1_c4 <= tile_9_filtered_output_c4(1);
   bh67_wm28_2_c4 <= tile_9_filtered_output_c4(2);
   bh67_wm27_3_c4 <= tile_9_filtered_output_c4(3);
   bh67_wm26_4_c4 <= tile_9_filtered_output_c4(4);
   tile_10_X_c4 <= X(24 downto 23);
   tile_10_Y_c4 <= Y(17 downto 16);
   tile_10_mult: IntMultiplierLUT_2_signedx2_Freq300_uid116
      port map ( clk  => clk,
                 X => tile_10_X_c4,
                 Y => tile_10_Y_c4,
                 R => tile_10_output_c4);

   tile_10_filtered_output_c4 <= signed(tile_10_output_c4(3 downto 0));
   bh67_wm26_5_c4 <= tile_10_filtered_output_c4(0);
   bh67_wm25_5_c4 <= tile_10_filtered_output_c4(1);
   bh67_wm24_5_c4 <= tile_10_filtered_output_c4(2);
   bh67_wm23_5_c4 <= not tile_10_filtered_output_c4(3);
   tile_11_X_c4 <= X(22 downto 20);
   tile_11_Y_c4 <= Y(17 downto 16);
   tile_11_mult: IntMultiplierLUT_3x2_Freq300_uid121
      port map ( clk  => clk,
                 X => tile_11_X_c4,
                 Y => tile_11_Y_c4,
                 R => tile_11_output_c4);

   tile_11_filtered_output_c4 <= unsigned(tile_11_output_c4(4 downto 0));
   bh67_wm29_2_c4 <= tile_11_filtered_output_c4(0);
   bh67_wm28_3_c4 <= tile_11_filtered_output_c4(1);
   bh67_wm27_4_c4 <= tile_11_filtered_output_c4(2);
   bh67_wm26_6_c4 <= tile_11_filtered_output_c4(3);
   bh67_wm25_6_c4 <= tile_11_filtered_output_c4(4);
   tile_12_X_c4 <= X(19 downto 17);
   tile_12_Y_c4 <= Y(17 downto 16);
   tile_12_mult: IntMultiplierLUT_3x2_Freq300_uid126
      port map ( clk  => clk,
                 X => tile_12_X_c4,
                 Y => tile_12_Y_c4,
                 R => tile_12_output_c4);

   tile_12_filtered_output_c4 <= unsigned(tile_12_output_c4(4 downto 0));
   bh67_wm32_1_c4 <= tile_12_filtered_output_c4(0);
   bh67_wm31_1_c4 <= tile_12_filtered_output_c4(1);
   bh67_wm30_2_c4 <= tile_12_filtered_output_c4(2);
   bh67_wm29_3_c4 <= tile_12_filtered_output_c4(3);
   bh67_wm28_4_c4 <= tile_12_filtered_output_c4(4);
   tile_13_X_c4 <= X(24 downto 23);
   tile_13_Y_c4 <= Y(15 downto 14);
   tile_13_mult: IntMultiplierLUT_2_signedx2_Freq300_uid131
      port map ( clk  => clk,
                 X => tile_13_X_c4,
                 Y => tile_13_Y_c4,
                 R => tile_13_output_c4);

   tile_13_filtered_output_c4 <= signed(tile_13_output_c4(3 downto 0));
   bh67_wm28_5_c4 <= tile_13_filtered_output_c4(0);
   bh67_wm27_5_c4 <= tile_13_filtered_output_c4(1);
   bh67_wm26_7_c4 <= tile_13_filtered_output_c4(2);
   bh67_wm25_7_c4 <= not tile_13_filtered_output_c4(3);
   tile_14_X_c4 <= X(22 downto 20);
   tile_14_Y_c4 <= Y(15 downto 14);
   tile_14_mult: IntMultiplierLUT_3x2_Freq300_uid136
      port map ( clk  => clk,
                 X => tile_14_X_c4,
                 Y => tile_14_Y_c4,
                 R => tile_14_output_c4);

   tile_14_filtered_output_c4 <= unsigned(tile_14_output_c4(4 downto 0));
   bh67_wm31_2_c4 <= tile_14_filtered_output_c4(0);
   bh67_wm30_3_c4 <= tile_14_filtered_output_c4(1);
   bh67_wm29_4_c4 <= tile_14_filtered_output_c4(2);
   bh67_wm28_6_c4 <= tile_14_filtered_output_c4(3);
   bh67_wm27_6_c4 <= tile_14_filtered_output_c4(4);
   tile_15_X_c4 <= X(19 downto 17);
   tile_15_Y_c4 <= Y(15 downto 14);
   tile_15_mult: IntMultiplierLUT_3x2_Freq300_uid141
      port map ( clk  => clk,
                 X => tile_15_X_c4,
                 Y => tile_15_Y_c4,
                 R => tile_15_output_c4);

   tile_15_filtered_output_c4 <= unsigned(tile_15_output_c4(4 downto 0));
   bh67_wm34_1_c4 <= tile_15_filtered_output_c4(0);
   bh67_wm33_1_c4 <= tile_15_filtered_output_c4(1);
   bh67_wm32_2_c4 <= tile_15_filtered_output_c4(2);
   bh67_wm31_3_c4 <= tile_15_filtered_output_c4(3);
   bh67_wm30_4_c4 <= tile_15_filtered_output_c4(4);
   tile_16_X_c4 <= X(24 downto 23);
   tile_16_Y_c4 <= Y(13 downto 12);
   tile_16_mult: IntMultiplierLUT_2_signedx2_Freq300_uid146
      port map ( clk  => clk,
                 X => tile_16_X_c4,
                 Y => tile_16_Y_c4,
                 R => tile_16_output_c4);

   tile_16_filtered_output_c4 <= signed(tile_16_output_c4(3 downto 0));
   bh67_wm30_5_c4 <= tile_16_filtered_output_c4(0);
   bh67_wm29_5_c4 <= tile_16_filtered_output_c4(1);
   bh67_wm28_7_c4 <= tile_16_filtered_output_c4(2);
   bh67_wm27_7_c4 <= not tile_16_filtered_output_c4(3);
   tile_17_X_c4 <= X(22 downto 20);
   tile_17_Y_c4 <= Y(13 downto 12);
   tile_17_mult: IntMultiplierLUT_3x2_Freq300_uid151
      port map ( clk  => clk,
                 X => tile_17_X_c4,
                 Y => tile_17_Y_c4,
                 R => tile_17_output_c4);

   tile_17_filtered_output_c4 <= unsigned(tile_17_output_c4(4 downto 0));
   bh67_wm33_2_c4 <= tile_17_filtered_output_c4(0);
   bh67_wm32_3_c4 <= tile_17_filtered_output_c4(1);
   bh67_wm31_4_c4 <= tile_17_filtered_output_c4(2);
   bh67_wm30_6_c4 <= tile_17_filtered_output_c4(3);
   bh67_wm29_6_c4 <= tile_17_filtered_output_c4(4);
   tile_18_X_c4 <= X(19 downto 17);
   tile_18_Y_c4 <= Y(13 downto 12);
   tile_18_mult: IntMultiplierLUT_3x2_Freq300_uid156
      port map ( clk  => clk,
                 X => tile_18_X_c4,
                 Y => tile_18_Y_c4,
                 R => tile_18_output_c4);

   tile_18_filtered_output_c4 <= unsigned(tile_18_output_c4(4 downto 0));
   bh67_wm36_1_c4 <= tile_18_filtered_output_c4(0);
   bh67_wm35_1_c4 <= tile_18_filtered_output_c4(1);
   bh67_wm34_2_c4 <= tile_18_filtered_output_c4(2);
   bh67_wm33_3_c4 <= tile_18_filtered_output_c4(3);
   bh67_wm32_4_c4 <= tile_18_filtered_output_c4(4);
   tile_19_X_c4 <= X(24 downto 23);
   tile_19_Y_c4 <= Y(11 downto 10);
   tile_19_mult: IntMultiplierLUT_2_signedx2_Freq300_uid161
      port map ( clk  => clk,
                 X => tile_19_X_c4,
                 Y => tile_19_Y_c4,
                 R => tile_19_output_c4);

   tile_19_filtered_output_c4 <= signed(tile_19_output_c4(3 downto 0));
   bh67_wm32_5_c4 <= tile_19_filtered_output_c4(0);
   bh67_wm31_5_c4 <= tile_19_filtered_output_c4(1);
   bh67_wm30_7_c4 <= tile_19_filtered_output_c4(2);
   bh67_wm29_7_c4 <= not tile_19_filtered_output_c4(3);
   tile_20_X_c4 <= X(22 downto 20);
   tile_20_Y_c4 <= Y(11 downto 10);
   tile_20_mult: IntMultiplierLUT_3x2_Freq300_uid166
      port map ( clk  => clk,
                 X => tile_20_X_c4,
                 Y => tile_20_Y_c4,
                 R => tile_20_output_c4);

   tile_20_filtered_output_c4 <= unsigned(tile_20_output_c4(4 downto 0));
   bh67_wm35_2_c4 <= tile_20_filtered_output_c4(0);
   bh67_wm34_3_c4 <= tile_20_filtered_output_c4(1);
   bh67_wm33_4_c4 <= tile_20_filtered_output_c4(2);
   bh67_wm32_6_c4 <= tile_20_filtered_output_c4(3);
   bh67_wm31_6_c4 <= tile_20_filtered_output_c4(4);
   tile_21_X_c4 <= X(19 downto 17);
   tile_21_Y_c4 <= Y(11 downto 10);
   tile_21_mult: IntMultiplierLUT_3x2_Freq300_uid171
      port map ( clk  => clk,
                 X => tile_21_X_c4,
                 Y => tile_21_Y_c4,
                 R => tile_21_output_c4);

   tile_21_filtered_output_c4 <= unsigned(tile_21_output_c4(4 downto 0));
   bh67_wm38_1_c4 <= tile_21_filtered_output_c4(0);
   bh67_wm37_1_c4 <= tile_21_filtered_output_c4(1);
   bh67_wm36_2_c4 <= tile_21_filtered_output_c4(2);
   bh67_wm35_3_c4 <= tile_21_filtered_output_c4(3);
   bh67_wm34_4_c4 <= tile_21_filtered_output_c4(4);
   tile_22_X_c4 <= X(24 downto 23);
   tile_22_Y_c4 <= Y(9 downto 8);
   tile_22_mult: IntMultiplierLUT_2_signedx2_Freq300_uid176
      port map ( clk  => clk,
                 X => tile_22_X_c4,
                 Y => tile_22_Y_c4,
                 R => tile_22_output_c4);

   tile_22_filtered_output_c4 <= signed(tile_22_output_c4(3 downto 0));
   bh67_wm34_5_c4 <= tile_22_filtered_output_c4(0);
   bh67_wm33_5_c4 <= tile_22_filtered_output_c4(1);
   bh67_wm32_7_c4 <= tile_22_filtered_output_c4(2);
   bh67_wm31_7_c4 <= not tile_22_filtered_output_c4(3);
   tile_23_X_c4 <= X(22 downto 20);
   tile_23_Y_c4 <= Y(9 downto 8);
   tile_23_mult: IntMultiplierLUT_3x2_Freq300_uid181
      port map ( clk  => clk,
                 X => tile_23_X_c4,
                 Y => tile_23_Y_c4,
                 R => tile_23_output_c4);

   tile_23_filtered_output_c4 <= unsigned(tile_23_output_c4(4 downto 0));
   bh67_wm37_2_c4 <= tile_23_filtered_output_c4(0);
   bh67_wm36_3_c4 <= tile_23_filtered_output_c4(1);
   bh67_wm35_4_c4 <= tile_23_filtered_output_c4(2);
   bh67_wm34_6_c4 <= tile_23_filtered_output_c4(3);
   bh67_wm33_6_c4 <= tile_23_filtered_output_c4(4);
   tile_24_X_c4 <= X(19 downto 17);
   tile_24_Y_c4 <= Y(9 downto 8);
   tile_24_mult: IntMultiplierLUT_3x2_Freq300_uid186
      port map ( clk  => clk,
                 X => tile_24_X_c4,
                 Y => tile_24_Y_c4,
                 R => tile_24_output_c4);

   tile_24_filtered_output_c4 <= unsigned(tile_24_output_c4(4 downto 0));
   bh67_wm40_1_c4 <= tile_24_filtered_output_c4(0);
   bh67_wm39_1_c4 <= tile_24_filtered_output_c4(1);
   bh67_wm38_2_c4 <= tile_24_filtered_output_c4(2);
   bh67_wm37_3_c4 <= tile_24_filtered_output_c4(3);
   bh67_wm36_4_c4 <= tile_24_filtered_output_c4(4);
   tile_25_X_c4 <= X(24 downto 23);
   tile_25_Y_c4 <= Y(7 downto 6);
   tile_25_mult: IntMultiplierLUT_2_signedx2_Freq300_uid191
      port map ( clk  => clk,
                 X => tile_25_X_c4,
                 Y => tile_25_Y_c4,
                 R => tile_25_output_c4);

   tile_25_filtered_output_c4 <= signed(tile_25_output_c4(3 downto 0));
   bh67_wm36_5_c4 <= tile_25_filtered_output_c4(0);
   bh67_wm35_5_c4 <= tile_25_filtered_output_c4(1);
   bh67_wm34_7_c4 <= tile_25_filtered_output_c4(2);
   bh67_wm33_7_c4 <= not tile_25_filtered_output_c4(3);
   tile_26_X_c4 <= X(22 downto 20);
   tile_26_Y_c4 <= Y(7 downto 6);
   tile_26_mult: IntMultiplierLUT_3x2_Freq300_uid196
      port map ( clk  => clk,
                 X => tile_26_X_c4,
                 Y => tile_26_Y_c4,
                 R => tile_26_output_c4);

   tile_26_filtered_output_c4 <= unsigned(tile_26_output_c4(4 downto 0));
   bh67_wm39_2_c4 <= tile_26_filtered_output_c4(0);
   bh67_wm38_3_c4 <= tile_26_filtered_output_c4(1);
   bh67_wm37_4_c4 <= tile_26_filtered_output_c4(2);
   bh67_wm36_6_c4 <= tile_26_filtered_output_c4(3);
   bh67_wm35_6_c4 <= tile_26_filtered_output_c4(4);
   tile_27_X_c4 <= X(19 downto 17);
   tile_27_Y_c4 <= Y(7 downto 6);
   tile_27_mult: IntMultiplierLUT_3x2_Freq300_uid201
      port map ( clk  => clk,
                 X => tile_27_X_c4,
                 Y => tile_27_Y_c4,
                 R => tile_27_output_c4);

   tile_27_filtered_output_c4 <= unsigned(tile_27_output_c4(4 downto 0));
   bh67_wm42_1_c4 <= tile_27_filtered_output_c4(0);
   bh67_wm41_1_c4 <= tile_27_filtered_output_c4(1);
   bh67_wm40_2_c4 <= tile_27_filtered_output_c4(2);
   bh67_wm39_3_c4 <= tile_27_filtered_output_c4(3);
   bh67_wm38_4_c4 <= tile_27_filtered_output_c4(4);
   tile_28_X_c4 <= X(24 downto 23);
   tile_28_Y_c4 <= Y(5 downto 4);
   tile_28_mult: IntMultiplierLUT_2_signedx2_Freq300_uid206
      port map ( clk  => clk,
                 X => tile_28_X_c4,
                 Y => tile_28_Y_c4,
                 R => tile_28_output_c4);

   tile_28_filtered_output_c4 <= signed(tile_28_output_c4(3 downto 0));
   bh67_wm38_5_c4 <= tile_28_filtered_output_c4(0);
   bh67_wm37_5_c4 <= tile_28_filtered_output_c4(1);
   bh67_wm36_7_c4 <= tile_28_filtered_output_c4(2);
   bh67_wm35_7_c4 <= not tile_28_filtered_output_c4(3);
   tile_29_X_c4 <= X(22 downto 20);
   tile_29_Y_c4 <= Y(5 downto 4);
   tile_29_mult: IntMultiplierLUT_3x2_Freq300_uid211
      port map ( clk  => clk,
                 X => tile_29_X_c4,
                 Y => tile_29_Y_c4,
                 R => tile_29_output_c4);

   tile_29_filtered_output_c4 <= unsigned(tile_29_output_c4(4 downto 0));
   bh67_wm41_2_c4 <= tile_29_filtered_output_c4(0);
   bh67_wm40_3_c4 <= tile_29_filtered_output_c4(1);
   bh67_wm39_4_c4 <= tile_29_filtered_output_c4(2);
   bh67_wm38_6_c4 <= tile_29_filtered_output_c4(3);
   bh67_wm37_6_c4 <= tile_29_filtered_output_c4(4);
   tile_30_X_c4 <= X(19 downto 17);
   tile_30_Y_c4 <= Y(5 downto 4);
   tile_30_mult: IntMultiplierLUT_3x2_Freq300_uid216
      port map ( clk  => clk,
                 X => tile_30_X_c4,
                 Y => tile_30_Y_c4,
                 R => tile_30_output_c4);

   tile_30_filtered_output_c4 <= unsigned(tile_30_output_c4(4 downto 0));
   bh67_wm44_1_c4 <= tile_30_filtered_output_c4(0);
   bh67_wm43_1_c4 <= tile_30_filtered_output_c4(1);
   bh67_wm42_2_c4 <= tile_30_filtered_output_c4(2);
   bh67_wm41_3_c4 <= tile_30_filtered_output_c4(3);
   bh67_wm40_4_c4 <= tile_30_filtered_output_c4(4);
   tile_31_X_c4 <= X(24 downto 23);
   tile_31_Y_c4 <= Y(3 downto 2);
   tile_31_mult: IntMultiplierLUT_2_signedx2_Freq300_uid221
      port map ( clk  => clk,
                 X => tile_31_X_c4,
                 Y => tile_31_Y_c4,
                 R => tile_31_output_c4);

   tile_31_filtered_output_c4 <= signed(tile_31_output_c4(3 downto 0));
   bh67_wm40_5_c4 <= tile_31_filtered_output_c4(0);
   bh67_wm39_5_c4 <= tile_31_filtered_output_c4(1);
   bh67_wm38_7_c4 <= tile_31_filtered_output_c4(2);
   bh67_wm37_7_c4 <= not tile_31_filtered_output_c4(3);
   tile_32_X_c4 <= X(22 downto 20);
   tile_32_Y_c4 <= Y(3 downto 2);
   tile_32_mult: IntMultiplierLUT_3x2_Freq300_uid226
      port map ( clk  => clk,
                 X => tile_32_X_c4,
                 Y => tile_32_Y_c4,
                 R => tile_32_output_c4);

   tile_32_filtered_output_c4 <= unsigned(tile_32_output_c4(4 downto 0));
   bh67_wm43_2_c4 <= tile_32_filtered_output_c4(0);
   bh67_wm42_3_c4 <= tile_32_filtered_output_c4(1);
   bh67_wm41_4_c4 <= tile_32_filtered_output_c4(2);
   bh67_wm40_6_c4 <= tile_32_filtered_output_c4(3);
   bh67_wm39_6_c4 <= tile_32_filtered_output_c4(4);
   tile_33_X_c4 <= X(19 downto 17);
   tile_33_Y_c4 <= Y(3 downto 2);
   tile_33_mult: IntMultiplierLUT_3x2_Freq300_uid231
      port map ( clk  => clk,
                 X => tile_33_X_c4,
                 Y => tile_33_Y_c4,
                 R => tile_33_output_c4);

   tile_33_filtered_output_c4 <= unsigned(tile_33_output_c4(4 downto 0));
   bh67_wm46_1_c4 <= tile_33_filtered_output_c4(0);
   bh67_wm45_1_c4 <= tile_33_filtered_output_c4(1);
   bh67_wm44_2_c4 <= tile_33_filtered_output_c4(2);
   bh67_wm43_3_c4 <= tile_33_filtered_output_c4(3);
   bh67_wm42_4_c4 <= tile_33_filtered_output_c4(4);
   tile_34_X_c4 <= X(24 downto 23);
   tile_34_Y_c4 <= Y(1 downto 0);
   tile_34_mult: IntMultiplierLUT_2_signedx2_Freq300_uid236
      port map ( clk  => clk,
                 X => tile_34_X_c4,
                 Y => tile_34_Y_c4,
                 R => tile_34_output_c4);

   tile_34_filtered_output_c4 <= signed(tile_34_output_c4(3 downto 0));
   bh67_wm42_5_c4 <= tile_34_filtered_output_c4(0);
   bh67_wm41_5_c4 <= tile_34_filtered_output_c4(1);
   bh67_wm40_7_c4 <= tile_34_filtered_output_c4(2);
   bh67_wm39_7_c4 <= not tile_34_filtered_output_c4(3);
   tile_35_X_c4 <= X(22 downto 20);
   tile_35_Y_c4 <= Y(1 downto 0);
   tile_35_mult: IntMultiplierLUT_3x2_Freq300_uid241
      port map ( clk  => clk,
                 X => tile_35_X_c4,
                 Y => tile_35_Y_c4,
                 R => tile_35_output_c4);

   tile_35_filtered_output_c4 <= unsigned(tile_35_output_c4(4 downto 0));
   bh67_wm45_2_c4 <= tile_35_filtered_output_c4(0);
   bh67_wm44_3_c4 <= tile_35_filtered_output_c4(1);
   bh67_wm43_4_c4 <= tile_35_filtered_output_c4(2);
   bh67_wm42_6_c4 <= tile_35_filtered_output_c4(3);
   bh67_wm41_6_c4 <= tile_35_filtered_output_c4(4);
   tile_36_X_c4 <= X(19 downto 17);
   tile_36_Y_c4 <= Y(1 downto 0);
   tile_36_mult: IntMultiplierLUT_3x2_Freq300_uid246
      port map ( clk  => clk,
                 X => tile_36_X_c4,
                 Y => tile_36_Y_c4,
                 R => tile_36_output_c4);

   tile_36_filtered_output_c4 <= unsigned(tile_36_output_c4(4 downto 0));
   bh67_wm48_1_c4 <= tile_36_filtered_output_c4(0);
   bh67_wm47_1_c4 <= tile_36_filtered_output_c4(1);
   bh67_wm46_2_c4 <= tile_36_filtered_output_c4(2);
   bh67_wm45_3_c4 <= tile_36_filtered_output_c4(3);
   bh67_wm44_4_c4 <= tile_36_filtered_output_c4(4);
   tile_37_X_c4 <= X(16 downto 16);
   tile_37_Y_c4 <= Y(24 downto 24);
   tile_37_mult: IntMultiplierLUT_1x1_signed_Freq300_uid251
      port map ( clk  => clk,
                 X => tile_37_X_c4,
                 Y => tile_37_Y_c4,
                 R => tile_37_output_c4);

   tile_37_filtered_output_c4 <= signed(tile_37_output_c4(0 downto 0));
   bh67_wm25_8_c4 <= not tile_37_filtered_output_c4(0);
   tile_38_X_c4 <= X(15 downto 12);
   tile_38_Y_c4 <= Y(24 downto 24);
   tile_38_mult: IntMultiplierLUT_4x1_signed_Freq300_uid253
      port map ( clk  => clk,
                 X => tile_38_X_c4,
                 Y => tile_38_Y_c4,
                 R => tile_38_output_c4);

   tile_38_filtered_output_c4 <= signed(tile_38_output_c4(4 downto 0));
   bh67_wm29_8_c4 <= tile_38_filtered_output_c4(0);
   bh67_wm28_8_c4 <= tile_38_filtered_output_c4(1);
   bh67_wm27_8_c4 <= tile_38_filtered_output_c4(2);
   bh67_wm26_8_c4 <= tile_38_filtered_output_c4(3);
   bh67_wm25_9_c4 <= not tile_38_filtered_output_c4(4);
   tile_39_X_c4 <= X(11 downto 8);
   tile_39_Y_c4 <= Y(24 downto 24);
   tile_39_mult: IntMultiplierLUT_4x1_signed_Freq300_uid258
      port map ( clk  => clk,
                 X => tile_39_X_c4,
                 Y => tile_39_Y_c4,
                 R => tile_39_output_c4);

   tile_39_filtered_output_c4 <= signed(tile_39_output_c4(4 downto 0));
   bh67_wm33_8_c4 <= tile_39_filtered_output_c4(0);
   bh67_wm32_8_c4 <= tile_39_filtered_output_c4(1);
   bh67_wm31_8_c4 <= tile_39_filtered_output_c4(2);
   bh67_wm30_8_c4 <= tile_39_filtered_output_c4(3);
   bh67_wm29_9_c4 <= not tile_39_filtered_output_c4(4);
   tile_40_X_c4 <= X(7 downto 4);
   tile_40_Y_c4 <= Y(24 downto 24);
   tile_40_mult: IntMultiplierLUT_4x1_signed_Freq300_uid263
      port map ( clk  => clk,
                 X => tile_40_X_c4,
                 Y => tile_40_Y_c4,
                 R => tile_40_output_c4);

   tile_40_filtered_output_c4 <= signed(tile_40_output_c4(4 downto 0));
   bh67_wm37_8_c4 <= tile_40_filtered_output_c4(0);
   bh67_wm36_8_c4 <= tile_40_filtered_output_c4(1);
   bh67_wm35_8_c4 <= tile_40_filtered_output_c4(2);
   bh67_wm34_8_c4 <= tile_40_filtered_output_c4(3);
   bh67_wm33_9_c4 <= not tile_40_filtered_output_c4(4);
   tile_41_X_c4 <= X(3 downto 0);
   tile_41_Y_c4 <= Y(24 downto 24);
   tile_41_mult: IntMultiplierLUT_4x1_signed_Freq300_uid268
      port map ( clk  => clk,
                 X => tile_41_X_c4,
                 Y => tile_41_Y_c4,
                 R => tile_41_output_c4);

   tile_41_filtered_output_c4 <= signed(tile_41_output_c4(4 downto 0));
   bh67_wm41_7_c4 <= tile_41_filtered_output_c4(0);
   bh67_wm40_8_c4 <= tile_41_filtered_output_c4(1);
   bh67_wm39_8_c4 <= tile_41_filtered_output_c4(2);
   bh67_wm38_8_c4 <= tile_41_filtered_output_c4(3);
   bh67_wm37_9_c4 <= not tile_41_filtered_output_c4(4);
   tile_42_X_c4 <= X(24 downto 21);
   tile_42_Y_c4 <= Y(24 downto 24);
   tile_42_mult: IntMultiplierLUT_4_signedx1_signed_Freq300_uid273
      port map ( clk  => clk,
                 X => tile_42_X_c4,
                 Y => tile_42_Y_c4,
                 R => tile_42_output_c4);

   tile_42_filtered_output_c4 <= signed(tile_42_output_c4(4 downto 0));
   bh67_wm20_3_c4 <= tile_42_filtered_output_c4(0);
   bh67_wm19_3_c4 <= tile_42_filtered_output_c4(1);
   bh67_wm18_1_c4 <= tile_42_filtered_output_c4(2);
   bh67_wm17_1_c4 <= tile_42_filtered_output_c4(3);
   bh67_wm16_0_c4 <= not tile_42_filtered_output_c4(4);
   tile_43_X_c4 <= X(20 downto 17);
   tile_43_Y_c4 <= Y(24 downto 24);
   tile_43_mult: IntMultiplierLUT_4x1_signed_Freq300_uid278
      port map ( clk  => clk,
                 X => tile_43_X_c4,
                 Y => tile_43_Y_c4,
                 R => tile_43_output_c4);

   tile_43_filtered_output_c4 <= signed(tile_43_output_c4(4 downto 0));
   bh67_wm24_6_c4 <= tile_43_filtered_output_c4(0);
   bh67_wm23_6_c4 <= tile_43_filtered_output_c4(1);
   bh67_wm22_5_c4 <= tile_43_filtered_output_c4(2);
   bh67_wm21_4_c4 <= tile_43_filtered_output_c4(3);
   bh67_wm20_4_c4 <= not tile_43_filtered_output_c4(4);
   bh67_wm41_8_c4 <= AA_c4(0);
   bh67_wm40_9_c4 <= AA_c4(1);
   bh67_wm39_9_c4 <= AA_c4(2);
   bh67_wm38_9_c4 <= AA_c4(3);
   bh67_wm37_10_c4 <= AA_c4(4);
   bh67_wm36_9_c4 <= AA_c4(5);
   bh67_wm35_9_c4 <= AA_c4(6);
   bh67_wm34_9_c4 <= AA_c4(7);
   bh67_wm33_10_c4 <= AA_c4(8);
   bh67_wm32_9_c4 <= AA_c4(9);
   bh67_wm31_9_c4 <= AA_c4(10);
   bh67_wm30_9_c4 <= AA_c4(11);
   bh67_wm29_10_c4 <= AA_c4(12);
   bh67_wm28_9_c4 <= AA_c4(13);
   bh67_wm27_9_c4 <= AA_c4(14);
   bh67_wm26_9_c4 <= AA_c4(15);
   bh67_wm25_10_c4 <= AA_c4(16);
   bh67_wm24_7_c4 <= AA_c4(17);
   bh67_wm23_7_c4 <= AA_c4(18);
   bh67_wm22_6_c4 <= AA_c4(19);
   bh67_wm21_5_c4 <= AA_c4(20);
   bh67_wm20_5_c4 <= AA_c4(21);
   bh67_wm19_4_c4 <= AA_c4(22);
   bh67_wm18_2_c4 <= AA_c4(23);
   bh67_wm17_2_c4 <= AA_c4(24);
   bh67_wm16_1_c4 <= AA_c4(25);
   bh67_wm15_0_c4 <= AA_c4(26);
   bh67_wm14_0_c4 <= AA_c4(27);
   bh67_wm13_0_c4 <= AA_c4(28);
   bh67_wm12_0_c4 <= AA_c4(29);
   bh67_wm11_0_c4 <= AA_c4(30);
   bh67_wm10_0_c4 <= AA_c4(31);
   bh67_wm9_0_c4 <= AA_c4(32);

   -- Adding the constant bits 
   bh67_wm42_7_c0 <= '1';
   bh67_wm39_10_c0 <= '1';
   bh67_wm38_10_c0 <= '1';
   bh67_wm37_11_c0 <= '1';
   bh67_wm34_10_c0 <= '1';
   bh67_wm33_11_c0 <= '1';
   bh67_wm30_10_c0 <= '1';
   bh67_wm29_11_c0 <= '1';
   bh67_wm26_10_c0 <= '1';
   bh67_wm22_7_c0 <= '1';
   bh67_wm18_3_c0 <= '1';
   bh67_wm15_1_c0 <= '1';
   bh67_wm14_1_c0 <= '1';
   bh67_wm13_1_c0 <= '1';
   bh67_wm12_1_c0 <= '1';
   bh67_wm11_1_c0 <= '1';
   bh67_wm10_1_c0 <= '1';
   bh67_wm9_1_c0 <= '1';


   Compressor_23_3_Freq300_uid284_bh67_uid285_In0_c5 <= "" & bh67_wm48_0_c5 & bh67_wm48_1_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid285_In1_c5 <= "" & bh67_wm47_0_c5 & bh67_wm47_1_c5;
   bh67_wm48_2_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid285_Out0_c5(0);
   bh67_wm47_2_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid285_Out0_c5(1);
   bh67_wm46_3_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid285_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid285: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid285_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid285_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid285_Out0_copy286_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid285_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid285_Out0_copy286_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid289_In0_c5 <= "" & bh67_wm46_0_c5 & bh67_wm46_1_c5 & bh67_wm46_2_c5;
   bh67_wm46_4_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid289_Out0_c5(0);
   bh67_wm45_4_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid289_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid289: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid289_In0_c5,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid289_Out0_copy290_c5);
   Compressor_3_2_Freq300_uid288_bh67_uid289_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid289_Out0_copy290_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid293_In0_c5 <= "" & bh67_wm45_0_c5 & bh67_wm45_1_c5 & bh67_wm45_2_c5 & bh67_wm45_3_c5;
   Compressor_14_3_Freq300_uid292_bh67_uid293_In1_c5 <= "" & bh67_wm44_0_c5;
   bh67_wm45_5_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid293_Out0_c5(0);
   bh67_wm44_5_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid293_Out0_c5(1);
   bh67_wm43_5_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid293_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid293: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid293_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid293_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid293_Out0_copy294_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid293_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid293_Out0_copy294_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid295_In0_c4 <= "" & bh67_wm44_1_c4 & bh67_wm44_2_c4 & bh67_wm44_3_c4 & bh67_wm44_4_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid295_In1_c5 <= "" & bh67_wm43_0_c5;
   bh67_wm44_6_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid295_Out0_c5(0);
   bh67_wm43_6_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid295_Out0_c5(1);
   bh67_wm42_8_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid295_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid295: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid295_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid295_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid295_Out0_copy296_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid295_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid295_Out0_copy296_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid297_In0_c4 <= "" & bh67_wm43_1_c4 & bh67_wm43_2_c4 & bh67_wm43_3_c4 & bh67_wm43_4_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid297_In1_c5 <= "" & bh67_wm42_0_c5;
   bh67_wm43_7_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid297_Out0_c5(0);
   bh67_wm42_9_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid297_Out0_c5(1);
   bh67_wm41_9_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid297_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid297: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid297_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid297_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid297_Out0_copy298_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid297_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid297_Out0_copy298_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid301_In0_c4 <= "" & bh67_wm42_1_c4 & bh67_wm42_2_c4 & bh67_wm42_3_c4 & bh67_wm42_4_c4 & bh67_wm42_5_c4 & bh67_wm42_6_c4;
   bh67_wm42_10_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid301_Out0_c4(0);
   bh67_wm41_10_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid301_Out0_c4(1);
   bh67_wm40_10_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid301_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid301: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid301_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid301_Out0_copy302_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid301_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid301_Out0_copy302_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid303_In0_c5 <= "" & bh67_wm41_0_c5 & bh67_wm41_1_c5 & bh67_wm41_2_c5 & bh67_wm41_3_c5 & bh67_wm41_4_c5 & bh67_wm41_5_c5;
   bh67_wm41_11_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid303_Out0_c5(0);
   bh67_wm40_11_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid303_Out0_c5(1);
   bh67_wm39_11_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid303_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid303: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid303_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid303_Out0_copy304_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid303_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid303_Out0_copy304_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid305_In0_c4 <= "" & bh67_wm41_6_c4 & bh67_wm41_7_c4 & bh67_wm41_8_c4;
   bh67_wm41_12_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid305_Out0_c4(0);
   bh67_wm40_12_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid305_Out0_c4(1);
   Compressor_3_2_Freq300_uid288_uid305: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid305_In0_c4,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid305_Out0_copy306_c4);
   Compressor_3_2_Freq300_uid288_bh67_uid305_Out0_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid305_Out0_copy306_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid307_In0_c5 <= "" & bh67_wm40_0_c5 & bh67_wm40_1_c5 & bh67_wm40_2_c5 & bh67_wm40_3_c5 & bh67_wm40_4_c5 & bh67_wm40_5_c5;
   bh67_wm40_13_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid307_Out0_c5(0);
   bh67_wm39_12_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid307_Out0_c5(1);
   bh67_wm38_11_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid307_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid307: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid307_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid307_Out0_copy308_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid307_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid307_Out0_copy308_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid309_In0_c4 <= "" & bh67_wm40_6_c4 & bh67_wm40_7_c4 & bh67_wm40_8_c4 & bh67_wm40_9_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid309_In1_c5 <= "" & bh67_wm39_0_c5;
   bh67_wm40_14_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid309_Out0_c5(0);
   bh67_wm39_13_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid309_Out0_c5(1);
   bh67_wm38_12_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid309_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid309: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid309_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid309_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid309_Out0_copy310_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid309_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid309_Out0_copy310_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid311_In0_c4 <= "" & bh67_wm39_1_c4 & bh67_wm39_2_c4 & bh67_wm39_3_c4 & bh67_wm39_4_c4 & bh67_wm39_5_c4 & bh67_wm39_6_c4;
   bh67_wm39_14_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid311_Out0_c4(0);
   bh67_wm38_13_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid311_Out0_c4(1);
   bh67_wm37_12_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid311_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid311: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid311_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid311_Out0_copy312_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid311_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid311_Out0_copy312_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid313_In0_c4 <= "" & bh67_wm39_7_c4 & bh67_wm39_8_c4 & bh67_wm39_9_c4 & bh67_wm39_10_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid313_In1_c5 <= "" & bh67_wm38_0_c5;
   bh67_wm39_15_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid313_Out0_c5(0);
   bh67_wm38_14_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid313_Out0_c5(1);
   bh67_wm37_13_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid313_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid313: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid313_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid313_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid313_Out0_copy314_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid313_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid313_Out0_copy314_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid315_In0_c4 <= "" & bh67_wm38_1_c4 & bh67_wm38_2_c4 & bh67_wm38_3_c4 & bh67_wm38_4_c4 & bh67_wm38_5_c4 & bh67_wm38_6_c4;
   bh67_wm38_15_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid315_Out0_c4(0);
   bh67_wm37_14_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid315_Out0_c4(1);
   bh67_wm36_10_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid315_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid315: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid315_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid315_Out0_copy316_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid315_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid315_Out0_copy316_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid317_In0_c4 <= "" & bh67_wm38_7_c4 & bh67_wm38_8_c4 & bh67_wm38_9_c4;
   bh67_wm38_16_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid317_Out0_c4(0);
   bh67_wm37_15_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid317_Out0_c4(1);
   Compressor_3_2_Freq300_uid288_uid317: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid317_In0_c4,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid317_Out0_copy318_c4);
   Compressor_3_2_Freq300_uid288_bh67_uid317_Out0_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid317_Out0_copy318_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid319_In0_c5 <= "" & bh67_wm37_0_c5 & bh67_wm37_1_c5 & bh67_wm37_2_c5 & bh67_wm37_3_c5 & bh67_wm37_4_c5 & bh67_wm37_5_c5;
   bh67_wm37_16_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid319_Out0_c5(0);
   bh67_wm36_11_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid319_Out0_c5(1);
   bh67_wm35_10_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid319_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid319: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid319_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid319_Out0_copy320_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid319_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid319_Out0_copy320_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid321_In0_c4 <= "" & bh67_wm37_8_c4 & bh67_wm37_11_c4 & bh67_wm37_10_c4 & bh67_wm37_9_c4 & bh67_wm37_7_c4 & bh67_wm37_6_c4;
   bh67_wm37_17_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid321_Out0_c4(0);
   bh67_wm36_12_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid321_Out0_c4(1);
   bh67_wm35_11_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid321_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid321: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid321_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid321_Out0_copy322_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid321_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid321_Out0_copy322_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid323_In0_c5 <= "" & bh67_wm36_0_c5 & bh67_wm36_1_c5 & bh67_wm36_2_c5 & bh67_wm36_3_c5 & bh67_wm36_4_c5 & bh67_wm36_5_c5;
   bh67_wm36_13_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid323_Out0_c5(0);
   bh67_wm35_12_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid323_Out0_c5(1);
   bh67_wm34_11_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid323_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid323: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid323_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid323_Out0_copy324_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid323_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid323_Out0_copy324_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid325_In0_c4 <= "" & bh67_wm36_6_c4 & bh67_wm36_7_c4 & bh67_wm36_8_c4 & bh67_wm36_9_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid325_In1_c5 <= "" & bh67_wm35_0_c5;
   bh67_wm36_14_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid325_Out0_c5(0);
   bh67_wm35_13_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid325_Out0_c5(1);
   bh67_wm34_12_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid325_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid325: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid325_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid325_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid325_Out0_copy326_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid325_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid325_Out0_copy326_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid327_In0_c4 <= "" & bh67_wm35_1_c4 & bh67_wm35_2_c4 & bh67_wm35_3_c4 & bh67_wm35_4_c4 & bh67_wm35_5_c4 & bh67_wm35_6_c4;
   bh67_wm35_14_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid327_Out0_c4(0);
   bh67_wm34_13_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid327_Out0_c4(1);
   bh67_wm33_12_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid327_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid327: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid327_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid327_Out0_copy328_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid327_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid327_Out0_copy328_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid329_In0_c4 <= "" & bh67_wm35_7_c4 & bh67_wm35_8_c4 & bh67_wm35_9_c4;
   bh67_wm35_15_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid329_Out0_c4(0);
   bh67_wm34_14_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid329_Out0_c4(1);
   Compressor_3_2_Freq300_uid288_uid329: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid329_In0_c4,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid329_Out0_copy330_c4);
   Compressor_3_2_Freq300_uid288_bh67_uid329_Out0_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid329_Out0_copy330_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid331_In0_c5 <= "" & bh67_wm34_0_c5 & bh67_wm34_1_c5 & bh67_wm34_2_c5 & bh67_wm34_3_c5 & bh67_wm34_4_c5 & bh67_wm34_5_c5;
   bh67_wm34_15_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid331_Out0_c5(0);
   bh67_wm33_13_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid331_Out0_c5(1);
   bh67_wm32_10_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid331_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid331: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid331_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid331_Out0_copy332_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid331_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid331_Out0_copy332_c5; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid334_bh67_uid335_In0_c4 <= "" & bh67_wm34_6_c4 & bh67_wm34_7_c4 & bh67_wm34_8_c4 & bh67_wm34_9_c4 & bh67_wm34_10_c4;
   bh67_wm34_16_c4 <= Compressor_5_3_Freq300_uid334_bh67_uid335_Out0_c4(0);
   bh67_wm33_14_c4 <= Compressor_5_3_Freq300_uid334_bh67_uid335_Out0_c4(1);
   bh67_wm32_11_c4 <= Compressor_5_3_Freq300_uid334_bh67_uid335_Out0_c4(2);
   Compressor_5_3_Freq300_uid334_uid335: Compressor_5_3_Freq300_uid334
      port map ( X0 => Compressor_5_3_Freq300_uid334_bh67_uid335_In0_c4,
                 R => Compressor_5_3_Freq300_uid334_bh67_uid335_Out0_copy336_c4);
   Compressor_5_3_Freq300_uid334_bh67_uid335_Out0_c4 <= Compressor_5_3_Freq300_uid334_bh67_uid335_Out0_copy336_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid337_In0_c5 <= "" & bh67_wm33_0_c5 & bh67_wm33_1_c5 & bh67_wm33_2_c5 & bh67_wm33_3_c5 & bh67_wm33_4_c5 & bh67_wm33_5_c5;
   bh67_wm33_15_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid337_Out0_c5(0);
   bh67_wm32_12_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid337_Out0_c5(1);
   bh67_wm31_10_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid337_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid337: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid337_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid337_Out0_copy338_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid337_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid337_Out0_copy338_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid339_In0_c4 <= "" & bh67_wm33_6_c4 & bh67_wm33_7_c4 & bh67_wm33_8_c4 & bh67_wm33_9_c4 & bh67_wm33_10_c4 & bh67_wm33_11_c4;
   bh67_wm33_16_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid339_Out0_c4(0);
   bh67_wm32_13_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid339_Out0_c4(1);
   bh67_wm31_11_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid339_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid339: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid339_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid339_Out0_copy340_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid339_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid339_Out0_copy340_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid341_In0_c5 <= "" & bh67_wm32_0_c5 & bh67_wm32_1_c5 & bh67_wm32_2_c5 & bh67_wm32_3_c5 & bh67_wm32_4_c5 & bh67_wm32_5_c5;
   bh67_wm32_14_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid341_Out0_c5(0);
   bh67_wm31_12_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid341_Out0_c5(1);
   bh67_wm30_11_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid341_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid341: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid341_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid341_Out0_copy342_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid341_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid341_Out0_copy342_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid343_In0_c4 <= "" & bh67_wm32_6_c4 & bh67_wm32_7_c4 & bh67_wm32_8_c4 & bh67_wm32_9_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid343_In1_c5 <= "" & bh67_wm31_0_c5;
   bh67_wm32_15_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid343_Out0_c5(0);
   bh67_wm31_13_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid343_Out0_c5(1);
   bh67_wm30_12_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid343_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid343: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid343_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid343_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid343_Out0_copy344_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid343_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid343_Out0_copy344_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid345_In0_c4 <= "" & bh67_wm31_1_c4 & bh67_wm31_2_c4 & bh67_wm31_3_c4 & bh67_wm31_4_c4 & bh67_wm31_5_c4 & bh67_wm31_6_c4;
   bh67_wm31_14_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid345_Out0_c4(0);
   bh67_wm30_13_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid345_Out0_c4(1);
   bh67_wm29_12_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid345_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid345: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid345_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid345_Out0_copy346_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid345_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid345_Out0_copy346_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid347_In0_c4 <= "" & bh67_wm31_7_c4 & bh67_wm31_8_c4 & bh67_wm31_9_c4;
   bh67_wm31_15_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid347_Out0_c4(0);
   bh67_wm30_14_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid347_Out0_c4(1);
   Compressor_3_2_Freq300_uid288_uid347: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid347_In0_c4,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid347_Out0_copy348_c4);
   Compressor_3_2_Freq300_uid288_bh67_uid347_Out0_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid347_Out0_copy348_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid349_In0_c5 <= "" & bh67_wm30_0_c5 & bh67_wm30_1_c5 & bh67_wm30_2_c5 & bh67_wm30_3_c5 & bh67_wm30_4_c5 & bh67_wm30_5_c5;
   bh67_wm30_15_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid349_Out0_c5(0);
   bh67_wm29_13_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid349_Out0_c5(1);
   bh67_wm28_10_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid349_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid349: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid349_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid349_Out0_copy350_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid349_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid349_Out0_copy350_c5; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid334_bh67_uid351_In0_c4 <= "" & bh67_wm30_6_c4 & bh67_wm30_7_c4 & bh67_wm30_8_c4 & bh67_wm30_9_c4 & bh67_wm30_10_c4;
   bh67_wm30_16_c4 <= Compressor_5_3_Freq300_uid334_bh67_uid351_Out0_c4(0);
   bh67_wm29_14_c4 <= Compressor_5_3_Freq300_uid334_bh67_uid351_Out0_c4(1);
   bh67_wm28_11_c4 <= Compressor_5_3_Freq300_uid334_bh67_uid351_Out0_c4(2);
   Compressor_5_3_Freq300_uid334_uid351: Compressor_5_3_Freq300_uid334
      port map ( X0 => Compressor_5_3_Freq300_uid334_bh67_uid351_In0_c4,
                 R => Compressor_5_3_Freq300_uid334_bh67_uid351_Out0_copy352_c4);
   Compressor_5_3_Freq300_uid334_bh67_uid351_Out0_c4 <= Compressor_5_3_Freq300_uid334_bh67_uid351_Out0_copy352_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid353_In0_c5 <= "" & bh67_wm29_0_c5 & bh67_wm29_1_c5 & bh67_wm29_2_c5 & bh67_wm29_3_c5 & bh67_wm29_4_c5 & bh67_wm29_5_c5;
   bh67_wm29_15_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid353_Out0_c5(0);
   bh67_wm28_12_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid353_Out0_c5(1);
   bh67_wm27_10_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid353_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid353: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid353_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid353_Out0_copy354_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid353_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid353_Out0_copy354_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid355_In0_c4 <= "" & bh67_wm29_6_c4 & bh67_wm29_7_c4 & bh67_wm29_8_c4 & bh67_wm29_9_c4 & bh67_wm29_10_c4 & bh67_wm29_11_c4;
   bh67_wm29_16_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid355_Out0_c4(0);
   bh67_wm28_13_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid355_Out0_c4(1);
   bh67_wm27_11_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid355_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid355: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid355_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid355_Out0_copy356_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid355_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid355_Out0_copy356_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid357_In0_c5 <= "" & bh67_wm28_0_c5 & bh67_wm28_1_c5 & bh67_wm28_2_c5 & bh67_wm28_3_c5 & bh67_wm28_4_c5 & bh67_wm28_5_c5;
   bh67_wm28_14_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid357_Out0_c5(0);
   bh67_wm27_12_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid357_Out0_c5(1);
   bh67_wm26_11_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid357_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid357: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid357_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid357_Out0_copy358_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid357_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid357_Out0_copy358_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid359_In0_c4 <= "" & bh67_wm28_6_c4 & bh67_wm28_7_c4 & bh67_wm28_8_c4 & bh67_wm28_9_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid359_In1_c5 <= "" & bh67_wm27_0_c5;
   bh67_wm28_15_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid359_Out0_c5(0);
   bh67_wm27_13_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid359_Out0_c5(1);
   bh67_wm26_12_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid359_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid359: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid359_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid359_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid359_Out0_copy360_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid359_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid359_Out0_copy360_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid361_In0_c4 <= "" & bh67_wm27_1_c4 & bh67_wm27_2_c4 & bh67_wm27_3_c4 & bh67_wm27_4_c4 & bh67_wm27_5_c4 & bh67_wm27_6_c4;
   bh67_wm27_14_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid361_Out0_c4(0);
   bh67_wm26_13_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid361_Out0_c4(1);
   bh67_wm25_11_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid361_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid361: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid361_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid361_Out0_copy362_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid361_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid361_Out0_copy362_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid363_In0_c4 <= "" & bh67_wm27_7_c4 & bh67_wm27_8_c4 & bh67_wm27_9_c4;
   bh67_wm27_15_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid363_Out0_c4(0);
   bh67_wm26_14_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid363_Out0_c4(1);
   Compressor_3_2_Freq300_uid288_uid363: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid363_In0_c4,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid363_Out0_copy364_c4);
   Compressor_3_2_Freq300_uid288_bh67_uid363_Out0_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid363_Out0_copy364_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid365_In0_c5 <= "" & bh67_wm26_0_c5 & bh67_wm26_1_c5 & bh67_wm26_2_c5 & bh67_wm26_3_c5 & bh67_wm26_4_c5 & bh67_wm26_5_c5;
   bh67_wm26_15_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid365_Out0_c5(0);
   bh67_wm25_12_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid365_Out0_c5(1);
   bh67_wm24_8_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid365_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid365: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid365_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid365_Out0_copy366_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid365_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid365_Out0_copy366_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid367_In0_c4 <= "" & bh67_wm26_6_c4 & bh67_wm26_7_c4 & bh67_wm26_8_c4 & bh67_wm26_9_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid367_In1_c5 <= "" & bh67_wm25_0_c5;
   bh67_wm26_16_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid367_Out0_c5(0);
   bh67_wm25_13_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid367_Out0_c5(1);
   bh67_wm24_9_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid367_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid367: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid367_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid367_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid367_Out0_copy368_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid367_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid367_Out0_copy368_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid369_In0_c4 <= "" & bh67_wm25_1_c4 & bh67_wm25_2_c4 & bh67_wm25_3_c4 & bh67_wm25_4_c4 & bh67_wm25_5_c4 & bh67_wm25_6_c4;
   bh67_wm25_14_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid369_Out0_c4(0);
   bh67_wm24_10_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid369_Out0_c4(1);
   bh67_wm23_8_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid369_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid369: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid369_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid369_Out0_copy370_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid369_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid369_Out0_copy370_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid371_In0_c4 <= "" & bh67_wm25_7_c4 & bh67_wm25_8_c4 & bh67_wm25_9_c4 & bh67_wm25_10_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid371_In1_c4 <= "" & bh67_wm24_0_c4;
   bh67_wm25_15_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid371_Out0_c4(0);
   bh67_wm24_11_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid371_Out0_c4(1);
   bh67_wm23_9_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid371_Out0_c4(2);
   Compressor_14_3_Freq300_uid292_uid371: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid371_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid371_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid371_Out0_copy372_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid371_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid371_Out0_copy372_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid373_In0_c4 <= "" & bh67_wm24_1_c4 & bh67_wm24_2_c4 & bh67_wm24_3_c4 & bh67_wm24_4_c4 & bh67_wm24_5_c4 & bh67_wm24_6_c4;
   bh67_wm24_12_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid373_Out0_c4(0);
   bh67_wm23_10_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid373_Out0_c4(1);
   bh67_wm22_8_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid373_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid373: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid373_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid373_Out0_copy374_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid373_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid373_Out0_copy374_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid375_In0_c4 <= "" & bh67_wm23_0_c4 & bh67_wm23_1_c4 & bh67_wm23_2_c4 & bh67_wm23_3_c4 & bh67_wm23_4_c4 & "0";
   bh67_wm23_11_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid375_Out0_c4(0);
   bh67_wm22_9_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid375_Out0_c4(1);
   bh67_wm21_6_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid375_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid375: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid375_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid375_Out0_copy376_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid375_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid375_Out0_copy376_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid377_In0_c4 <= "" & bh67_wm23_5_c4 & bh67_wm23_6_c4 & bh67_wm23_7_c4;
   Compressor_23_3_Freq300_uid284_bh67_uid377_In1_c4 <= "" & bh67_wm22_0_c4 & bh67_wm22_1_c4;
   bh67_wm23_12_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid377_Out0_c4(0);
   bh67_wm22_10_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid377_Out0_c4(1);
   bh67_wm21_7_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid377_Out0_c4(2);
   Compressor_23_3_Freq300_uid284_uid377: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid377_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid377_In1_c4,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid377_Out0_copy378_c4);
   Compressor_23_3_Freq300_uid284_bh67_uid377_Out0_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid377_Out0_copy378_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid379_In0_c4 <= "" & bh67_wm22_2_c4 & bh67_wm22_3_c4 & bh67_wm22_4_c4 & bh67_wm22_5_c4 & bh67_wm22_6_c4 & bh67_wm22_7_c4;
   bh67_wm22_11_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid379_Out0_c4(0);
   bh67_wm21_8_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid379_Out0_c4(1);
   bh67_wm20_6_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid379_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid379: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid379_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid379_Out0_copy380_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid379_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid379_Out0_copy380_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid381_In0_c4 <= "" & bh67_wm21_0_c4 & bh67_wm21_1_c4 & bh67_wm21_2_c4 & bh67_wm21_3_c4 & bh67_wm21_4_c4 & bh67_wm21_5_c4;
   bh67_wm21_9_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid381_Out0_c4(0);
   bh67_wm20_7_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid381_Out0_c4(1);
   bh67_wm19_5_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid381_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid381: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid381_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid381_Out0_copy382_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid381_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid381_Out0_copy382_c4; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid383_In0_c4 <= "" & bh67_wm20_0_c4 & bh67_wm20_1_c4 & bh67_wm20_2_c4 & bh67_wm20_3_c4 & bh67_wm20_4_c4 & bh67_wm20_5_c4;
   bh67_wm20_8_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid383_Out0_c4(0);
   bh67_wm19_6_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid383_Out0_c4(1);
   bh67_wm18_4_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid383_Out0_c4(2);
   Compressor_6_3_Freq300_uid300_uid383: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid383_In0_c4,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid383_Out0_copy384_c4);
   Compressor_6_3_Freq300_uid300_bh67_uid383_Out0_c4 <= Compressor_6_3_Freq300_uid300_bh67_uid383_Out0_copy384_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid385_In0_c4 <= "" & bh67_wm19_0_c4 & bh67_wm19_1_c4 & bh67_wm19_2_c4 & bh67_wm19_3_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid385_In1_c4 <= "" & bh67_wm18_0_c4;
   bh67_wm19_7_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid385_Out0_c4(0);
   bh67_wm18_5_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid385_Out0_c4(1);
   bh67_wm17_3_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid385_Out0_c4(2);
   Compressor_14_3_Freq300_uid292_uid385: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid385_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid385_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid385_Out0_copy386_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid385_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid385_Out0_copy386_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid387_In0_c4 <= "" & bh67_wm18_1_c4 & bh67_wm18_2_c4 & bh67_wm18_3_c4;
   Compressor_23_3_Freq300_uid284_bh67_uid387_In1_c4 <= "" & bh67_wm17_0_c4 & bh67_wm17_1_c4;
   bh67_wm18_6_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid387_Out0_c4(0);
   bh67_wm17_4_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid387_Out0_c4(1);
   bh67_wm16_2_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid387_Out0_c4(2);
   Compressor_23_3_Freq300_uid284_uid387: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid387_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid387_In1_c4,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid387_Out0_copy388_c4);
   Compressor_23_3_Freq300_uid284_bh67_uid387_Out0_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid387_Out0_copy388_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid389_In0_c4 <= "" & bh67_wm16_0_c4 & bh67_wm16_1_c4 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid389_In1_c4 <= "" & bh67_wm15_0_c4 & bh67_wm15_1_c4;
   bh67_wm16_3_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid389_Out0_c4(0);
   bh67_wm15_2_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid389_Out0_c4(1);
   bh67_wm14_2_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid389_Out0_c4(2);
   Compressor_23_3_Freq300_uid284_uid389: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid389_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid389_In1_c4,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid389_Out0_copy390_c4);
   Compressor_23_3_Freq300_uid284_bh67_uid389_Out0_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid389_Out0_copy390_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid391_In0_c4 <= "" & bh67_wm14_0_c4 & bh67_wm14_1_c4 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid391_In1_c4 <= "" & bh67_wm13_0_c4 & bh67_wm13_1_c4;
   bh67_wm14_3_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid391_Out0_c4(0);
   bh67_wm13_2_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid391_Out0_c4(1);
   bh67_wm12_2_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid391_Out0_c4(2);
   Compressor_23_3_Freq300_uid284_uid391: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid391_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid391_In1_c4,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid391_Out0_copy392_c4);
   Compressor_23_3_Freq300_uid284_bh67_uid391_Out0_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid391_Out0_copy392_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid393_In0_c4 <= "" & bh67_wm12_0_c4 & bh67_wm12_1_c4 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid393_In1_c4 <= "" & bh67_wm11_0_c4 & bh67_wm11_1_c4;
   bh67_wm12_3_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid393_Out0_c4(0);
   bh67_wm11_2_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid393_Out0_c4(1);
   bh67_wm10_2_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid393_Out0_c4(2);
   Compressor_23_3_Freq300_uid284_uid393: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid393_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid393_In1_c4,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid393_Out0_copy394_c4);
   Compressor_23_3_Freq300_uid284_bh67_uid393_Out0_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid393_Out0_copy394_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid395_In0_c4 <= "" & bh67_wm10_0_c4 & bh67_wm10_1_c4 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid395_In1_c4 <= "" & bh67_wm9_0_c4 & bh67_wm9_1_c4;
   bh67_wm10_3_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid395_Out0_c4(0);
   bh67_wm9_2_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid395_Out0_c4(1);
   Compressor_23_3_Freq300_uid284_uid395: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid395_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid395_In1_c4,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid395_Out0_copy396_c4);
   Compressor_23_3_Freq300_uid284_bh67_uid395_Out0_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid395_Out0_copy396_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid397_In0_c5 <= "" & bh67_wm46_3_c5 & bh67_wm46_4_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid397_In1_c5 <= "" & bh67_wm45_4_c5 & bh67_wm45_5_c5;
   bh67_wm46_5_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid397_Out0_c5(0);
   bh67_wm45_6_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid397_Out0_c5(1);
   bh67_wm44_7_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid397_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid397: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid397_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid397_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid397_Out0_copy398_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid397_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid397_Out0_copy398_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid399_In0_c5 <= "" & bh67_wm44_5_c5 & bh67_wm44_6_c5 & "0";
   bh67_wm44_8_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid399_Out0_c5(0);
   bh67_wm43_8_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid399_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid399: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid399_In0_c5,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid399_Out0_copy400_c5);
   Compressor_3_2_Freq300_uid288_bh67_uid399_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid399_Out0_copy400_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid401_In0_c5 <= "" & bh67_wm43_5_c5 & bh67_wm43_6_c5 & bh67_wm43_7_c5;
   bh67_wm43_9_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid401_Out0_c5(0);
   bh67_wm42_11_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid401_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid401: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid401_In0_c5,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid401_Out0_copy402_c5);
   Compressor_3_2_Freq300_uid288_bh67_uid401_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid401_Out0_copy402_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid403_In0_c5 <= "" & bh67_wm42_7_c5 & bh67_wm42_8_c5 & bh67_wm42_9_c5 & bh67_wm42_10_c5;
   Compressor_14_3_Freq300_uid292_bh67_uid403_In1_c5 <= "" & bh67_wm41_9_c5;
   bh67_wm42_12_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid403_Out0_c5(0);
   bh67_wm41_13_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid403_Out0_c5(1);
   bh67_wm40_15_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid403_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid403: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid403_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid403_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid403_Out0_copy404_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid403_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid403_Out0_copy404_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid405_In0_c5 <= "" & bh67_wm41_10_c5 & bh67_wm41_11_c5 & bh67_wm41_12_c5;
   bh67_wm41_14_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid405_Out0_c5(0);
   bh67_wm40_16_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid405_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid405: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid405_In0_c5,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid405_Out0_copy406_c5);
   Compressor_3_2_Freq300_uid288_bh67_uid405_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid405_Out0_copy406_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid407_In0_c5 <= "" & bh67_wm40_10_c5 & bh67_wm40_11_c5 & bh67_wm40_12_c5 & bh67_wm40_13_c5;
   Compressor_14_3_Freq300_uid292_bh67_uid407_In1_c5 <= "" & bh67_wm39_11_c5;
   bh67_wm40_17_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid407_Out0_c5(0);
   bh67_wm39_16_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid407_Out0_c5(1);
   bh67_wm38_17_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid407_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid407: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid407_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid407_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid407_Out0_copy408_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid407_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid407_Out0_copy408_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid409_In0_c5 <= "" & bh67_wm39_12_c5 & bh67_wm39_13_c5 & bh67_wm39_14_c5 & bh67_wm39_15_c5;
   Compressor_14_3_Freq300_uid292_bh67_uid409_In1_c4 <= "" & bh67_wm38_16_c4;
   bh67_wm39_17_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid409_Out0_c5(0);
   bh67_wm38_18_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid409_Out0_c5(1);
   bh67_wm37_18_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid409_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid409: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid409_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid409_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid409_Out0_copy410_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid409_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid409_Out0_copy410_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid411_In0_c5 <= "" & bh67_wm38_15_c5 & bh67_wm38_14_c5 & bh67_wm38_13_c5 & bh67_wm38_12_c5 & bh67_wm38_11_c5 & bh67_wm38_10_c5;
   bh67_wm38_19_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid411_Out0_c5(0);
   bh67_wm37_19_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid411_Out0_c5(1);
   bh67_wm36_15_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid411_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid411: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid411_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid411_Out0_copy412_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid411_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid411_Out0_copy412_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid413_In0_c5 <= "" & bh67_wm37_17_c5 & bh67_wm37_12_c5 & bh67_wm37_13_c5 & bh67_wm37_14_c5 & bh67_wm37_15_c5 & bh67_wm37_16_c5;
   bh67_wm37_20_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid413_Out0_c5(0);
   bh67_wm36_16_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid413_Out0_c5(1);
   bh67_wm35_16_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid413_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid413: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid413_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid413_Out0_copy414_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid413_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid413_Out0_copy414_c5; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid334_bh67_uid415_In0_c5 <= "" & bh67_wm36_10_c5 & bh67_wm36_11_c5 & bh67_wm36_12_c5 & bh67_wm36_13_c5 & bh67_wm36_14_c5;
   bh67_wm36_17_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid415_Out0_c5(0);
   bh67_wm35_17_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid415_Out0_c5(1);
   bh67_wm34_17_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid415_Out0_c5(2);
   Compressor_5_3_Freq300_uid334_uid415: Compressor_5_3_Freq300_uid334
      port map ( X0 => Compressor_5_3_Freq300_uid334_bh67_uid415_In0_c5,
                 R => Compressor_5_3_Freq300_uid334_bh67_uid415_Out0_copy416_c5);
   Compressor_5_3_Freq300_uid334_bh67_uid415_Out0_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid415_Out0_copy416_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid417_In0_c5 <= "" & bh67_wm35_10_c5 & bh67_wm35_11_c5 & bh67_wm35_12_c5 & bh67_wm35_13_c5 & bh67_wm35_14_c5 & bh67_wm35_15_c5;
   bh67_wm35_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid417_Out0_c5(0);
   bh67_wm34_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid417_Out0_c5(1);
   bh67_wm33_17_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid417_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid417: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid417_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid417_Out0_copy418_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid417_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid417_Out0_copy418_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid419_In0_c5 <= "" & bh67_wm34_16_c5 & bh67_wm34_15_c5 & bh67_wm34_14_c5 & bh67_wm34_13_c5 & bh67_wm34_12_c5 & bh67_wm34_11_c5;
   bh67_wm34_19_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid419_Out0_c5(0);
   bh67_wm33_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid419_Out0_c5(1);
   bh67_wm32_16_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid419_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid419: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid419_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid419_Out0_copy420_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid419_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid419_Out0_copy420_c5; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid334_bh67_uid421_In0_c5 <= "" & bh67_wm33_16_c5 & bh67_wm33_15_c5 & bh67_wm33_14_c5 & bh67_wm33_13_c5 & bh67_wm33_12_c5;
   bh67_wm33_19_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid421_Out0_c5(0);
   bh67_wm32_17_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid421_Out0_c5(1);
   bh67_wm31_16_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid421_Out0_c5(2);
   Compressor_5_3_Freq300_uid334_uid421: Compressor_5_3_Freq300_uid334
      port map ( X0 => Compressor_5_3_Freq300_uid334_bh67_uid421_In0_c5,
                 R => Compressor_5_3_Freq300_uid334_bh67_uid421_Out0_copy422_c5);
   Compressor_5_3_Freq300_uid334_bh67_uid421_Out0_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid421_Out0_copy422_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid423_In0_c5 <= "" & bh67_wm32_10_c5 & bh67_wm32_11_c5 & bh67_wm32_12_c5 & bh67_wm32_13_c5 & bh67_wm32_14_c5 & bh67_wm32_15_c5;
   bh67_wm32_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid423_Out0_c5(0);
   bh67_wm31_17_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid423_Out0_c5(1);
   bh67_wm30_17_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid423_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid423: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid423_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid423_Out0_copy424_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid423_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid423_Out0_copy424_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid425_In0_c5 <= "" & bh67_wm31_10_c5 & bh67_wm31_11_c5 & bh67_wm31_12_c5 & bh67_wm31_13_c5 & bh67_wm31_14_c5 & bh67_wm31_15_c5;
   bh67_wm31_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid425_Out0_c5(0);
   bh67_wm30_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid425_Out0_c5(1);
   bh67_wm29_17_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid425_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid425: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid425_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid425_Out0_copy426_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid425_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid425_Out0_copy426_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid427_In0_c5 <= "" & bh67_wm30_16_c5 & bh67_wm30_15_c5 & bh67_wm30_14_c5 & bh67_wm30_13_c5 & bh67_wm30_12_c5 & bh67_wm30_11_c5;
   bh67_wm30_19_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid427_Out0_c5(0);
   bh67_wm29_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid427_Out0_c5(1);
   bh67_wm28_16_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid427_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid427: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid427_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid427_Out0_copy428_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid427_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid427_Out0_copy428_c5; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid334_bh67_uid429_In0_c5 <= "" & bh67_wm29_16_c5 & bh67_wm29_15_c5 & bh67_wm29_14_c5 & bh67_wm29_13_c5 & bh67_wm29_12_c5;
   bh67_wm29_19_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid429_Out0_c5(0);
   bh67_wm28_17_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid429_Out0_c5(1);
   bh67_wm27_16_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid429_Out0_c5(2);
   Compressor_5_3_Freq300_uid334_uid429: Compressor_5_3_Freq300_uid334
      port map ( X0 => Compressor_5_3_Freq300_uid334_bh67_uid429_In0_c5,
                 R => Compressor_5_3_Freq300_uid334_bh67_uid429_Out0_copy430_c5);
   Compressor_5_3_Freq300_uid334_bh67_uid429_Out0_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid429_Out0_copy430_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid431_In0_c5 <= "" & bh67_wm28_10_c5 & bh67_wm28_11_c5 & bh67_wm28_12_c5 & bh67_wm28_13_c5 & bh67_wm28_14_c5 & bh67_wm28_15_c5;
   bh67_wm28_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid431_Out0_c5(0);
   bh67_wm27_17_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid431_Out0_c5(1);
   bh67_wm26_17_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid431_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid431: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid431_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid431_Out0_copy432_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid431_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid431_Out0_copy432_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid433_In0_c5 <= "" & bh67_wm27_10_c5 & bh67_wm27_11_c5 & bh67_wm27_12_c5 & bh67_wm27_13_c5 & bh67_wm27_14_c5 & bh67_wm27_15_c5;
   bh67_wm27_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid433_Out0_c5(0);
   bh67_wm26_18_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid433_Out0_c5(1);
   bh67_wm25_16_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid433_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid433: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid433_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid433_Out0_copy434_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid433_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid433_Out0_copy434_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid435_In0_c5 <= "" & bh67_wm26_16_c5 & bh67_wm26_15_c5 & bh67_wm26_14_c5 & bh67_wm26_13_c5 & bh67_wm26_12_c5 & bh67_wm26_11_c5;
   bh67_wm26_19_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid435_Out0_c5(0);
   bh67_wm25_17_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid435_Out0_c5(1);
   bh67_wm24_13_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid435_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid435: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid435_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid435_Out0_copy436_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid435_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid435_Out0_copy436_c5; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid334_bh67_uid437_In0_c5 <= "" & bh67_wm25_11_c5 & bh67_wm25_12_c5 & bh67_wm25_13_c5 & bh67_wm25_14_c5 & bh67_wm25_15_c5;
   bh67_wm25_18_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid437_Out0_c5(0);
   bh67_wm24_14_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid437_Out0_c5(1);
   bh67_wm23_13_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid437_Out0_c5(2);
   Compressor_5_3_Freq300_uid334_uid437: Compressor_5_3_Freq300_uid334
      port map ( X0 => Compressor_5_3_Freq300_uid334_bh67_uid437_In0_c5,
                 R => Compressor_5_3_Freq300_uid334_bh67_uid437_Out0_copy438_c5);
   Compressor_5_3_Freq300_uid334_bh67_uid437_Out0_c5 <= Compressor_5_3_Freq300_uid334_bh67_uid437_Out0_copy438_c5; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid300_bh67_uid439_In0_c5 <= "" & bh67_wm24_7_c5 & bh67_wm24_8_c5 & bh67_wm24_9_c5 & bh67_wm24_10_c5 & bh67_wm24_11_c5 & bh67_wm24_12_c5;
   bh67_wm24_15_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid439_Out0_c5(0);
   bh67_wm23_14_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid439_Out0_c5(1);
   bh67_wm22_12_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid439_Out0_c5(2);
   Compressor_6_3_Freq300_uid300_uid439: Compressor_6_3_Freq300_uid300
      port map ( X0 => Compressor_6_3_Freq300_uid300_bh67_uid439_In0_c5,
                 R => Compressor_6_3_Freq300_uid300_bh67_uid439_Out0_copy440_c5);
   Compressor_6_3_Freq300_uid300_bh67_uid439_Out0_c5 <= Compressor_6_3_Freq300_uid300_bh67_uid439_Out0_copy440_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid441_In0_c4 <= "" & bh67_wm23_8_c4 & bh67_wm23_9_c4 & bh67_wm23_10_c4 & bh67_wm23_11_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid441_In1_c4 <= "" & bh67_wm22_8_c4;
   bh67_wm23_15_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid441_Out0_c4(0);
   bh67_wm22_13_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid441_Out0_c4(1);
   bh67_wm21_10_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid441_Out0_c4(2);
   Compressor_14_3_Freq300_uid292_uid441: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid441_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid441_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid441_Out0_copy442_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid441_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid441_Out0_copy442_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid443_In0_c4 <= "" & bh67_wm22_9_c4 & bh67_wm22_10_c4 & bh67_wm22_11_c4;
   bh67_wm22_14_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid443_Out0_c4(0);
   bh67_wm21_11_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid443_Out0_c4(1);
   Compressor_3_2_Freq300_uid288_uid443: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid443_In0_c4,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid443_Out0_copy444_c4);
   Compressor_3_2_Freq300_uid288_bh67_uid443_Out0_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid443_Out0_copy444_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid445_In0_c4 <= "" & bh67_wm21_6_c4 & bh67_wm21_7_c4 & bh67_wm21_8_c4 & bh67_wm21_9_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid445_In1_c0 <= "" & "0";
   bh67_wm21_12_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid445_Out0_c4(0);
   bh67_wm20_9_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid445_Out0_c4(1);
   bh67_wm19_8_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid445_Out0_c4(2);
   Compressor_14_3_Freq300_uid292_uid445: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid445_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid445_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid445_Out0_copy446_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid445_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid445_Out0_copy446_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid447_In0_c4 <= "" & bh67_wm20_6_c4 & bh67_wm20_7_c4 & bh67_wm20_8_c4;
   bh67_wm20_10_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid447_Out0_c4(0);
   bh67_wm19_9_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid447_Out0_c4(1);
   Compressor_3_2_Freq300_uid288_uid447: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid447_In0_c4,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid447_Out0_copy448_c4);
   Compressor_3_2_Freq300_uid288_bh67_uid447_Out0_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid447_Out0_copy448_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid449_In0_c4 <= "" & bh67_wm19_4_c4 & bh67_wm19_5_c4 & bh67_wm19_6_c4 & bh67_wm19_7_c4;
   Compressor_14_3_Freq300_uid292_bh67_uid449_In1_c0 <= "" & "0";
   bh67_wm19_10_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid449_Out0_c4(0);
   bh67_wm18_7_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid449_Out0_c4(1);
   bh67_wm17_5_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid449_Out0_c4(2);
   Compressor_14_3_Freq300_uid292_uid449: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid449_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid449_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid449_Out0_copy450_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid449_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid449_Out0_copy450_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid451_In0_c4 <= "" & bh67_wm18_4_c4 & bh67_wm18_5_c4 & bh67_wm18_6_c4;
   bh67_wm18_8_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid451_Out0_c4(0);
   bh67_wm17_6_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid451_Out0_c4(1);
   Compressor_3_2_Freq300_uid288_uid451: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid451_In0_c4,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid451_Out0_copy452_c4);
   Compressor_3_2_Freq300_uid288_bh67_uid451_Out0_c4 <= Compressor_3_2_Freq300_uid288_bh67_uid451_Out0_copy452_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid453_In0_c4 <= "" & bh67_wm17_2_c4 & bh67_wm17_3_c4 & bh67_wm17_4_c4;
   Compressor_23_3_Freq300_uid284_bh67_uid453_In1_c4 <= "" & bh67_wm16_2_c4 & bh67_wm16_3_c4;
   bh67_wm17_7_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid453_Out0_c4(0);
   bh67_wm16_4_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid453_Out0_c4(1);
   bh67_wm15_3_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid453_Out0_c4(2);
   Compressor_23_3_Freq300_uid284_uid453: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid453_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid453_In1_c4,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid453_Out0_copy454_c4);
   Compressor_23_3_Freq300_uid284_bh67_uid453_Out0_c4 <= Compressor_23_3_Freq300_uid284_bh67_uid453_Out0_copy454_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid455_In0_c4 <= "" & bh67_wm14_2_c4 & bh67_wm14_3_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid455_In1_c4 <= "" & bh67_wm13_2_c4;
   bh67_wm14_4_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid455_Out0_c4(0);
   bh67_wm13_3_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid455_Out0_c4(1);
   bh67_wm12_4_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid455_Out0_c4(2);
   Compressor_14_3_Freq300_uid292_uid455: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid455_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid455_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid455_Out0_copy456_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid455_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid455_Out0_copy456_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid457_In0_c4 <= "" & bh67_wm12_2_c4 & bh67_wm12_3_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid457_In1_c4 <= "" & bh67_wm11_2_c4;
   bh67_wm12_5_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid457_Out0_c4(0);
   bh67_wm11_3_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid457_Out0_c4(1);
   bh67_wm10_4_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid457_Out0_c4(2);
   Compressor_14_3_Freq300_uid292_uid457: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid457_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid457_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid457_Out0_copy458_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid457_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid457_Out0_copy458_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid459_In0_c4 <= "" & bh67_wm10_2_c4 & bh67_wm10_3_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid459_In1_c4 <= "" & bh67_wm9_2_c4;
   bh67_wm10_5_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid459_Out0_c4(0);
   bh67_wm9_3_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid459_Out0_c4(1);
   Compressor_14_3_Freq300_uid292_uid459: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid459_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid459_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid459_Out0_copy460_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid459_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid459_Out0_copy460_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid461_In0_c5 <= "" & bh67_wm44_7_c5 & bh67_wm44_8_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid461_In1_c5 <= "" & bh67_wm43_8_c5 & bh67_wm43_9_c5;
   bh67_wm44_9_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid461_Out0_c5(0);
   bh67_wm43_10_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid461_Out0_c5(1);
   bh67_wm42_13_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid461_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid461: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid461_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid461_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid461_Out0_copy462_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid461_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid461_Out0_copy462_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid463_In0_c5 <= "" & bh67_wm42_11_c5 & bh67_wm42_12_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid463_In1_c5 <= "" & bh67_wm41_13_c5 & bh67_wm41_14_c5;
   bh67_wm42_14_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid463_Out0_c5(0);
   bh67_wm41_15_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid463_Out0_c5(1);
   bh67_wm40_18_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid463_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid463: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid463_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid463_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid463_Out0_copy464_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid463_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid463_Out0_copy464_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid465_In0_c5 <= "" & bh67_wm40_14_c5 & bh67_wm40_15_c5 & bh67_wm40_16_c5 & bh67_wm40_17_c5;
   Compressor_14_3_Freq300_uid292_bh67_uid465_In1_c5 <= "" & bh67_wm39_16_c5;
   bh67_wm40_19_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid465_Out0_c5(0);
   bh67_wm39_18_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid465_Out0_c5(1);
   bh67_wm38_20_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid465_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid465: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid465_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid465_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid465_Out0_copy466_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid465_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid465_Out0_copy466_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid467_In0_c5 <= "" & bh67_wm38_17_c5 & bh67_wm38_18_c5 & bh67_wm38_19_c5;
   Compressor_23_3_Freq300_uid284_bh67_uid467_In1_c5 <= "" & bh67_wm37_18_c5 & bh67_wm37_19_c5;
   bh67_wm38_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid467_Out0_c5(0);
   bh67_wm37_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid467_Out0_c5(1);
   bh67_wm36_18_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid467_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid467: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid467_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid467_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid467_Out0_copy468_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid467_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid467_Out0_copy468_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid469_In0_c5 <= "" & bh67_wm36_15_c5 & bh67_wm36_16_c5 & bh67_wm36_17_c5;
   Compressor_23_3_Freq300_uid284_bh67_uid469_In1_c5 <= "" & bh67_wm35_16_c5 & bh67_wm35_17_c5;
   bh67_wm36_19_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid469_Out0_c5(0);
   bh67_wm35_19_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid469_Out0_c5(1);
   bh67_wm34_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid469_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid469: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid469_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid469_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid469_Out0_copy470_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid469_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid469_Out0_copy470_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid471_In0_c5 <= "" & bh67_wm34_17_c5 & bh67_wm34_18_c5 & bh67_wm34_19_c5;
   Compressor_23_3_Freq300_uid284_bh67_uid471_In1_c5 <= "" & bh67_wm33_17_c5 & bh67_wm33_18_c5;
   bh67_wm34_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid471_Out0_c5(0);
   bh67_wm33_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid471_Out0_c5(1);
   bh67_wm32_19_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid471_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid471: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid471_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid471_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid471_Out0_copy472_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid471_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid471_Out0_copy472_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid473_In0_c5 <= "" & bh67_wm32_16_c5 & bh67_wm32_17_c5 & bh67_wm32_18_c5;
   Compressor_23_3_Freq300_uid284_bh67_uid473_In1_c5 <= "" & bh67_wm31_16_c5 & bh67_wm31_17_c5;
   bh67_wm32_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid473_Out0_c5(0);
   bh67_wm31_19_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid473_Out0_c5(1);
   bh67_wm30_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid473_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid473: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid473_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid473_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid473_Out0_copy474_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid473_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid473_Out0_copy474_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid475_In0_c5 <= "" & bh67_wm30_17_c5 & bh67_wm30_18_c5 & bh67_wm30_19_c5;
   Compressor_23_3_Freq300_uid284_bh67_uid475_In1_c5 <= "" & bh67_wm29_17_c5 & bh67_wm29_18_c5;
   bh67_wm30_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid475_Out0_c5(0);
   bh67_wm29_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid475_Out0_c5(1);
   bh67_wm28_19_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid475_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid475: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid475_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid475_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid475_Out0_copy476_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid475_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid475_Out0_copy476_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid477_In0_c5 <= "" & bh67_wm28_16_c5 & bh67_wm28_17_c5 & bh67_wm28_18_c5;
   Compressor_23_3_Freq300_uid284_bh67_uid477_In1_c5 <= "" & bh67_wm27_16_c5 & bh67_wm27_17_c5;
   bh67_wm28_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid477_Out0_c5(0);
   bh67_wm27_19_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid477_Out0_c5(1);
   bh67_wm26_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid477_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid477: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid477_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid477_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid477_Out0_copy478_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid477_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid477_Out0_copy478_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid479_In0_c5 <= "" & bh67_wm26_10_c5 & bh67_wm26_17_c5 & bh67_wm26_18_c5 & bh67_wm26_19_c5;
   Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c0 <= "" & "0";
   bh67_wm26_21_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid479_Out0_c5(0);
   bh67_wm25_19_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid479_Out0_c5(1);
   bh67_wm24_16_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid479_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid479: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid479_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid479_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid479_Out0_copy480_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid479_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid479_Out0_copy480_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid481_In0_c5 <= "" & bh67_wm25_16_c5 & bh67_wm25_17_c5 & bh67_wm25_18_c5;
   bh67_wm25_20_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid481_Out0_c5(0);
   bh67_wm24_17_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid481_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid481: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid481_In0_c5,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid481_Out0_copy482_c5);
   Compressor_3_2_Freq300_uid288_bh67_uid481_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid481_Out0_copy482_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid483_In0_c5 <= "" & bh67_wm24_13_c5 & bh67_wm24_14_c5 & bh67_wm24_15_c5;
   bh67_wm24_18_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid483_Out0_c5(0);
   bh67_wm23_16_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid483_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid483: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid483_In0_c5,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid483_Out0_copy484_c5);
   Compressor_3_2_Freq300_uid288_bh67_uid483_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid483_Out0_copy484_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid485_In0_c5 <= "" & bh67_wm23_12_c5 & bh67_wm23_13_c5 & bh67_wm23_14_c5 & bh67_wm23_15_c5;
   Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c0 <= "" & "0";
   bh67_wm23_17_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid485_Out0_c5(0);
   bh67_wm22_15_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid485_Out0_c5(1);
   bh67_wm21_13_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid485_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid485: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid485_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid485_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid485_Out0_copy486_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid485_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid485_Out0_copy486_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid487_In0_c5 <= "" & bh67_wm22_12_c5 & bh67_wm22_13_c5 & bh67_wm22_14_c5;
   bh67_wm22_16_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid487_Out0_c5(0);
   bh67_wm21_14_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid487_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid487: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid487_In0_c5,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid487_Out0_copy488_c5);
   Compressor_3_2_Freq300_uid288_bh67_uid487_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid487_Out0_copy488_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid489_In0_c4 <= "" & bh67_wm21_10_c4 & bh67_wm21_11_c4 & bh67_wm21_12_c4;
   Compressor_23_3_Freq300_uid284_bh67_uid489_In1_c4 <= "" & bh67_wm20_9_c4 & bh67_wm20_10_c4;
   bh67_wm21_15_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_c5(0);
   bh67_wm20_11_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_c5(1);
   bh67_wm19_11_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid489: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid489_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid489_In1_c4,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_copy490_c4);
   Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid489_Out0_copy490_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid491_In0_c4 <= "" & bh67_wm19_8_c4 & bh67_wm19_9_c4 & bh67_wm19_10_c4;
   Compressor_23_3_Freq300_uid284_bh67_uid491_In1_c4 <= "" & bh67_wm18_7_c4 & bh67_wm18_8_c4;
   bh67_wm19_12_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_c5(0);
   bh67_wm18_9_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_c5(1);
   bh67_wm17_8_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid491: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid491_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid491_In1_c4,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_copy492_c4);
   Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid491_Out0_copy492_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid493_In0_c4 <= "" & bh67_wm17_5_c4 & bh67_wm17_6_c4 & bh67_wm17_7_c4;
   bh67_wm17_9_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_c5(0);
   bh67_wm16_5_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid493: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid493_In0_c4,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_copy494_c4);
   Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid493_Out0_copy494_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid495_In0_c4 <= "" & bh67_wm15_2_c4 & bh67_wm15_3_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid495_In1_c4 <= "" & bh67_wm14_4_c4;
   bh67_wm15_4_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid495_Out0_c4(0);
   bh67_wm14_5_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid495_Out0_c4(1);
   bh67_wm13_4_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid495_Out0_c4(2);
   Compressor_14_3_Freq300_uid292_uid495: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid495_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid495_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid495_Out0_copy496_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid495_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid495_Out0_copy496_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid497_In0_c4 <= "" & bh67_wm12_4_c4 & bh67_wm12_5_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid497_In1_c4 <= "" & bh67_wm11_3_c4;
   bh67_wm12_6_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid497_Out0_c4(0);
   bh67_wm11_4_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid497_Out0_c4(1);
   bh67_wm10_6_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid497_Out0_c4(2);
   Compressor_14_3_Freq300_uid292_uid497: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid497_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid497_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid497_Out0_copy498_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid497_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid497_Out0_copy498_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid499_In0_c4 <= "" & bh67_wm10_4_c4 & bh67_wm10_5_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid499_In1_c4 <= "" & bh67_wm9_3_c4;
   bh67_wm10_7_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid499_Out0_c4(0);
   bh67_wm9_4_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid499_Out0_c4(1);
   Compressor_14_3_Freq300_uid292_uid499: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid499_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid499_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid499_Out0_copy500_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid499_Out0_c4 <= Compressor_14_3_Freq300_uid292_bh67_uid499_Out0_copy500_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid501_In0_c5 <= "" & bh67_wm42_13_c5 & bh67_wm42_14_c5 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid501_In1_c5 <= "" & bh67_wm41_15_c5;
   bh67_wm42_15_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid501_Out0_c5(0);
   bh67_wm41_16_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid501_Out0_c5(1);
   bh67_wm40_20_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid501_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid501: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid501_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid501_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid501_Out0_copy502_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid501_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid501_Out0_copy502_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid503_In0_c5 <= "" & bh67_wm40_18_c5 & bh67_wm40_19_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid503_In1_c5 <= "" & bh67_wm39_17_c5 & bh67_wm39_18_c5;
   bh67_wm40_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid503_Out0_c5(0);
   bh67_wm39_19_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid503_Out0_c5(1);
   bh67_wm38_22_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid503_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid503: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid503_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid503_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid503_Out0_copy504_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid503_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid503_Out0_copy504_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid505_In0_c5 <= "" & bh67_wm38_20_c5 & bh67_wm38_21_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid505_In1_c5 <= "" & bh67_wm37_20_c5 & bh67_wm37_21_c5;
   bh67_wm38_23_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid505_Out0_c5(0);
   bh67_wm37_22_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid505_Out0_c5(1);
   bh67_wm36_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid505_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid505: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid505_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid505_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid505_Out0_copy506_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid505_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid505_Out0_copy506_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid507_In0_c5 <= "" & bh67_wm36_18_c5 & bh67_wm36_19_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid507_In1_c5 <= "" & bh67_wm35_18_c5 & bh67_wm35_19_c5;
   bh67_wm36_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid507_Out0_c5(0);
   bh67_wm35_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid507_Out0_c5(1);
   bh67_wm34_22_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid507_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid507: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid507_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid507_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid507_Out0_copy508_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid507_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid507_Out0_copy508_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid509_In0_c5 <= "" & bh67_wm34_20_c5 & bh67_wm34_21_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid509_In1_c5 <= "" & bh67_wm33_19_c5 & bh67_wm33_20_c5;
   bh67_wm34_23_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid509_Out0_c5(0);
   bh67_wm33_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid509_Out0_c5(1);
   bh67_wm32_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid509_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid509: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid509_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid509_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid509_Out0_copy510_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid509_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid509_Out0_copy510_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid511_In0_c5 <= "" & bh67_wm32_19_c5 & bh67_wm32_20_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid511_In1_c5 <= "" & bh67_wm31_18_c5 & bh67_wm31_19_c5;
   bh67_wm32_22_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid511_Out0_c5(0);
   bh67_wm31_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid511_Out0_c5(1);
   bh67_wm30_22_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid511_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid511: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid511_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid511_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid511_Out0_copy512_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid511_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid511_Out0_copy512_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid513_In0_c5 <= "" & bh67_wm30_20_c5 & bh67_wm30_21_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid513_In1_c5 <= "" & bh67_wm29_19_c5 & bh67_wm29_20_c5;
   bh67_wm30_23_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid513_Out0_c5(0);
   bh67_wm29_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid513_Out0_c5(1);
   bh67_wm28_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid513_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid513: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid513_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid513_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid513_Out0_copy514_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid513_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid513_Out0_copy514_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid515_In0_c5 <= "" & bh67_wm28_19_c5 & bh67_wm28_20_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid515_In1_c5 <= "" & bh67_wm27_18_c5 & bh67_wm27_19_c5;
   bh67_wm28_22_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid515_Out0_c5(0);
   bh67_wm27_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid515_Out0_c5(1);
   bh67_wm26_22_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid515_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid515: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid515_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid515_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid515_Out0_copy516_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid515_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid515_Out0_copy516_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid517_In0_c5 <= "" & bh67_wm26_20_c5 & bh67_wm26_21_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid517_In1_c5 <= "" & bh67_wm25_19_c5 & bh67_wm25_20_c5;
   bh67_wm26_23_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid517_Out0_c5(0);
   bh67_wm25_21_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid517_Out0_c5(1);
   bh67_wm24_19_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid517_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid517: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid517_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid517_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid517_Out0_copy518_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid517_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid517_Out0_copy518_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid519_In0_c5 <= "" & bh67_wm24_16_c5 & bh67_wm24_17_c5 & bh67_wm24_18_c5;
   Compressor_23_3_Freq300_uid284_bh67_uid519_In1_c5 <= "" & bh67_wm23_16_c5 & bh67_wm23_17_c5;
   bh67_wm24_20_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid519_Out0_c5(0);
   bh67_wm23_18_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid519_Out0_c5(1);
   bh67_wm22_17_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid519_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid519: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid519_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid519_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid519_Out0_copy520_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid519_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid519_Out0_copy520_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid521_In0_c5 <= "" & bh67_wm22_15_c5 & bh67_wm22_16_c5 & "0";
   bh67_wm22_18_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid521_Out0_c5(0);
   bh67_wm21_16_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid521_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid521: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid521_In0_c5,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid521_Out0_copy522_c5);
   Compressor_3_2_Freq300_uid288_bh67_uid521_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid521_Out0_copy522_c5; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid288_bh67_uid523_In0_c5 <= "" & bh67_wm21_13_c5 & bh67_wm21_14_c5 & bh67_wm21_15_c5;
   bh67_wm21_17_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid523_Out0_c5(0);
   bh67_wm20_12_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid523_Out0_c5(1);
   Compressor_3_2_Freq300_uid288_uid523: Compressor_3_2_Freq300_uid288
      port map ( X0 => Compressor_3_2_Freq300_uid288_bh67_uid523_In0_c5,
                 R => Compressor_3_2_Freq300_uid288_bh67_uid523_Out0_copy524_c5);
   Compressor_3_2_Freq300_uid288_bh67_uid523_Out0_c5 <= Compressor_3_2_Freq300_uid288_bh67_uid523_Out0_copy524_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid525_In0_c5 <= "" & bh67_wm19_11_c5 & bh67_wm19_12_c5 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid525_In1_c5 <= "" & bh67_wm18_9_c5;
   bh67_wm19_13_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid525_Out0_c5(0);
   bh67_wm18_10_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid525_Out0_c5(1);
   bh67_wm17_10_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid525_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid525: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid525_In0_c5,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid525_In1_c5,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid525_Out0_copy526_c5);
   Compressor_14_3_Freq300_uid292_bh67_uid525_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid525_Out0_copy526_c5; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid284_bh67_uid527_In0_c5 <= "" & bh67_wm17_8_c5 & bh67_wm17_9_c5 & "0";
   Compressor_23_3_Freq300_uid284_bh67_uid527_In1_c5 <= "" & bh67_wm16_4_c5 & bh67_wm16_5_c5;
   bh67_wm17_11_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid527_Out0_c5(0);
   bh67_wm16_6_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid527_Out0_c5(1);
   bh67_wm15_5_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid527_Out0_c5(2);
   Compressor_23_3_Freq300_uid284_uid527: Compressor_23_3_Freq300_uid284
      port map ( X0 => Compressor_23_3_Freq300_uid284_bh67_uid527_In0_c5,
                 X1 => Compressor_23_3_Freq300_uid284_bh67_uid527_In1_c5,
                 R => Compressor_23_3_Freq300_uid284_bh67_uid527_Out0_copy528_c5);
   Compressor_23_3_Freq300_uid284_bh67_uid527_Out0_c5 <= Compressor_23_3_Freq300_uid284_bh67_uid527_Out0_copy528_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid529_In0_c4 <= "" & bh67_wm13_3_c4 & bh67_wm13_4_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid529_In1_c4 <= "" & bh67_wm12_6_c4;
   bh67_wm13_5_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_c5(0);
   bh67_wm12_7_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_c5(1);
   bh67_wm11_5_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_c5(2);
   Compressor_14_3_Freq300_uid292_uid529: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid529_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid529_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_copy530_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid529_Out0_copy530_c5; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid292_bh67_uid531_In0_c4 <= "" & bh67_wm10_6_c4 & bh67_wm10_7_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid292_bh67_uid531_In1_c4 <= "" & bh67_wm9_4_c4;
   bh67_wm10_8_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_c5(0);
   bh67_wm9_5_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_c5(1);
   Compressor_14_3_Freq300_uid292_uid531: Compressor_14_3_Freq300_uid292
      port map ( X0 => Compressor_14_3_Freq300_uid292_bh67_uid531_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid292_bh67_uid531_In1_c4,
                 R => Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_copy532_c4);
   Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_c5 <= Compressor_14_3_Freq300_uid292_bh67_uid531_Out0_copy532_c5; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh67_24_c5 <= bh67_wm41_16_c5 & bh67_wm42_15_c5 & bh67_wm43_10_c5 & bh67_wm44_9_c5 & bh67_wm45_6_c5 & bh67_wm46_5_c5 & bh67_wm47_2_c5 & bh67_wm48_2_c5 & bh67_wm49_0_c5 & bh67_wm50_0_c5 & bh67_wm51_0_c5 & bh67_wm52_0_c5 & bh67_wm53_0_c5 & bh67_wm54_0_c5 & bh67_wm55_0_c5 & bh67_wm56_0_c5 & bh67_wm57_0_c5 & bh67_wm58_0_c5 & bh67_wm59_0_c5 & bh67_wm60_0_c5 & bh67_wm61_0_c5 & bh67_wm62_0_c5 & bh67_wm63_0_c5 & bh67_wm64_0_c5 & bh67_wm65_0_c5;

   bitheapFinalAdd_bh67_In0_c5 <= "0" & bh67_wm9_5_c5 & bh67_wm10_8_c5 & bh67_wm11_4_c5 & bh67_wm12_7_c5 & bh67_wm13_5_c5 & bh67_wm14_5_c5 & bh67_wm15_4_c5 & bh67_wm16_6_c5 & bh67_wm17_10_c5 & bh67_wm18_10_c5 & bh67_wm19_13_c5 & bh67_wm20_11_c5 & bh67_wm21_16_c5 & bh67_wm22_17_c5 & bh67_wm23_18_c5 & bh67_wm24_19_c5 & bh67_wm25_21_c5 & bh67_wm26_22_c5 & bh67_wm27_20_c5 & bh67_wm28_21_c5 & bh67_wm29_21_c5 & bh67_wm30_22_c5 & bh67_wm31_20_c5 & bh67_wm32_21_c5 & bh67_wm33_21_c5 & bh67_wm34_22_c5 & bh67_wm35_20_c5 & bh67_wm36_20_c5 & bh67_wm37_22_c5 & bh67_wm38_22_c5 & bh67_wm39_19_c5 & bh67_wm40_20_c5;
   bitheapFinalAdd_bh67_In1_c5 <= "0" & "0" & "0" & bh67_wm11_5_c5 & "0" & "0" & "0" & bh67_wm15_5_c5 & "0" & bh67_wm17_11_c5 & "0" & "0" & bh67_wm20_12_c5 & bh67_wm21_17_c5 & bh67_wm22_18_c5 & "0" & bh67_wm24_20_c5 & "0" & bh67_wm26_23_c5 & "0" & bh67_wm28_22_c5 & "0" & bh67_wm30_23_c5 & "0" & bh67_wm32_22_c5 & "0" & bh67_wm34_23_c5 & "0" & bh67_wm36_21_c5 & "0" & bh67_wm38_23_c5 & "0" & bh67_wm40_21_c5;
   bitheapFinalAdd_bh67_Cin_c0 <= '0';

   bitheapFinalAdd_bh67: IntAdder_33_Freq300_uid534
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 Cin => bitheapFinalAdd_bh67_Cin_c0,
                 X => bitheapFinalAdd_bh67_In0_c5,
                 Y => bitheapFinalAdd_bh67_In1_c5,
                 R => bitheapFinalAdd_bh67_Out_c6);
   bitheapResult_bh67_c6 <= bitheapFinalAdd_bh67_Out_c6(31 downto 0) & tmp_bitheapResult_bh67_24_c6;
   RR_c6 <= signed(bitheapResult_bh67_c6(56 downto 24));
R <= std_logic_vector(RR_c6);  
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x24_Freq300_uid539
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid539 is
    port (clk, ce_5, ce_6, ce_7 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid539 is
signal Mfull_c6, Mfull_c7 :  std_logic_vector(40 downto 0);
signal M_c7 :  std_logic_vector(40 downto 0);
signal X_c5, X_c6 :  std_logic_vector(16 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
            if ce_7 = '1' then
               Mfull_c7 <= Mfull_c6;
            end if;
         end if;
      end process;
   Mfull_c6 <= std_logic_vector(unsigned(X_c6) * unsigned(Y)); -- multiplier
   M_c7 <= Mfull_c7(40 downto 0);
   R <= M_c7;
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_12x24_Freq300_uid541
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_12x24_Freq300_uid541 is
    port (clk, ce_5, ce_6, ce_7 : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(35 downto 0)   );
end entity;

architecture arch of DSPBlock_12x24_Freq300_uid541 is
signal Mfull_c6, Mfull_c7 :  std_logic_vector(36 downto 0);
signal M_c7 :  std_logic_vector(35 downto 0);
signal X_c5, X_c6 :  std_logic_vector(11 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
            if ce_7 = '1' then
               Mfull_c7 <= Mfull_c6;
            end if;
         end if;
      end process;
   Mfull_c6 <= std_logic_vector(signed(X_c6) * signed('0' & Y)); -- multiplier
   M_c7 <= Mfull_c7(35 downto 0);
   R <= M_c7;
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_1x1_signed_Freq300_uid543
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_signed_Freq300_uid543 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_signed_Freq300_uid543 is
signal replicated_c4, replicated_c5, replicated_c6 :  std_logic_vector(0 downto 0);
signal prod_c6 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               replicated_c5 <= replicated_c4;
            end if;
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
         end if;
      end process;
   replicated_c4 <= (0 downto 0 => X(0));
   prod_c6 <= Y and replicated_c6;
   R <= prod_c6;
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid545
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid545 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid545 is
   component MultTable_Freq300_uid547 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy548_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid547
      port map ( X => Xtable_c6,
                 Y => Y1_copy548_c6);
   Y1_c6 <= Y1_copy548_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid550
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid550 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid550 is
   component MultTable_Freq300_uid552 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy553_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid552
      port map ( X => Xtable_c6,
                 Y => Y1_copy553_c6);
   Y1_c6 <= Y1_copy553_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid555
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid555 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid555 is
   component MultTable_Freq300_uid557 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy558_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid557
      port map ( X => Xtable_c6,
                 Y => Y1_copy558_c6);
   Y1_c6 <= Y1_copy558_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid560
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid560 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid560 is
   component MultTable_Freq300_uid562 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy563_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid562
      port map ( X => Xtable_c6,
                 Y => Y1_copy563_c6);
   Y1_c6 <= Y1_copy563_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid565
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid565 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid565 is
   component MultTable_Freq300_uid567 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(3 downto 0);
signal Y1_c6 :  std_logic_vector(3 downto 0);
signal Y1_copy568_c6 :  std_logic_vector(3 downto 0);
signal X_c5, X_c6 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid567
      port map ( X => Xtable_c6,
                 Y => Y1_copy568_c6);
   Y1_c6 <= Y1_copy568_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid570
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid570 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid570 is
   component MultTable_Freq300_uid572 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy573_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid572
      port map ( X => Xtable_c6,
                 Y => Y1_copy573_c6);
   Y1_c6 <= Y1_copy573_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid575
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid575 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid575 is
   component MultTable_Freq300_uid577 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy578_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid577
      port map ( X => Xtable_c6,
                 Y => Y1_copy578_c6);
   Y1_c6 <= Y1_copy578_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid580
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid580 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid580 is
   component MultTable_Freq300_uid582 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy583_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid582
      port map ( X => Xtable_c6,
                 Y => Y1_copy583_c6);
   Y1_c6 <= Y1_copy583_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid585
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid585 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid585 is
   component MultTable_Freq300_uid587 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy588_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid587
      port map ( X => Xtable_c6,
                 Y => Y1_copy588_c6);
   Y1_c6 <= Y1_copy588_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid590
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid590 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid590 is
   component MultTable_Freq300_uid592 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy593_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid592
      port map ( X => Xtable_c6,
                 Y => Y1_copy593_c6);
   Y1_c6 <= Y1_copy593_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid595
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid595 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid595 is
   component MultTable_Freq300_uid597 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(3 downto 0);
signal Y1_c6 :  std_logic_vector(3 downto 0);
signal Y1_copy598_c6 :  std_logic_vector(3 downto 0);
signal X_c5, X_c6 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid597
      port map ( X => Xtable_c6,
                 Y => Y1_copy598_c6);
   Y1_c6 <= Y1_copy598_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid600
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid600 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid600 is
   component MultTable_Freq300_uid602 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy603_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid602
      port map ( X => Xtable_c6,
                 Y => Y1_copy603_c6);
   Y1_c6 <= Y1_copy603_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid605
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid605 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid605 is
   component MultTable_Freq300_uid607 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy608_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid607
      port map ( X => Xtable_c6,
                 Y => Y1_copy608_c6);
   Y1_c6 <= Y1_copy608_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid610
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid610 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid610 is
   component MultTable_Freq300_uid612 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy613_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid612
      port map ( X => Xtable_c6,
                 Y => Y1_copy613_c6);
   Y1_c6 <= Y1_copy613_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid615
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid615 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid615 is
   component MultTable_Freq300_uid617 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy618_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid617
      port map ( X => Xtable_c6,
                 Y => Y1_copy618_c6);
   Y1_c6 <= Y1_copy618_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid620
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid620 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid620 is
   component MultTable_Freq300_uid622 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy623_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid622
      port map ( X => Xtable_c6,
                 Y => Y1_copy623_c6);
   Y1_c6 <= Y1_copy623_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid625
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid625 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid625 is
   component MultTable_Freq300_uid627 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(3 downto 0);
signal Y1_c6 :  std_logic_vector(3 downto 0);
signal Y1_copy628_c6 :  std_logic_vector(3 downto 0);
signal X_c5, X_c6 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid627
      port map ( X => Xtable_c6,
                 Y => Y1_copy628_c6);
   Y1_c6 <= Y1_copy628_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid630
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid630 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid630 is
   component MultTable_Freq300_uid632 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy633_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid632
      port map ( X => Xtable_c6,
                 Y => Y1_copy633_c6);
   Y1_c6 <= Y1_copy633_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid635
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid635 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid635 is
   component MultTable_Freq300_uid637 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy638_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid637
      port map ( X => Xtable_c6,
                 Y => Y1_copy638_c6);
   Y1_c6 <= Y1_copy638_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid640
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid640 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid640 is
   component MultTable_Freq300_uid642 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy643_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid642
      port map ( X => Xtable_c6,
                 Y => Y1_copy643_c6);
   Y1_c6 <= Y1_copy643_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid645
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid645 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid645 is
   component MultTable_Freq300_uid647 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy648_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid647
      port map ( X => Xtable_c6,
                 Y => Y1_copy648_c6);
   Y1_c6 <= Y1_copy648_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid650
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid650 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid650 is
   component MultTable_Freq300_uid652 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy653_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid652
      port map ( X => Xtable_c6,
                 Y => Y1_copy653_c6);
   Y1_c6 <= Y1_copy653_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid655
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid655 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid655 is
   component MultTable_Freq300_uid657 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(3 downto 0);
signal Y1_c6 :  std_logic_vector(3 downto 0);
signal Y1_copy658_c6 :  std_logic_vector(3 downto 0);
signal X_c5, X_c6 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid657
      port map ( X => Xtable_c6,
                 Y => Y1_copy658_c6);
   Y1_c6 <= Y1_copy658_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid660
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid660 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid660 is
   component MultTable_Freq300_uid662 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy663_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid662
      port map ( X => Xtable_c6,
                 Y => Y1_copy663_c6);
   Y1_c6 <= Y1_copy663_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid665
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid665 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid665 is
   component MultTable_Freq300_uid667 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy668_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid667
      port map ( X => Xtable_c6,
                 Y => Y1_copy668_c6);
   Y1_c6 <= Y1_copy668_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid670
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid670 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid670 is
   component MultTable_Freq300_uid672 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy673_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid672
      port map ( X => Xtable_c6,
                 Y => Y1_copy673_c6);
   Y1_c6 <= Y1_copy673_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid675
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid675 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid675 is
   component MultTable_Freq300_uid677 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy678_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid677
      port map ( X => Xtable_c6,
                 Y => Y1_copy678_c6);
   Y1_c6 <= Y1_copy678_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid680
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid680 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid680 is
   component MultTable_Freq300_uid682 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy683_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid682
      port map ( X => Xtable_c6,
                 Y => Y1_copy683_c6);
   Y1_c6 <= Y1_copy683_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--             IntMultiplierLUT_4_signedx1_signed_Freq300_uid685
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4_signedx1_signed_Freq300_uid685 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4_signedx1_signed_Freq300_uid685 is
   component MultTable_Freq300_uid687 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy688_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid687
      port map ( X => Xtable_c6,
                 Y => Y1_copy688_c6);
   Y1_c6 <= Y1_copy688_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid690
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid690 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid690 is
   component MultTable_Freq300_uid692 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy693_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid692
      port map ( X => Xtable_c6,
                 Y => Y1_copy693_c6);
   Y1_c6 <= Y1_copy693_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_4x1_signed_Freq300_uid695
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_signed_Freq300_uid695 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_signed_Freq300_uid695 is
   component MultTable_Freq300_uid697 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy698_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(3 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid697
      port map ( X => Xtable_c6,
                 Y => Y1_copy698_c6);
   Y1_c6 <= Y1_copy698_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_3_signedx2_Freq300_uid700
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3_signedx2_Freq300_uid700 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3_signedx2_Freq300_uid700 is
   component MultTable_Freq300_uid702 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy703_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid702
      port map ( X => Xtable_c6,
                 Y => Y1_copy703_c6);
   Y1_c6 <= Y1_copy703_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid705
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid705 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid705 is
   component MultTable_Freq300_uid707 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy708_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid707
      port map ( X => Xtable_c6,
                 Y => Y1_copy708_c6);
   Y1_c6 <= Y1_copy708_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid710
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid710 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid710 is
   component MultTable_Freq300_uid712 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy713_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid712
      port map ( X => Xtable_c6,
                 Y => Y1_copy713_c6);
   Y1_c6 <= Y1_copy713_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid715
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid715 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid715 is
   component MultTable_Freq300_uid717 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy718_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid717
      port map ( X => Xtable_c6,
                 Y => Y1_copy718_c6);
   Y1_c6 <= Y1_copy718_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_3_signedx2_Freq300_uid720
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3_signedx2_Freq300_uid720 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3_signedx2_Freq300_uid720 is
   component MultTable_Freq300_uid722 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy723_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid722
      port map ( X => Xtable_c6,
                 Y => Y1_copy723_c6);
   Y1_c6 <= Y1_copy723_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid725
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid725 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid725 is
   component MultTable_Freq300_uid727 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy728_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid727
      port map ( X => Xtable_c6,
                 Y => Y1_copy728_c6);
   Y1_c6 <= Y1_copy728_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid730
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid730 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid730 is
   component MultTable_Freq300_uid732 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy733_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid732
      port map ( X => Xtable_c6,
                 Y => Y1_copy733_c6);
   Y1_c6 <= Y1_copy733_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid735
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid735 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid735 is
   component MultTable_Freq300_uid737 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy738_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid737
      port map ( X => Xtable_c6,
                 Y => Y1_copy738_c6);
   Y1_c6 <= Y1_copy738_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_3_signedx2_Freq300_uid740
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3_signedx2_Freq300_uid740 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3_signedx2_Freq300_uid740 is
   component MultTable_Freq300_uid742 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy743_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid742
      port map ( X => Xtable_c6,
                 Y => Y1_copy743_c6);
   Y1_c6 <= Y1_copy743_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid745
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid745 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid745 is
   component MultTable_Freq300_uid747 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy748_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid747
      port map ( X => Xtable_c6,
                 Y => Y1_copy748_c6);
   Y1_c6 <= Y1_copy748_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid750
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid750 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid750 is
   component MultTable_Freq300_uid752 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy753_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid752
      port map ( X => Xtable_c6,
                 Y => Y1_copy753_c6);
   Y1_c6 <= Y1_copy753_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid755
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid755 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid755 is
   component MultTable_Freq300_uid757 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy758_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid757
      port map ( X => Xtable_c6,
                 Y => Y1_copy758_c6);
   Y1_c6 <= Y1_copy758_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                 IntMultiplierLUT_3_signedx2_Freq300_uid760
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3_signedx2_Freq300_uid760 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3_signedx2_Freq300_uid760 is
   component MultTable_Freq300_uid762 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy763_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid762
      port map ( X => Xtable_c6,
                 Y => Y1_copy763_c6);
   Y1_c6 <= Y1_copy763_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid765
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid765 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid765 is
   component MultTable_Freq300_uid767 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy768_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid767
      port map ( X => Xtable_c6,
                 Y => Y1_copy768_c6);
   Y1_c6 <= Y1_copy768_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid770
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid770 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid770 is
   component MultTable_Freq300_uid772 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy773_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid772
      port map ( X => Xtable_c6,
                 Y => Y1_copy773_c6);
   Y1_c6 <= Y1_copy773_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid775
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid775 is
    port (clk, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid775 is
   component MultTable_Freq300_uid777 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c6 :  std_logic_vector(4 downto 0);
signal Y1_c6 :  std_logic_vector(4 downto 0);
signal Y1_copy778_c6 :  std_logic_vector(4 downto 0);
signal X_c5, X_c6 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               X_c5 <= X;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
            end if;
         end if;
      end process;
Xtable_c6 <= Y & X_c6;
   R <= Y1_c6;
   TableMult: MultTable_Freq300_uid777
      port map ( X => Xtable_c6,
                 Y => Y1_copy778_c6);
   Y1_c6 <= Y1_copy778_c6; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_45_Freq300_uid1105
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 8 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_45_Freq300_uid1105 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
          X : in  std_logic_vector(44 downto 0);
          Y : in  std_logic_vector(44 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(44 downto 0)   );
end entity;

architecture arch of IntAdder_45_Freq300_uid1105 is
signal Rtmp_c8 :  std_logic_vector(44 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
         end if;
      end process;
   Rtmp_c8 <= X + Y + Cin_c8;
   R <= Rtmp_c8;
end architecture;

--------------------------------------------------------------------------------
--    FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid536
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Matei Istoan, 2012-2014, 2024
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y A
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid536 is
    port (clk, ce_5, ce_6, ce_7, ce_8 : in std_logic;
          X : in  std_logic_vector(28 downto 0);
          Y : in  std_logic_vector(32 downto 0);
          A : in  std_logic_vector(39 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid536 is
   component DSPBlock_17x24_Freq300_uid539 is
      port ( clk, ce_5, ce_6, ce_7 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_12x24_Freq300_uid541 is
      port ( clk, ce_5, ce_6, ce_7 : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(35 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_signed_Freq300_uid543 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid545 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid550 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid555 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid560 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid565 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid570 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid575 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid580 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid585 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid590 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid595 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid600 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid605 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid610 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid615 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid620 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid625 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid630 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid635 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid640 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid645 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid650 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid655 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid660 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid665 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid670 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid675 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid680 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4_signedx1_signed_Freq300_uid685 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid690 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_signed_Freq300_uid695 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3_signedx2_Freq300_uid700 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid705 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid710 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid715 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3_signedx2_Freq300_uid720 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid725 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid730 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid735 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3_signedx2_Freq300_uid740 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid745 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid750 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid755 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3_signedx2_Freq300_uid760 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid765 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid770 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid775 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid781 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid789 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid797 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid813 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq300_uid839 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_45_Freq300_uid1105 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
             X : in  std_logic_vector(44 downto 0);
             Y : in  std_logic_vector(44 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(44 downto 0)   );
   end component;

signal XX_c4 :  signed(0+28 downto 0);
signal YY_c6 :  signed(-9+41 downto 0);
signal AA_c4 :  signed(-2+41 downto 0);
signal tile_0_X_c4 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c6 :  std_logic_vector(23 downto 0);
signal tile_0_output_c7 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c7 :  unsigned(40-0 downto 0);
signal bh537_wm69_0_c7, bh537_wm69_0_c8 :  std_logic;
signal bh537_wm68_0_c7, bh537_wm68_0_c8 :  std_logic;
signal bh537_wm67_0_c7, bh537_wm67_0_c8 :  std_logic;
signal bh537_wm66_0_c7, bh537_wm66_0_c8 :  std_logic;
signal bh537_wm65_0_c7, bh537_wm65_0_c8 :  std_logic;
signal bh537_wm64_0_c7, bh537_wm64_0_c8 :  std_logic;
signal bh537_wm63_0_c7, bh537_wm63_0_c8 :  std_logic;
signal bh537_wm62_0_c7, bh537_wm62_0_c8 :  std_logic;
signal bh537_wm61_0_c7, bh537_wm61_0_c8 :  std_logic;
signal bh537_wm60_0_c7, bh537_wm60_0_c8 :  std_logic;
signal bh537_wm59_0_c7, bh537_wm59_0_c8 :  std_logic;
signal bh537_wm58_0_c7, bh537_wm58_0_c8 :  std_logic;
signal bh537_wm57_0_c7, bh537_wm57_0_c8 :  std_logic;
signal bh537_wm56_0_c7, bh537_wm56_0_c8 :  std_logic;
signal bh537_wm55_0_c7, bh537_wm55_0_c8 :  std_logic;
signal bh537_wm54_0_c7, bh537_wm54_0_c8 :  std_logic;
signal bh537_wm53_0_c7, bh537_wm53_0_c8 :  std_logic;
signal bh537_wm52_0_c7 :  std_logic;
signal bh537_wm51_0_c7 :  std_logic;
signal bh537_wm50_0_c7 :  std_logic;
signal bh537_wm49_0_c7 :  std_logic;
signal bh537_wm48_0_c7 :  std_logic;
signal bh537_wm47_0_c7 :  std_logic;
signal bh537_wm46_0_c7 :  std_logic;
signal bh537_wm45_0_c7 :  std_logic;
signal bh537_wm44_0_c7 :  std_logic;
signal bh537_wm43_0_c7 :  std_logic;
signal bh537_wm42_0_c7 :  std_logic;
signal bh537_wm41_0_c7 :  std_logic;
signal bh537_wm40_0_c7 :  std_logic;
signal bh537_wm39_0_c7 :  std_logic;
signal bh537_wm38_0_c7 :  std_logic;
signal bh537_wm37_0_c7 :  std_logic;
signal bh537_wm36_0_c7 :  std_logic;
signal bh537_wm35_0_c7 :  std_logic;
signal bh537_wm34_0_c7 :  std_logic;
signal bh537_wm33_0_c7 :  std_logic;
signal bh537_wm32_0_c7 :  std_logic;
signal bh537_wm31_0_c7 :  std_logic;
signal bh537_wm30_0_c7 :  std_logic;
signal bh537_wm29_0_c7 :  std_logic;
signal tile_1_X_c4 :  std_logic_vector(11 downto 0);
signal tile_1_Y_c6 :  std_logic_vector(23 downto 0);
signal tile_1_output_c7 :  std_logic_vector(35 downto 0);
signal tile_1_filtered_output_c7 :  signed(35-0 downto 0);
signal bh537_wm52_1_c7 :  std_logic;
signal bh537_wm51_1_c7 :  std_logic;
signal bh537_wm50_1_c7 :  std_logic;
signal bh537_wm49_1_c7 :  std_logic;
signal bh537_wm48_1_c7 :  std_logic;
signal bh537_wm47_1_c7 :  std_logic;
signal bh537_wm46_1_c7 :  std_logic;
signal bh537_wm45_1_c7 :  std_logic;
signal bh537_wm44_1_c7 :  std_logic;
signal bh537_wm43_1_c7 :  std_logic;
signal bh537_wm42_1_c7 :  std_logic;
signal bh537_wm41_1_c7 :  std_logic;
signal bh537_wm40_1_c7 :  std_logic;
signal bh537_wm39_1_c7 :  std_logic;
signal bh537_wm38_1_c7 :  std_logic;
signal bh537_wm37_1_c7 :  std_logic;
signal bh537_wm36_1_c7 :  std_logic;
signal bh537_wm35_1_c7 :  std_logic;
signal bh537_wm34_1_c7 :  std_logic;
signal bh537_wm33_1_c7 :  std_logic;
signal bh537_wm32_1_c7 :  std_logic;
signal bh537_wm31_1_c7 :  std_logic;
signal bh537_wm30_1_c7 :  std_logic;
signal bh537_wm29_1_c7 :  std_logic;
signal bh537_wm28_0_c7 :  std_logic;
signal bh537_wm27_0_c7 :  std_logic;
signal bh537_wm26_0_c7 :  std_logic;
signal bh537_wm25_0_c7 :  std_logic;
signal bh537_wm24_0_c7 :  std_logic;
signal bh537_wm23_0_c7 :  std_logic;
signal bh537_wm22_0_c7 :  std_logic;
signal bh537_wm21_0_c7 :  std_logic;
signal bh537_wm20_0_c7 :  std_logic;
signal bh537_wm19_0_c7 :  std_logic;
signal bh537_wm18_0_c7 :  std_logic;
signal bh537_wm17_0_c7 :  std_logic;
signal tile_2_X_c4 :  std_logic_vector(0 downto 0);
signal tile_2_Y_c6 :  std_logic_vector(0 downto 0);
signal tile_2_output_c6 :  std_logic_vector(0 downto 0);
signal tile_2_filtered_output_c6 :  signed(0-0 downto 0);
signal bh537_wm21_1_c6, bh537_wm21_1_c7 :  std_logic;
signal tile_3_X_c4 :  std_logic_vector(3 downto 0);
signal tile_3_Y_c6 :  std_logic_vector(0 downto 0);
signal tile_3_output_c6 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm25_1_c6 :  std_logic;
signal bh537_wm24_1_c6 :  std_logic;
signal bh537_wm23_1_c6 :  std_logic;
signal bh537_wm22_1_c6 :  std_logic;
signal bh537_wm21_2_c6, bh537_wm21_2_c7 :  std_logic;
signal tile_4_X_c4 :  std_logic_vector(3 downto 0);
signal tile_4_Y_c6 :  std_logic_vector(0 downto 0);
signal tile_4_output_c6 :  std_logic_vector(4 downto 0);
signal tile_4_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm29_2_c6, bh537_wm29_2_c7 :  std_logic;
signal bh537_wm28_1_c6, bh537_wm28_1_c7 :  std_logic;
signal bh537_wm27_1_c6 :  std_logic;
signal bh537_wm26_1_c6 :  std_logic;
signal bh537_wm25_2_c6 :  std_logic;
signal tile_5_X_c4 :  std_logic_vector(3 downto 0);
signal tile_5_Y_c6 :  std_logic_vector(0 downto 0);
signal tile_5_output_c6 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm33_2_c6, bh537_wm33_2_c7 :  std_logic;
signal bh537_wm32_2_c6, bh537_wm32_2_c7 :  std_logic;
signal bh537_wm31_2_c6, bh537_wm31_2_c7 :  std_logic;
signal bh537_wm30_2_c6, bh537_wm30_2_c7 :  std_logic;
signal bh537_wm29_3_c6, bh537_wm29_3_c7 :  std_logic;
signal tile_6_X_c4 :  std_logic_vector(3 downto 0);
signal tile_6_Y_c6 :  std_logic_vector(0 downto 0);
signal tile_6_output_c6 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm37_2_c6, bh537_wm37_2_c7 :  std_logic;
signal bh537_wm36_2_c6, bh537_wm36_2_c7 :  std_logic;
signal bh537_wm35_2_c6, bh537_wm35_2_c7 :  std_logic;
signal bh537_wm34_2_c6, bh537_wm34_2_c7 :  std_logic;
signal bh537_wm33_3_c6, bh537_wm33_3_c7 :  std_logic;
signal tile_7_X_c4 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_7_output_c6 :  std_logic_vector(3 downto 0);
signal tile_7_filtered_output_c6 :  unsigned(3-0 downto 0);
signal bh537_wm24_2_c6 :  std_logic;
signal bh537_wm23_2_c6 :  std_logic;
signal bh537_wm22_2_c6 :  std_logic;
signal bh537_wm21_3_c6, bh537_wm21_3_c7 :  std_logic;
signal tile_8_X_c4 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_8_output_c6 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm27_2_c6 :  std_logic;
signal bh537_wm26_2_c6 :  std_logic;
signal bh537_wm25_3_c6 :  std_logic;
signal bh537_wm24_3_c6 :  std_logic;
signal bh537_wm23_3_c6 :  std_logic;
signal tile_9_X_c4 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_9_output_c6 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm30_3_c6, bh537_wm30_3_c7 :  std_logic;
signal bh537_wm29_4_c6, bh537_wm29_4_c7 :  std_logic;
signal bh537_wm28_2_c6, bh537_wm28_2_c7 :  std_logic;
signal bh537_wm27_3_c6 :  std_logic;
signal bh537_wm26_3_c6 :  std_logic;
signal tile_10_X_c4 :  std_logic_vector(2 downto 0);
signal tile_10_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_10_output_c6 :  std_logic_vector(4 downto 0);
signal tile_10_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm33_4_c6, bh537_wm33_4_c7 :  std_logic;
signal bh537_wm32_3_c6, bh537_wm32_3_c7 :  std_logic;
signal bh537_wm31_3_c6, bh537_wm31_3_c7 :  std_logic;
signal bh537_wm30_4_c6, bh537_wm30_4_c7 :  std_logic;
signal bh537_wm29_5_c6, bh537_wm29_5_c7 :  std_logic;
signal tile_11_X_c4 :  std_logic_vector(2 downto 0);
signal tile_11_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_11_output_c6 :  std_logic_vector(4 downto 0);
signal tile_11_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm36_3_c6, bh537_wm36_3_c7 :  std_logic;
signal bh537_wm35_3_c6, bh537_wm35_3_c7 :  std_logic;
signal bh537_wm34_3_c6, bh537_wm34_3_c7 :  std_logic;
signal bh537_wm33_5_c6, bh537_wm33_5_c7 :  std_logic;
signal bh537_wm32_4_c6, bh537_wm32_4_c7 :  std_logic;
signal tile_12_X_c4 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_12_output_c6 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm39_2_c6, bh537_wm39_2_c7 :  std_logic;
signal bh537_wm38_2_c6 :  std_logic;
signal bh537_wm37_3_c6, bh537_wm37_3_c7 :  std_logic;
signal bh537_wm36_4_c6, bh537_wm36_4_c7 :  std_logic;
signal bh537_wm35_4_c6, bh537_wm35_4_c7 :  std_logic;
signal tile_13_X_c4 :  std_logic_vector(1 downto 0);
signal tile_13_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_13_output_c6 :  std_logic_vector(3 downto 0);
signal tile_13_filtered_output_c6 :  unsigned(3-0 downto 0);
signal bh537_wm26_4_c6 :  std_logic;
signal bh537_wm25_4_c6 :  std_logic;
signal bh537_wm24_4_c6 :  std_logic;
signal bh537_wm23_4_c6 :  std_logic;
signal tile_14_X_c4 :  std_logic_vector(2 downto 0);
signal tile_14_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_14_output_c6 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm29_6_c6 :  std_logic;
signal bh537_wm28_3_c6, bh537_wm28_3_c7 :  std_logic;
signal bh537_wm27_4_c6 :  std_logic;
signal bh537_wm26_5_c6 :  std_logic;
signal bh537_wm25_5_c6 :  std_logic;
signal tile_15_X_c4 :  std_logic_vector(2 downto 0);
signal tile_15_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_15_output_c6 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm32_5_c6, bh537_wm32_5_c7 :  std_logic;
signal bh537_wm31_4_c6, bh537_wm31_4_c7 :  std_logic;
signal bh537_wm30_5_c6, bh537_wm30_5_c7 :  std_logic;
signal bh537_wm29_7_c6 :  std_logic;
signal bh537_wm28_4_c6, bh537_wm28_4_c7 :  std_logic;
signal tile_16_X_c4 :  std_logic_vector(2 downto 0);
signal tile_16_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_16_output_c6 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm35_5_c6, bh537_wm35_5_c7 :  std_logic;
signal bh537_wm34_4_c6, bh537_wm34_4_c7 :  std_logic;
signal bh537_wm33_6_c6, bh537_wm33_6_c7 :  std_logic;
signal bh537_wm32_6_c6 :  std_logic;
signal bh537_wm31_5_c6, bh537_wm31_5_c7 :  std_logic;
signal tile_17_X_c4 :  std_logic_vector(2 downto 0);
signal tile_17_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_17_output_c6 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm38_3_c6 :  std_logic;
signal bh537_wm37_4_c6, bh537_wm37_4_c7 :  std_logic;
signal bh537_wm36_5_c6, bh537_wm36_5_c7 :  std_logic;
signal bh537_wm35_6_c6, bh537_wm35_6_c7 :  std_logic;
signal bh537_wm34_5_c6, bh537_wm34_5_c7 :  std_logic;
signal tile_18_X_c4 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_18_output_c6 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm41_2_c6, bh537_wm41_2_c7 :  std_logic;
signal bh537_wm40_2_c6, bh537_wm40_2_c7 :  std_logic;
signal bh537_wm39_3_c6, bh537_wm39_3_c7 :  std_logic;
signal bh537_wm38_4_c6 :  std_logic;
signal bh537_wm37_5_c6, bh537_wm37_5_c7 :  std_logic;
signal tile_19_X_c4 :  std_logic_vector(1 downto 0);
signal tile_19_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_19_output_c6 :  std_logic_vector(3 downto 0);
signal tile_19_filtered_output_c6 :  unsigned(3-0 downto 0);
signal bh537_wm28_5_c6, bh537_wm28_5_c7 :  std_logic;
signal bh537_wm27_5_c6 :  std_logic;
signal bh537_wm26_6_c6 :  std_logic;
signal bh537_wm25_6_c6 :  std_logic;
signal tile_20_X_c4 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_20_output_c6 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm31_6_c6 :  std_logic;
signal bh537_wm30_6_c6 :  std_logic;
signal bh537_wm29_8_c6 :  std_logic;
signal bh537_wm28_6_c6 :  std_logic;
signal bh537_wm27_6_c6 :  std_logic;
signal tile_21_X_c4 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_21_output_c6 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm34_6_c6, bh537_wm34_6_c7 :  std_logic;
signal bh537_wm33_7_c6, bh537_wm33_7_c7 :  std_logic;
signal bh537_wm32_7_c6 :  std_logic;
signal bh537_wm31_7_c6 :  std_logic;
signal bh537_wm30_7_c6 :  std_logic;
signal tile_22_X_c4 :  std_logic_vector(2 downto 0);
signal tile_22_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_22_output_c6 :  std_logic_vector(4 downto 0);
signal tile_22_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm37_6_c6 :  std_logic;
signal bh537_wm36_6_c6, bh537_wm36_6_c7 :  std_logic;
signal bh537_wm35_7_c6 :  std_logic;
signal bh537_wm34_7_c6 :  std_logic;
signal bh537_wm33_8_c6, bh537_wm33_8_c7 :  std_logic;
signal tile_23_X_c4 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_23_output_c6 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm40_3_c6, bh537_wm40_3_c7 :  std_logic;
signal bh537_wm39_4_c6, bh537_wm39_4_c7 :  std_logic;
signal bh537_wm38_5_c6 :  std_logic;
signal bh537_wm37_7_c6 :  std_logic;
signal bh537_wm36_7_c6 :  std_logic;
signal tile_24_X_c4 :  std_logic_vector(2 downto 0);
signal tile_24_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_24_output_c6 :  std_logic_vector(4 downto 0);
signal tile_24_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm43_2_c6, bh537_wm43_2_c7 :  std_logic;
signal bh537_wm42_2_c6, bh537_wm42_2_c7 :  std_logic;
signal bh537_wm41_3_c6, bh537_wm41_3_c7 :  std_logic;
signal bh537_wm40_4_c6, bh537_wm40_4_c7 :  std_logic;
signal bh537_wm39_5_c6, bh537_wm39_5_c7 :  std_logic;
signal tile_25_X_c4 :  std_logic_vector(1 downto 0);
signal tile_25_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_25_output_c6 :  std_logic_vector(3 downto 0);
signal tile_25_filtered_output_c6 :  unsigned(3-0 downto 0);
signal bh537_wm30_8_c6 :  std_logic;
signal bh537_wm29_9_c6 :  std_logic;
signal bh537_wm28_7_c6 :  std_logic;
signal bh537_wm27_7_c6 :  std_logic;
signal tile_26_X_c4 :  std_logic_vector(2 downto 0);
signal tile_26_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_26_output_c6 :  std_logic_vector(4 downto 0);
signal tile_26_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm33_9_c6, bh537_wm33_9_c7 :  std_logic;
signal bh537_wm32_8_c6 :  std_logic;
signal bh537_wm31_8_c6 :  std_logic;
signal bh537_wm30_9_c6 :  std_logic;
signal bh537_wm29_10_c6 :  std_logic;
signal tile_27_X_c4 :  std_logic_vector(2 downto 0);
signal tile_27_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_27_output_c6 :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm36_8_c6 :  std_logic;
signal bh537_wm35_8_c6 :  std_logic;
signal bh537_wm34_8_c6 :  std_logic;
signal bh537_wm33_10_c6, bh537_wm33_10_c7 :  std_logic;
signal bh537_wm32_9_c6 :  std_logic;
signal tile_28_X_c4 :  std_logic_vector(2 downto 0);
signal tile_28_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_28_output_c6 :  std_logic_vector(4 downto 0);
signal tile_28_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm39_6_c6 :  std_logic;
signal bh537_wm38_6_c6 :  std_logic;
signal bh537_wm37_8_c6 :  std_logic;
signal bh537_wm36_9_c6 :  std_logic;
signal bh537_wm35_9_c6 :  std_logic;
signal tile_29_X_c4 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_29_output_c6 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm42_3_c6, bh537_wm42_3_c7 :  std_logic;
signal bh537_wm41_4_c6, bh537_wm41_4_c7 :  std_logic;
signal bh537_wm40_5_c6, bh537_wm40_5_c7 :  std_logic;
signal bh537_wm39_7_c6 :  std_logic;
signal bh537_wm38_7_c6 :  std_logic;
signal tile_30_X_c4 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_30_output_c6 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm45_2_c6, bh537_wm45_2_c7 :  std_logic;
signal bh537_wm44_2_c6, bh537_wm44_2_c7 :  std_logic;
signal bh537_wm43_3_c6, bh537_wm43_3_c7 :  std_logic;
signal bh537_wm42_4_c6, bh537_wm42_4_c7 :  std_logic;
signal bh537_wm41_5_c6, bh537_wm41_5_c7 :  std_logic;
signal tile_31_X_c4 :  std_logic_vector(3 downto 0);
signal tile_31_Y_c6 :  std_logic_vector(0 downto 0);
signal tile_31_output_c6 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm12_0_c6 :  std_logic;
signal bh537_wm11_0_c6 :  std_logic;
signal bh537_wm10_0_c6 :  std_logic;
signal bh537_wm9_0_c6 :  std_logic;
signal bh537_wm8_0_c6 :  std_logic;
signal tile_32_X_c4 :  std_logic_vector(3 downto 0);
signal tile_32_Y_c6 :  std_logic_vector(0 downto 0);
signal tile_32_output_c6 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm16_0_c6 :  std_logic;
signal bh537_wm15_0_c6 :  std_logic;
signal bh537_wm14_0_c6 :  std_logic;
signal bh537_wm13_0_c6 :  std_logic;
signal bh537_wm12_1_c6 :  std_logic;
signal tile_33_X_c4 :  std_logic_vector(3 downto 0);
signal tile_33_Y_c6 :  std_logic_vector(0 downto 0);
signal tile_33_output_c6 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm20_1_c6, bh537_wm20_1_c7 :  std_logic;
signal bh537_wm19_1_c6, bh537_wm19_1_c7 :  std_logic;
signal bh537_wm18_1_c6 :  std_logic;
signal bh537_wm17_1_c6, bh537_wm17_1_c7 :  std_logic;
signal bh537_wm16_1_c6 :  std_logic;
signal tile_34_X_c4 :  std_logic_vector(2 downto 0);
signal tile_34_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_34_output_c6 :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm13_1_c6 :  std_logic;
signal bh537_wm12_2_c6 :  std_logic;
signal bh537_wm11_1_c6 :  std_logic;
signal bh537_wm10_1_c6 :  std_logic;
signal bh537_wm9_1_c6 :  std_logic;
signal tile_35_X_c4 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_35_output_c6 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm16_2_c6 :  std_logic;
signal bh537_wm15_1_c6 :  std_logic;
signal bh537_wm14_1_c6 :  std_logic;
signal bh537_wm13_2_c6 :  std_logic;
signal bh537_wm12_3_c6 :  std_logic;
signal tile_36_X_c4 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_36_output_c6 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm19_2_c6, bh537_wm19_2_c7 :  std_logic;
signal bh537_wm18_2_c6 :  std_logic;
signal bh537_wm17_2_c6, bh537_wm17_2_c7 :  std_logic;
signal bh537_wm16_3_c6 :  std_logic;
signal bh537_wm15_2_c6 :  std_logic;
signal tile_37_X_c4 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_37_output_c6 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm22_3_c6 :  std_logic;
signal bh537_wm21_4_c6, bh537_wm21_4_c7 :  std_logic;
signal bh537_wm20_2_c6, bh537_wm20_2_c7 :  std_logic;
signal bh537_wm19_3_c6, bh537_wm19_3_c7 :  std_logic;
signal bh537_wm18_3_c6 :  std_logic;
signal tile_38_X_c4 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_38_output_c6 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm15_3_c6 :  std_logic;
signal bh537_wm14_2_c6 :  std_logic;
signal bh537_wm13_3_c6 :  std_logic;
signal bh537_wm12_4_c6 :  std_logic;
signal bh537_wm11_2_c6 :  std_logic;
signal tile_39_X_c4 :  std_logic_vector(2 downto 0);
signal tile_39_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_39_output_c6 :  std_logic_vector(4 downto 0);
signal tile_39_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm18_4_c6 :  std_logic;
signal bh537_wm17_3_c6, bh537_wm17_3_c7 :  std_logic;
signal bh537_wm16_4_c6 :  std_logic;
signal bh537_wm15_4_c6 :  std_logic;
signal bh537_wm14_3_c6 :  std_logic;
signal tile_40_X_c4 :  std_logic_vector(2 downto 0);
signal tile_40_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_40_output_c6 :  std_logic_vector(4 downto 0);
signal tile_40_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm21_5_c6, bh537_wm21_5_c7 :  std_logic;
signal bh537_wm20_3_c6, bh537_wm20_3_c7 :  std_logic;
signal bh537_wm19_4_c6, bh537_wm19_4_c7 :  std_logic;
signal bh537_wm18_5_c6 :  std_logic;
signal bh537_wm17_4_c6, bh537_wm17_4_c7 :  std_logic;
signal tile_41_X_c4 :  std_logic_vector(2 downto 0);
signal tile_41_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_41_output_c6 :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm24_5_c6 :  std_logic;
signal bh537_wm23_5_c6 :  std_logic;
signal bh537_wm22_4_c6 :  std_logic;
signal bh537_wm21_6_c6 :  std_logic;
signal bh537_wm20_4_c6, bh537_wm20_4_c7 :  std_logic;
signal tile_42_X_c4 :  std_logic_vector(2 downto 0);
signal tile_42_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_42_output_c6 :  std_logic_vector(4 downto 0);
signal tile_42_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm17_5_c6, bh537_wm17_5_c7 :  std_logic;
signal bh537_wm16_5_c6 :  std_logic;
signal bh537_wm15_5_c6 :  std_logic;
signal bh537_wm14_4_c6 :  std_logic;
signal bh537_wm13_4_c6 :  std_logic;
signal tile_43_X_c4 :  std_logic_vector(2 downto 0);
signal tile_43_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_43_output_c6 :  std_logic_vector(4 downto 0);
signal tile_43_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm20_5_c6, bh537_wm20_5_c7 :  std_logic;
signal bh537_wm19_5_c6, bh537_wm19_5_c7 :  std_logic;
signal bh537_wm18_6_c6 :  std_logic;
signal bh537_wm17_6_c6 :  std_logic;
signal bh537_wm16_6_c6 :  std_logic;
signal tile_44_X_c4 :  std_logic_vector(2 downto 0);
signal tile_44_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_44_output_c6 :  std_logic_vector(4 downto 0);
signal tile_44_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm23_6_c6 :  std_logic;
signal bh537_wm22_5_c6 :  std_logic;
signal bh537_wm21_7_c6 :  std_logic;
signal bh537_wm20_6_c6 :  std_logic;
signal bh537_wm19_6_c6 :  std_logic;
signal tile_45_X_c4 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_45_output_c6 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm26_7_c6 :  std_logic;
signal bh537_wm25_7_c6 :  std_logic;
signal bh537_wm24_6_c6 :  std_logic;
signal bh537_wm23_7_c6 :  std_logic;
signal bh537_wm22_6_c6 :  std_logic;
signal tile_46_X_c4 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_46_output_c6 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c6 :  signed(4-0 downto 0);
signal bh537_wm19_7_c6 :  std_logic;
signal bh537_wm18_7_c6 :  std_logic;
signal bh537_wm17_7_c6 :  std_logic;
signal bh537_wm16_7_c6 :  std_logic;
signal bh537_wm15_6_c6 :  std_logic;
signal tile_47_X_c4 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_47_output_c6 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm22_7_c6 :  std_logic;
signal bh537_wm21_8_c6 :  std_logic;
signal bh537_wm20_7_c6 :  std_logic;
signal bh537_wm19_8_c6 :  std_logic;
signal bh537_wm18_8_c6 :  std_logic;
signal tile_48_X_c4 :  std_logic_vector(2 downto 0);
signal tile_48_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_48_output_c6 :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm25_8_c6 :  std_logic;
signal bh537_wm24_7_c6 :  std_logic;
signal bh537_wm23_8_c6 :  std_logic;
signal bh537_wm22_8_c6 :  std_logic;
signal bh537_wm21_9_c6 :  std_logic;
signal tile_49_X_c4 :  std_logic_vector(2 downto 0);
signal tile_49_Y_c6 :  std_logic_vector(1 downto 0);
signal tile_49_output_c6 :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output_c6 :  unsigned(4-0 downto 0);
signal bh537_wm28_8_c6 :  std_logic;
signal bh537_wm27_8_c6 :  std_logic;
signal bh537_wm26_8_c6 :  std_logic;
signal bh537_wm25_9_c6 :  std_logic;
signal bh537_wm24_8_c6 :  std_logic;
signal bh537_wm41_6_c4, bh537_wm41_6_c5, bh537_wm41_6_c6, bh537_wm41_6_c7 :  std_logic;
signal bh537_wm40_6_c4, bh537_wm40_6_c5, bh537_wm40_6_c6, bh537_wm40_6_c7 :  std_logic;
signal bh537_wm39_8_c4, bh537_wm39_8_c5, bh537_wm39_8_c6 :  std_logic;
signal bh537_wm38_8_c4, bh537_wm38_8_c5, bh537_wm38_8_c6, bh537_wm38_8_c7 :  std_logic;
signal bh537_wm37_9_c4, bh537_wm37_9_c5, bh537_wm37_9_c6 :  std_logic;
signal bh537_wm36_10_c4, bh537_wm36_10_c5, bh537_wm36_10_c6 :  std_logic;
signal bh537_wm35_10_c4, bh537_wm35_10_c5, bh537_wm35_10_c6 :  std_logic;
signal bh537_wm34_9_c4, bh537_wm34_9_c5, bh537_wm34_9_c6 :  std_logic;
signal bh537_wm33_11_c4, bh537_wm33_11_c5, bh537_wm33_11_c6, bh537_wm33_11_c7 :  std_logic;
signal bh537_wm32_10_c4, bh537_wm32_10_c5, bh537_wm32_10_c6 :  std_logic;
signal bh537_wm31_9_c4, bh537_wm31_9_c5, bh537_wm31_9_c6 :  std_logic;
signal bh537_wm30_10_c4, bh537_wm30_10_c5, bh537_wm30_10_c6 :  std_logic;
signal bh537_wm29_11_c4, bh537_wm29_11_c5, bh537_wm29_11_c6 :  std_logic;
signal bh537_wm28_9_c4, bh537_wm28_9_c5, bh537_wm28_9_c6 :  std_logic;
signal bh537_wm27_9_c4, bh537_wm27_9_c5, bh537_wm27_9_c6 :  std_logic;
signal bh537_wm26_9_c4, bh537_wm26_9_c5, bh537_wm26_9_c6 :  std_logic;
signal bh537_wm25_10_c4, bh537_wm25_10_c5, bh537_wm25_10_c6 :  std_logic;
signal bh537_wm24_9_c4, bh537_wm24_9_c5, bh537_wm24_9_c6 :  std_logic;
signal bh537_wm23_9_c4, bh537_wm23_9_c5, bh537_wm23_9_c6 :  std_logic;
signal bh537_wm22_9_c4, bh537_wm22_9_c5, bh537_wm22_9_c6 :  std_logic;
signal bh537_wm21_10_c4, bh537_wm21_10_c5, bh537_wm21_10_c6 :  std_logic;
signal bh537_wm20_8_c4, bh537_wm20_8_c5, bh537_wm20_8_c6 :  std_logic;
signal bh537_wm19_9_c4, bh537_wm19_9_c5, bh537_wm19_9_c6 :  std_logic;
signal bh537_wm18_9_c4, bh537_wm18_9_c5, bh537_wm18_9_c6 :  std_logic;
signal bh537_wm17_8_c4, bh537_wm17_8_c5, bh537_wm17_8_c6 :  std_logic;
signal bh537_wm16_8_c4, bh537_wm16_8_c5, bh537_wm16_8_c6 :  std_logic;
signal bh537_wm15_7_c4, bh537_wm15_7_c5, bh537_wm15_7_c6 :  std_logic;
signal bh537_wm14_5_c4, bh537_wm14_5_c5, bh537_wm14_5_c6 :  std_logic;
signal bh537_wm13_5_c4, bh537_wm13_5_c5, bh537_wm13_5_c6 :  std_logic;
signal bh537_wm12_5_c4, bh537_wm12_5_c5, bh537_wm12_5_c6 :  std_logic;
signal bh537_wm11_3_c4, bh537_wm11_3_c5, bh537_wm11_3_c6 :  std_logic;
signal bh537_wm10_2_c4, bh537_wm10_2_c5, bh537_wm10_2_c6 :  std_logic;
signal bh537_wm9_2_c4, bh537_wm9_2_c5, bh537_wm9_2_c6 :  std_logic;
signal bh537_wm8_1_c4, bh537_wm8_1_c5, bh537_wm8_1_c6 :  std_logic;
signal bh537_wm7_0_c4 :  std_logic;
signal bh537_wm6_0_c4 :  std_logic;
signal bh537_wm5_0_c4 :  std_logic;
signal bh537_wm4_0_c4 :  std_logic;
signal bh537_wm3_0_c4 :  std_logic;
signal bh537_wm2_0_c4 :  std_logic;
signal bh537_wm42_5_c0, bh537_wm42_5_c1, bh537_wm42_5_c2, bh537_wm42_5_c3, bh537_wm42_5_c4, bh537_wm42_5_c5, bh537_wm42_5_c6, bh537_wm42_5_c7 :  std_logic;
signal bh537_wm33_12_c0, bh537_wm33_12_c1, bh537_wm33_12_c2, bh537_wm33_12_c3, bh537_wm33_12_c4, bh537_wm33_12_c5, bh537_wm33_12_c6, bh537_wm33_12_c7 :  std_logic;
signal bh537_wm32_11_c0, bh537_wm32_11_c1, bh537_wm32_11_c2, bh537_wm32_11_c3, bh537_wm32_11_c4, bh537_wm32_11_c5, bh537_wm32_11_c6 :  std_logic;
signal bh537_wm31_10_c0, bh537_wm31_10_c1, bh537_wm31_10_c2, bh537_wm31_10_c3, bh537_wm31_10_c4, bh537_wm31_10_c5, bh537_wm31_10_c6 :  std_logic;
signal bh537_wm30_11_c0, bh537_wm30_11_c1, bh537_wm30_11_c2, bh537_wm30_11_c3, bh537_wm30_11_c4, bh537_wm30_11_c5, bh537_wm30_11_c6 :  std_logic;
signal bh537_wm28_10_c0, bh537_wm28_10_c1, bh537_wm28_10_c2, bh537_wm28_10_c3, bh537_wm28_10_c4, bh537_wm28_10_c5, bh537_wm28_10_c6, bh537_wm28_10_c7 :  std_logic;
signal bh537_wm27_10_c0, bh537_wm27_10_c1, bh537_wm27_10_c2, bh537_wm27_10_c3, bh537_wm27_10_c4, bh537_wm27_10_c5, bh537_wm27_10_c6 :  std_logic;
signal bh537_wm26_10_c0, bh537_wm26_10_c1, bh537_wm26_10_c2, bh537_wm26_10_c3, bh537_wm26_10_c4, bh537_wm26_10_c5, bh537_wm26_10_c6 :  std_logic;
signal bh537_wm24_10_c0, bh537_wm24_10_c1, bh537_wm24_10_c2, bh537_wm24_10_c3, bh537_wm24_10_c4, bh537_wm24_10_c5, bh537_wm24_10_c6 :  std_logic;
signal bh537_wm23_10_c0, bh537_wm23_10_c1, bh537_wm23_10_c2, bh537_wm23_10_c3, bh537_wm23_10_c4, bh537_wm23_10_c5, bh537_wm23_10_c6 :  std_logic;
signal bh537_wm22_10_c0, bh537_wm22_10_c1, bh537_wm22_10_c2, bh537_wm22_10_c3, bh537_wm22_10_c4, bh537_wm22_10_c5, bh537_wm22_10_c6, bh537_wm22_10_c7 :  std_logic;
signal bh537_wm21_11_c0, bh537_wm21_11_c1, bh537_wm21_11_c2, bh537_wm21_11_c3, bh537_wm21_11_c4, bh537_wm21_11_c5, bh537_wm21_11_c6 :  std_logic;
signal bh537_wm19_10_c0 :  std_logic;
signal bh537_wm18_10_c0, bh537_wm18_10_c1, bh537_wm18_10_c2, bh537_wm18_10_c3, bh537_wm18_10_c4, bh537_wm18_10_c5, bh537_wm18_10_c6 :  std_logic;
signal bh537_wm14_6_c0 :  std_logic;
signal bh537_wm10_3_c0, bh537_wm10_3_c1, bh537_wm10_3_c2, bh537_wm10_3_c3, bh537_wm10_3_c4, bh537_wm10_3_c5, bh537_wm10_3_c6 :  std_logic;
signal bh537_wm7_1_c0, bh537_wm7_1_c1, bh537_wm7_1_c2, bh537_wm7_1_c3, bh537_wm7_1_c4 :  std_logic;
signal bh537_wm6_1_c0, bh537_wm6_1_c1, bh537_wm6_1_c2, bh537_wm6_1_c3, bh537_wm6_1_c4 :  std_logic;
signal bh537_wm5_1_c0, bh537_wm5_1_c1, bh537_wm5_1_c2, bh537_wm5_1_c3, bh537_wm5_1_c4 :  std_logic;
signal bh537_wm4_1_c0, bh537_wm4_1_c1, bh537_wm4_1_c2, bh537_wm4_1_c3, bh537_wm4_1_c4 :  std_logic;
signal bh537_wm3_1_c0, bh537_wm3_1_c1, bh537_wm3_1_c2, bh537_wm3_1_c3, bh537_wm3_1_c4 :  std_logic;
signal bh537_wm1_0_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid782_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid782_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid782_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm52_2_c7, bh537_wm52_2_c8 :  std_logic;
signal bh537_wm51_2_c7, bh537_wm51_2_c8 :  std_logic;
signal bh537_wm50_2_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid782_Out0_copy783_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid784_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid784_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid784_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm50_3_c7 :  std_logic;
signal bh537_wm49_2_c7 :  std_logic;
signal bh537_wm48_2_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid784_Out0_copy785_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid786_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid786_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid786_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm48_3_c7 :  std_logic;
signal bh537_wm47_2_c7 :  std_logic;
signal bh537_wm46_2_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid786_Out0_copy787_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid790_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid790_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm46_3_c7 :  std_logic;
signal bh537_wm45_3_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid790_Out0_copy791_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid792_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid792_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid792_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm45_4_c7 :  std_logic;
signal bh537_wm44_3_c7 :  std_logic;
signal bh537_wm43_4_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid792_Out0_copy793_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid794_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid794_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm43_5_c7 :  std_logic;
signal bh537_wm42_6_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid794_Out0_copy795_c7 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid798_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid798_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm42_7_c7 :  std_logic;
signal bh537_wm41_7_c7 :  std_logic;
signal bh537_wm40_7_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid798_Out0_copy799_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid800_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid800_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm41_8_c7 :  std_logic;
signal bh537_wm40_8_c7 :  std_logic;
signal bh537_wm39_9_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid800_Out0_copy801_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid802_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid802_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm40_9_c7 :  std_logic;
signal bh537_wm39_10_c7 :  std_logic;
signal bh537_wm38_9_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid802_Out0_copy803_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid804_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid804_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm39_11_c7 :  std_logic;
signal bh537_wm38_10_c7 :  std_logic;
signal bh537_wm37_10_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid804_Out0_copy805_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid806_In0_c6, Compressor_23_3_Freq300_uid781_bh537_uid806_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid806_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid806_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm39_12_c7 :  std_logic;
signal bh537_wm38_11_c7 :  std_logic;
signal bh537_wm37_11_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid806_Out0_copy807_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid808_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid808_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm38_12_c6, bh537_wm38_12_c7 :  std_logic;
signal bh537_wm37_12_c6, bh537_wm37_12_c7 :  std_logic;
signal bh537_wm36_11_c6 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid808_Out0_copy809_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid810_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid810_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm37_13_c7 :  std_logic;
signal bh537_wm36_12_c7 :  std_logic;
signal bh537_wm35_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid810_Out0_copy811_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid814_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid814_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid814_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid814_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm37_14_c7 :  std_logic;
signal bh537_wm36_13_c7 :  std_logic;
signal bh537_wm35_12_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid814_Out0_copy815_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid816_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid816_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm36_14_c7 :  std_logic;
signal bh537_wm35_13_c7 :  std_logic;
signal bh537_wm34_10_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid816_Out0_copy817_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid818_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid818_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid818_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid818_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm36_15_c7 :  std_logic;
signal bh537_wm35_14_c7 :  std_logic;
signal bh537_wm34_11_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid818_Out0_copy819_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid820_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid820_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm35_15_c7 :  std_logic;
signal bh537_wm34_12_c7 :  std_logic;
signal bh537_wm33_13_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid820_Out0_copy821_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid822_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid822_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid822_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid822_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm35_16_c7 :  std_logic;
signal bh537_wm34_13_c7 :  std_logic;
signal bh537_wm33_14_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid822_Out0_copy823_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid824_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid824_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm34_14_c7 :  std_logic;
signal bh537_wm33_15_c7 :  std_logic;
signal bh537_wm32_12_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid824_Out0_copy825_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid826_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid826_Out0_c6 :  std_logic_vector(1 downto 0);
signal bh537_wm34_15_c6, bh537_wm34_15_c7 :  std_logic;
signal bh537_wm33_16_c6, bh537_wm33_16_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid826_Out0_copy827_c6 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid828_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid828_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm33_17_c7 :  std_logic;
signal bh537_wm32_13_c7 :  std_logic;
signal bh537_wm31_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid828_Out0_copy829_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid830_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid830_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm33_18_c7 :  std_logic;
signal bh537_wm32_14_c7 :  std_logic;
signal bh537_wm31_12_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid830_Out0_copy831_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid832_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid832_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm32_15_c7 :  std_logic;
signal bh537_wm31_13_c7 :  std_logic;
signal bh537_wm30_12_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid832_Out0_copy833_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid834_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid834_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm32_16_c6, bh537_wm32_16_c7 :  std_logic;
signal bh537_wm31_14_c6, bh537_wm31_14_c7 :  std_logic;
signal bh537_wm30_13_c6, bh537_wm30_13_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid834_Out0_copy835_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid836_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid836_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm31_15_c7 :  std_logic;
signal bh537_wm30_14_c7 :  std_logic;
signal bh537_wm29_12_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid836_Out0_copy837_c7 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid839_bh537_uid840_In0_c6 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid839_bh537_uid840_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm31_16_c6, bh537_wm31_16_c7 :  std_logic;
signal bh537_wm30_15_c6, bh537_wm30_15_c7 :  std_logic;
signal bh537_wm29_13_c6, bh537_wm29_13_c7 :  std_logic;
signal Compressor_5_3_Freq300_uid839_bh537_uid840_Out0_copy841_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid842_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid842_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm30_16_c7 :  std_logic;
signal bh537_wm29_14_c7 :  std_logic;
signal bh537_wm28_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid842_Out0_copy843_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid844_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid844_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm30_17_c6, bh537_wm30_17_c7 :  std_logic;
signal bh537_wm29_15_c6, bh537_wm29_15_c7 :  std_logic;
signal bh537_wm28_12_c6, bh537_wm28_12_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid844_Out0_copy845_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid846_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid846_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm29_16_c7 :  std_logic;
signal bh537_wm28_13_c7 :  std_logic;
signal bh537_wm27_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid846_Out0_copy847_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid848_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid848_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm29_17_c6, bh537_wm29_17_c7 :  std_logic;
signal bh537_wm28_14_c6, bh537_wm28_14_c7 :  std_logic;
signal bh537_wm27_12_c6, bh537_wm27_12_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid848_Out0_copy849_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid850_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid850_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm28_15_c7 :  std_logic;
signal bh537_wm27_13_c7 :  std_logic;
signal bh537_wm26_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid850_Out0_copy851_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid852_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid852_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid852_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid852_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm28_16_c7 :  std_logic;
signal bh537_wm27_14_c7 :  std_logic;
signal bh537_wm26_12_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid852_Out0_copy853_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid854_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid854_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm27_15_c6, bh537_wm27_15_c7 :  std_logic;
signal bh537_wm26_13_c6, bh537_wm26_13_c7 :  std_logic;
signal bh537_wm25_11_c6, bh537_wm25_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid854_Out0_copy855_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid856_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid856_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid856_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid856_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm27_16_c7 :  std_logic;
signal bh537_wm26_14_c7 :  std_logic;
signal bh537_wm25_12_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid856_Out0_copy857_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid858_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid858_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm26_15_c6, bh537_wm26_15_c7 :  std_logic;
signal bh537_wm25_13_c6, bh537_wm25_13_c7 :  std_logic;
signal bh537_wm24_11_c6, bh537_wm24_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid858_Out0_copy859_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid860_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid860_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid860_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid860_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm26_16_c7 :  std_logic;
signal bh537_wm25_14_c7 :  std_logic;
signal bh537_wm24_12_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid860_Out0_copy861_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid862_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid862_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm25_15_c6, bh537_wm25_15_c7 :  std_logic;
signal bh537_wm24_13_c6, bh537_wm24_13_c7 :  std_logic;
signal bh537_wm23_11_c6, bh537_wm23_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid862_Out0_copy863_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid864_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid864_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid864_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid864_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm25_16_c7 :  std_logic;
signal bh537_wm24_14_c7 :  std_logic;
signal bh537_wm23_12_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid864_Out0_copy865_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid866_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid866_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm24_15_c6, bh537_wm24_15_c7 :  std_logic;
signal bh537_wm23_13_c6, bh537_wm23_13_c7 :  std_logic;
signal bh537_wm22_11_c6, bh537_wm22_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid866_Out0_copy867_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid868_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid868_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid868_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid868_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm24_16_c7 :  std_logic;
signal bh537_wm23_14_c7 :  std_logic;
signal bh537_wm22_12_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid868_Out0_copy869_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid870_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid870_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm23_15_c6, bh537_wm23_15_c7 :  std_logic;
signal bh537_wm22_13_c6, bh537_wm22_13_c7 :  std_logic;
signal bh537_wm21_12_c6, bh537_wm21_12_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid870_Out0_copy871_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid872_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid872_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid872_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid872_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm23_16_c7 :  std_logic;
signal bh537_wm22_14_c7 :  std_logic;
signal bh537_wm21_13_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid872_Out0_copy873_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid874_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid874_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm22_15_c6, bh537_wm22_15_c7 :  std_logic;
signal bh537_wm21_14_c6, bh537_wm21_14_c7 :  std_logic;
signal bh537_wm20_9_c6, bh537_wm20_9_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid874_Out0_copy875_c6 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid876_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid876_Out0_c6 :  std_logic_vector(1 downto 0);
signal bh537_wm22_16_c6, bh537_wm22_16_c7 :  std_logic;
signal bh537_wm21_15_c6, bh537_wm21_15_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid876_Out0_copy877_c6 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid878_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid878_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm21_16_c7 :  std_logic;
signal bh537_wm20_10_c7 :  std_logic;
signal bh537_wm19_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid878_Out0_copy879_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid880_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid880_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm21_17_c6, bh537_wm21_17_c7 :  std_logic;
signal bh537_wm20_11_c6, bh537_wm20_11_c7 :  std_logic;
signal bh537_wm19_12_c6, bh537_wm19_12_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid880_Out0_copy881_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid882_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid882_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm20_12_c7 :  std_logic;
signal bh537_wm19_13_c7 :  std_logic;
signal bh537_wm18_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid882_Out0_copy883_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid884_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid884_Out0_c6 :  std_logic_vector(1 downto 0);
signal bh537_wm20_13_c6, bh537_wm20_13_c7 :  std_logic;
signal bh537_wm19_14_c6, bh537_wm19_14_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid884_Out0_copy885_c6 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid886_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid886_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm19_15_c7 :  std_logic;
signal bh537_wm18_12_c7 :  std_logic;
signal bh537_wm17_9_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid886_Out0_copy887_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid888_In0_c6, Compressor_14_3_Freq300_uid813_bh537_uid888_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid888_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid888_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm19_16_c7 :  std_logic;
signal bh537_wm18_13_c7 :  std_logic;
signal bh537_wm17_10_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid888_Out0_copy889_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid890_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid890_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm18_14_c6, bh537_wm18_14_c7 :  std_logic;
signal bh537_wm17_11_c6, bh537_wm17_11_c7 :  std_logic;
signal bh537_wm16_9_c6, bh537_wm16_9_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid890_Out0_copy891_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid892_In0_c6 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c6 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid892_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm18_15_c6, bh537_wm18_15_c7 :  std_logic;
signal bh537_wm17_12_c6, bh537_wm17_12_c7 :  std_logic;
signal bh537_wm16_10_c6, bh537_wm16_10_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid892_Out0_copy893_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid894_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid894_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm17_13_c7 :  std_logic;
signal bh537_wm16_11_c7 :  std_logic;
signal bh537_wm15_8_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid894_Out0_copy895_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid896_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid896_Out0_c6 :  std_logic_vector(1 downto 0);
signal bh537_wm17_14_c6, bh537_wm17_14_c7 :  std_logic;
signal bh537_wm16_12_c6, bh537_wm16_12_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid896_Out0_copy897_c6 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid898_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid898_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm16_13_c6, bh537_wm16_13_c7 :  std_logic;
signal bh537_wm15_9_c6, bh537_wm15_9_c7 :  std_logic;
signal bh537_wm14_7_c6 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid898_Out0_copy899_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid900_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid900_In1_c6 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid900_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm16_14_c6, bh537_wm16_14_c7 :  std_logic;
signal bh537_wm15_10_c6, bh537_wm15_10_c7 :  std_logic;
signal bh537_wm14_8_c6 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid900_Out0_copy901_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid902_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid902_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm15_11_c6, bh537_wm15_11_c7 :  std_logic;
signal bh537_wm14_9_c6 :  std_logic;
signal bh537_wm13_6_c6 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid902_Out0_copy903_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid904_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid904_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm14_10_c6 :  std_logic;
signal bh537_wm13_7_c6 :  std_logic;
signal bh537_wm12_6_c6 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid904_Out0_copy905_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid906_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid906_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm13_8_c6 :  std_logic;
signal bh537_wm12_7_c6 :  std_logic;
signal bh537_wm11_4_c6 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid906_Out0_copy907_c6 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid908_In0_c6 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid908_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm12_8_c6 :  std_logic;
signal bh537_wm11_5_c6 :  std_logic;
signal bh537_wm10_4_c6 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid908_Out0_copy909_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid910_In0_c6 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid910_In1_c6 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid910_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm11_6_c6 :  std_logic;
signal bh537_wm10_5_c6 :  std_logic;
signal bh537_wm9_3_c6 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid910_Out0_copy911_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid912_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid912_In1_c6 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid912_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm10_6_c6 :  std_logic;
signal bh537_wm9_4_c6 :  std_logic;
signal bh537_wm8_2_c6 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid912_Out0_copy913_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid914_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid914_In1_c4, Compressor_23_3_Freq300_uid781_bh537_uid914_In1_c5, Compressor_23_3_Freq300_uid781_bh537_uid914_In1_c6 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid914_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm8_3_c6 :  std_logic;
signal bh537_wm7_2_c6 :  std_logic;
signal bh537_wm6_2_c6 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid914_Out0_copy915_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid916_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid916_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid916_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh537_wm6_3_c4, bh537_wm6_3_c5, bh537_wm6_3_c6 :  std_logic;
signal bh537_wm5_2_c4 :  std_logic;
signal bh537_wm4_2_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid916_Out0_copy917_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid918_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid918_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid918_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh537_wm4_3_c4 :  std_logic;
signal bh537_wm3_2_c4 :  std_logic;
signal bh537_wm2_1_c4 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid918_Out0_copy919_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid920_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid920_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid920_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm50_4_c7, bh537_wm50_4_c8 :  std_logic;
signal bh537_wm49_3_c7, bh537_wm49_3_c8 :  std_logic;
signal bh537_wm48_4_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid920_Out0_copy921_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid922_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid922_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid922_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm48_5_c7 :  std_logic;
signal bh537_wm47_3_c7 :  std_logic;
signal bh537_wm46_4_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid922_Out0_copy923_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid924_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid924_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid924_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm46_5_c7 :  std_logic;
signal bh537_wm45_5_c7 :  std_logic;
signal bh537_wm44_4_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid924_Out0_copy925_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid926_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid926_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm44_5_c7 :  std_logic;
signal bh537_wm43_6_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid926_Out0_copy927_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid928_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid928_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid928_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm43_7_c7 :  std_logic;
signal bh537_wm42_8_c7 :  std_logic;
signal bh537_wm41_9_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid928_Out0_copy929_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid930_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid930_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm41_10_c7 :  std_logic;
signal bh537_wm40_10_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid930_Out0_copy931_c7 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid932_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid932_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid932_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm40_11_c7 :  std_logic;
signal bh537_wm39_13_c7 :  std_logic;
signal bh537_wm38_13_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid932_Out0_copy933_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid934_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid934_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm39_14_c7 :  std_logic;
signal bh537_wm38_14_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid934_Out0_copy935_c7 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid936_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid936_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid936_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm38_15_c7 :  std_logic;
signal bh537_wm37_15_c7 :  std_logic;
signal bh537_wm36_16_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid936_Out0_copy937_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid938_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid938_In1_c6, Compressor_14_3_Freq300_uid813_bh537_uid938_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid938_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm37_16_c7 :  std_logic;
signal bh537_wm36_17_c7 :  std_logic;
signal bh537_wm35_17_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid938_Out0_copy939_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid940_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid940_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm36_18_c7 :  std_logic;
signal bh537_wm35_18_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid940_Out0_copy941_c7 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid942_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid942_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm35_19_c7 :  std_logic;
signal bh537_wm34_16_c7 :  std_logic;
signal bh537_wm33_19_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid942_Out0_copy943_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid944_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid944_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm34_17_c7 :  std_logic;
signal bh537_wm33_20_c7 :  std_logic;
signal bh537_wm32_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid944_Out0_copy945_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid946_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid946_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm33_21_c7 :  std_logic;
signal bh537_wm32_18_c7 :  std_logic;
signal bh537_wm31_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid946_Out0_copy947_c7 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid839_bh537_uid948_In0_c7 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid839_bh537_uid948_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm32_19_c7 :  std_logic;
signal bh537_wm31_18_c7 :  std_logic;
signal bh537_wm30_18_c7 :  std_logic;
signal Compressor_5_3_Freq300_uid839_bh537_uid948_Out0_copy949_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid950_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid950_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm31_19_c7 :  std_logic;
signal bh537_wm30_19_c7 :  std_logic;
signal bh537_wm29_18_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid950_Out0_copy951_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid952_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid952_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm30_20_c7 :  std_logic;
signal bh537_wm29_19_c7 :  std_logic;
signal bh537_wm28_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid952_Out0_copy953_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid954_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid954_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm29_20_c7 :  std_logic;
signal bh537_wm28_18_c7 :  std_logic;
signal bh537_wm27_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid954_Out0_copy955_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid956_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid956_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm28_19_c7 :  std_logic;
signal bh537_wm27_18_c7 :  std_logic;
signal bh537_wm26_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid956_Out0_copy957_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid958_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid958_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm27_19_c7 :  std_logic;
signal bh537_wm26_18_c7 :  std_logic;
signal bh537_wm25_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid958_Out0_copy959_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid960_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid960_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm26_19_c7 :  std_logic;
signal bh537_wm25_18_c7 :  std_logic;
signal bh537_wm24_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid960_Out0_copy961_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid962_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid962_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm25_19_c7 :  std_logic;
signal bh537_wm24_18_c7 :  std_logic;
signal bh537_wm23_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid962_Out0_copy963_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid964_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid964_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm24_19_c7 :  std_logic;
signal bh537_wm23_18_c7 :  std_logic;
signal bh537_wm22_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid964_Out0_copy965_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid966_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid966_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm23_19_c7 :  std_logic;
signal bh537_wm22_18_c7 :  std_logic;
signal bh537_wm21_18_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid966_Out0_copy967_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid968_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid968_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm22_19_c7 :  std_logic;
signal bh537_wm21_19_c7 :  std_logic;
signal bh537_wm20_14_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid968_Out0_copy969_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid970_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid970_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm21_20_c7 :  std_logic;
signal bh537_wm20_15_c7 :  std_logic;
signal bh537_wm19_17_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid970_Out0_copy971_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid972_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c6, Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid972_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm20_16_c7 :  std_logic;
signal bh537_wm19_18_c7 :  std_logic;
signal bh537_wm18_16_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid972_Out0_copy973_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid974_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid974_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm19_19_c7 :  std_logic;
signal bh537_wm18_17_c7 :  std_logic;
signal bh537_wm17_15_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid974_Out0_copy975_c7 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid839_bh537_uid976_In0_c7 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid839_bh537_uid976_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm18_18_c7 :  std_logic;
signal bh537_wm17_16_c7 :  std_logic;
signal bh537_wm16_15_c7 :  std_logic;
signal Compressor_5_3_Freq300_uid839_bh537_uid976_Out0_copy977_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid978_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid978_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm17_17_c7 :  std_logic;
signal bh537_wm16_16_c7 :  std_logic;
signal bh537_wm15_12_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid978_Out0_copy979_c7 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid980_In0_c7 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid797_bh537_uid980_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm16_17_c7 :  std_logic;
signal bh537_wm15_13_c7 :  std_logic;
signal bh537_wm14_11_c7 :  std_logic;
signal Compressor_6_3_Freq300_uid797_bh537_uid980_Out0_copy981_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid982_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c6, Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid982_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm15_14_c7 :  std_logic;
signal bh537_wm14_12_c7 :  std_logic;
signal bh537_wm13_9_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid982_Out0_copy983_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid984_In0_c6 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c6 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid984_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm14_13_c6, bh537_wm14_13_c7 :  std_logic;
signal bh537_wm13_10_c6, bh537_wm13_10_c7 :  std_logic;
signal bh537_wm12_9_c6 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid984_Out0_copy985_c6 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid986_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid986_Out0_c6 :  std_logic_vector(1 downto 0);
signal bh537_wm13_11_c6, bh537_wm13_11_c7 :  std_logic;
signal bh537_wm12_10_c6 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid986_Out0_copy987_c6 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid988_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid988_In1_c6 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid988_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm12_11_c6 :  std_logic;
signal bh537_wm11_7_c6 :  std_logic;
signal bh537_wm10_7_c6 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid988_Out0_copy989_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid990_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid990_In1_c6 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid990_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm10_8_c6 :  std_logic;
signal bh537_wm9_5_c6 :  std_logic;
signal bh537_wm8_4_c6 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid990_Out0_copy991_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid992_In0_c6 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid992_In1_c6 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid992_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm8_5_c6 :  std_logic;
signal bh537_wm7_3_c6 :  std_logic;
signal bh537_wm6_4_c6 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid992_Out0_copy993_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid994_In0_c6 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid994_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid994_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid994_In1_c6 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid994_Out0_c6 :  std_logic_vector(2 downto 0);
signal bh537_wm6_5_c6 :  std_logic;
signal bh537_wm5_3_c6 :  std_logic;
signal bh537_wm4_4_c6 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid994_Out0_copy995_c6 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid996_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid996_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid996_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh537_wm4_5_c4, bh537_wm4_5_c5, bh537_wm4_5_c6 :  std_logic;
signal bh537_wm3_3_c4 :  std_logic;
signal bh537_wm2_2_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid996_Out0_copy997_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid998_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid998_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid998_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid998_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid998_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid998_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid998_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh537_wm2_3_c4 :  std_logic;
signal bh537_wm1_1_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid998_Out0_copy999_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1000_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1000_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1000_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm48_6_c7, bh537_wm48_6_c8 :  std_logic;
signal bh537_wm47_4_c7, bh537_wm47_4_c8 :  std_logic;
signal bh537_wm46_6_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1000_Out0_copy1001_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1002_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1002_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1002_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm46_7_c7 :  std_logic;
signal bh537_wm45_6_c7 :  std_logic;
signal bh537_wm44_6_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1002_Out0_copy1003_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1004_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1004_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1004_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm44_7_c7 :  std_logic;
signal bh537_wm43_8_c7 :  std_logic;
signal bh537_wm42_9_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1004_Out0_copy1005_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1006_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1006_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1006_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm41_11_c7 :  std_logic;
signal bh537_wm40_12_c7, bh537_wm40_12_c8 :  std_logic;
signal bh537_wm39_15_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1006_Out0_copy1007_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1008_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1008_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm39_16_c7 :  std_logic;
signal bh537_wm38_16_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid1008_Out0_copy1009_c7 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1010_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1010_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1010_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm38_17_c7 :  std_logic;
signal bh537_wm37_17_c7 :  std_logic;
signal bh537_wm36_19_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1010_Out0_copy1011_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1012_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c6, Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1012_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm36_20_c7 :  std_logic;
signal bh537_wm35_20_c7 :  std_logic;
signal bh537_wm34_18_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1012_Out0_copy1013_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1014_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1014_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1014_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm35_21_c7 :  std_logic;
signal bh537_wm34_19_c7 :  std_logic;
signal bh537_wm33_22_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1014_Out0_copy1015_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1016_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c6, Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1016_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm33_23_c7 :  std_logic;
signal bh537_wm32_20_c7 :  std_logic;
signal bh537_wm31_20_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1016_Out0_copy1017_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1018_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1018_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm32_21_c7 :  std_logic;
signal bh537_wm31_21_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid1018_Out0_copy1019_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1020_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1020_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1020_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm31_22_c7 :  std_logic;
signal bh537_wm30_21_c7 :  std_logic;
signal bh537_wm29_21_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1020_Out0_copy1021_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1022_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1022_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm29_22_c7 :  std_logic;
signal bh537_wm28_20_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid1022_Out0_copy1023_c7 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1024_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c6, Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1024_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm28_21_c7 :  std_logic;
signal bh537_wm27_20_c7 :  std_logic;
signal bh537_wm26_20_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1024_Out0_copy1025_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1026_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1026_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm27_21_c7 :  std_logic;
signal bh537_wm26_21_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid1026_Out0_copy1027_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1028_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1028_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1028_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm26_22_c7 :  std_logic;
signal bh537_wm25_20_c7 :  std_logic;
signal bh537_wm24_20_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1028_Out0_copy1029_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1030_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1030_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1030_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm24_21_c7 :  std_logic;
signal bh537_wm23_20_c7 :  std_logic;
signal bh537_wm22_20_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1030_Out0_copy1031_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1032_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c6, Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1032_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm22_21_c7 :  std_logic;
signal bh537_wm21_21_c7 :  std_logic;
signal bh537_wm20_17_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1032_Out0_copy1033_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1034_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1034_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm21_22_c7 :  std_logic;
signal bh537_wm20_18_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid1034_Out0_copy1035_c7 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1036_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c0, Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c1, Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c2, Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c3, Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c6, Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1036_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm20_19_c7 :  std_logic;
signal bh537_wm19_20_c7 :  std_logic;
signal bh537_wm18_19_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1036_Out0_copy1037_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1038_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1038_Out0_c7 :  std_logic_vector(1 downto 0);
signal bh537_wm19_21_c7 :  std_logic;
signal bh537_wm18_20_c7 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid1038_Out0_copy1039_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1040_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1040_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1040_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm18_21_c7 :  std_logic;
signal bh537_wm17_18_c7 :  std_logic;
signal bh537_wm16_18_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1040_Out0_copy1041_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1042_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1042_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1042_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm16_19_c7 :  std_logic;
signal bh537_wm15_15_c7 :  std_logic;
signal bh537_wm14_14_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1042_Out0_copy1043_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1044_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1044_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1044_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm14_15_c7 :  std_logic;
signal bh537_wm13_12_c7 :  std_logic;
signal bh537_wm12_12_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1044_Out0_copy1045_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1046_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1046_In1_c6 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm12_13_c7 :  std_logic;
signal bh537_wm11_8_c7 :  std_logic;
signal bh537_wm10_9_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_copy1047_c6, Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_copy1047_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1048_In0_c6 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1048_In1_c6 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm10_10_c7 :  std_logic;
signal bh537_wm9_6_c7 :  std_logic;
signal bh537_wm8_6_c7 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_copy1049_c6, Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_copy1049_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1050_In0_c6 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1050_In1_c6 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm8_7_c7 :  std_logic;
signal bh537_wm7_4_c7 :  std_logic;
signal bh537_wm6_6_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_copy1051_c6, Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_copy1051_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1052_In0_c6 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1052_In1_c6 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm6_7_c7 :  std_logic;
signal bh537_wm5_4_c7 :  std_logic;
signal bh537_wm4_6_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_copy1053_c6, Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_copy1053_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1054_In0_c6 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1054_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid1054_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid1054_In1_c6 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm4_7_c7 :  std_logic;
signal bh537_wm3_4_c7 :  std_logic;
signal bh537_wm2_4_c7 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_copy1055_c6, Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_copy1055_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1056_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1056_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1056_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh537_wm2_5_c4, bh537_wm2_5_c5, bh537_wm2_5_c6, bh537_wm2_5_c7 :  std_logic;
signal bh537_wm1_2_c4 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1056_Out0_copy1057_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1058_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1058_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm46_8_c8 :  std_logic;
signal bh537_wm45_7_c8 :  std_logic;
signal bh537_wm44_8_c8 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_copy1059_c7, Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_copy1059_c8 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1060_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1060_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm44_9_c8 :  std_logic;
signal bh537_wm43_9_c8 :  std_logic;
signal bh537_wm42_10_c8 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_copy1061_c7, Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_copy1061_c8 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1062_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1062_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm42_11_c8 :  std_logic;
signal bh537_wm41_12_c8 :  std_logic;
signal bh537_wm40_13_c8 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_copy1063_c7, Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_copy1063_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1064_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1064_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm39_17_c8 :  std_logic;
signal bh537_wm38_18_c8 :  std_logic;
signal bh537_wm37_18_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_copy1065_c7, Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_copy1065_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1066_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1066_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm37_19_c8 :  std_logic;
signal bh537_wm36_21_c8 :  std_logic;
signal bh537_wm35_22_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_copy1067_c7, Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_copy1067_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1068_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1068_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm35_23_c8 :  std_logic;
signal bh537_wm34_20_c8 :  std_logic;
signal bh537_wm33_24_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_copy1069_c7, Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_copy1069_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1070_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1070_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm33_25_c8 :  std_logic;
signal bh537_wm32_22_c8 :  std_logic;
signal bh537_wm31_23_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_copy1071_c7, Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_copy1071_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1072_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1072_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm31_24_c8 :  std_logic;
signal bh537_wm30_22_c8 :  std_logic;
signal bh537_wm29_23_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_copy1073_c7, Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_copy1073_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1074_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1074_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm29_24_c8 :  std_logic;
signal bh537_wm28_22_c8 :  std_logic;
signal bh537_wm27_22_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_copy1075_c7, Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_copy1075_c8 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1076_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_c8 :  std_logic_vector(1 downto 0);
signal bh537_wm27_23_c8 :  std_logic;
signal bh537_wm26_23_c8 :  std_logic;
signal Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_copy1077_c7, Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_copy1077_c8 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1078_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1078_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm26_24_c8 :  std_logic;
signal bh537_wm25_21_c8 :  std_logic;
signal bh537_wm24_22_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_copy1079_c7, Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_copy1079_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1080_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1080_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm24_23_c8 :  std_logic;
signal bh537_wm23_21_c8 :  std_logic;
signal bh537_wm22_22_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_copy1081_c7, Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_copy1081_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1082_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1082_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm22_23_c8 :  std_logic;
signal bh537_wm21_23_c8 :  std_logic;
signal bh537_wm20_20_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_copy1083_c7, Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_copy1083_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1084_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1084_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm20_21_c8 :  std_logic;
signal bh537_wm19_22_c8 :  std_logic;
signal bh537_wm18_22_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_copy1085_c7, Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_copy1085_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1086_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1086_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm18_23_c8 :  std_logic;
signal bh537_wm17_19_c8 :  std_logic;
signal bh537_wm16_20_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_copy1087_c7, Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_copy1087_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1088_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1088_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm16_21_c8 :  std_logic;
signal bh537_wm15_16_c8 :  std_logic;
signal bh537_wm14_16_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_copy1089_c7, Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_copy1089_c8 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1090_In0_c7 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1090_In1_c7 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm14_17_c8 :  std_logic;
signal bh537_wm13_13_c8 :  std_logic;
signal bh537_wm12_14_c8 :  std_logic;
signal Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_copy1091_c7, Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_copy1091_c8 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1092_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1092_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_c8 :  std_logic_vector(2 downto 0);
signal bh537_wm12_15_c8 :  std_logic;
signal bh537_wm11_9_c8 :  std_logic;
signal bh537_wm10_11_c8 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_copy1093_c7, Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_copy1093_c8 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1094_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1094_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1094_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm10_12_c7, bh537_wm10_12_c8 :  std_logic;
signal bh537_wm9_7_c7, bh537_wm9_7_c8 :  std_logic;
signal bh537_wm8_8_c7, bh537_wm8_8_c8 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1094_Out0_copy1095_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1096_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1096_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1096_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm8_9_c7, bh537_wm8_9_c8 :  std_logic;
signal bh537_wm7_5_c7, bh537_wm7_5_c8 :  std_logic;
signal bh537_wm6_8_c7, bh537_wm6_8_c8 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1096_Out0_copy1097_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1098_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1098_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1098_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm6_9_c7, bh537_wm6_9_c8 :  std_logic;
signal bh537_wm5_5_c7, bh537_wm5_5_c8 :  std_logic;
signal bh537_wm4_8_c7, bh537_wm4_8_c8 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1098_Out0_copy1099_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1100_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1100_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1100_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm4_9_c7, bh537_wm4_9_c8 :  std_logic;
signal bh537_wm3_5_c7, bh537_wm3_5_c8 :  std_logic;
signal bh537_wm2_6_c7, bh537_wm2_6_c8 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1100_Out0_copy1101_c7 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1102_In0_c7 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c4, Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c5, Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c6, Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c7 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid813_bh537_uid1102_Out0_c7 :  std_logic_vector(2 downto 0);
signal bh537_wm2_7_c7, bh537_wm2_7_c8 :  std_logic;
signal bh537_wm1_3_c7, bh537_wm1_3_c8 :  std_logic;
signal Compressor_14_3_Freq300_uid813_bh537_uid1102_Out0_copy1103_c7 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh537_24_c8 :  std_logic_vector(24 downto 0);
signal bitheapFinalAdd_bh537_In0_c8 :  std_logic_vector(44 downto 0);
signal bitheapFinalAdd_bh537_In1_c8 :  std_logic_vector(44 downto 0);
signal bitheapFinalAdd_bh537_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh537_Out_c8 :  std_logic_vector(44 downto 0);
signal bitheapResult_bh537_c8 :  std_logic_vector(68 downto 0);
signal RR_c8 :  signed(-1+41 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               bh537_wm41_6_c5 <= bh537_wm41_6_c4;
               bh537_wm40_6_c5 <= bh537_wm40_6_c4;
               bh537_wm39_8_c5 <= bh537_wm39_8_c4;
               bh537_wm38_8_c5 <= bh537_wm38_8_c4;
               bh537_wm37_9_c5 <= bh537_wm37_9_c4;
               bh537_wm36_10_c5 <= bh537_wm36_10_c4;
               bh537_wm35_10_c5 <= bh537_wm35_10_c4;
               bh537_wm34_9_c5 <= bh537_wm34_9_c4;
               bh537_wm33_11_c5 <= bh537_wm33_11_c4;
               bh537_wm32_10_c5 <= bh537_wm32_10_c4;
               bh537_wm31_9_c5 <= bh537_wm31_9_c4;
               bh537_wm30_10_c5 <= bh537_wm30_10_c4;
               bh537_wm29_11_c5 <= bh537_wm29_11_c4;
               bh537_wm28_9_c5 <= bh537_wm28_9_c4;
               bh537_wm27_9_c5 <= bh537_wm27_9_c4;
               bh537_wm26_9_c5 <= bh537_wm26_9_c4;
               bh537_wm25_10_c5 <= bh537_wm25_10_c4;
               bh537_wm24_9_c5 <= bh537_wm24_9_c4;
               bh537_wm23_9_c5 <= bh537_wm23_9_c4;
               bh537_wm22_9_c5 <= bh537_wm22_9_c4;
               bh537_wm21_10_c5 <= bh537_wm21_10_c4;
               bh537_wm20_8_c5 <= bh537_wm20_8_c4;
               bh537_wm19_9_c5 <= bh537_wm19_9_c4;
               bh537_wm18_9_c5 <= bh537_wm18_9_c4;
               bh537_wm17_8_c5 <= bh537_wm17_8_c4;
               bh537_wm16_8_c5 <= bh537_wm16_8_c4;
               bh537_wm15_7_c5 <= bh537_wm15_7_c4;
               bh537_wm14_5_c5 <= bh537_wm14_5_c4;
               bh537_wm13_5_c5 <= bh537_wm13_5_c4;
               bh537_wm12_5_c5 <= bh537_wm12_5_c4;
               bh537_wm11_3_c5 <= bh537_wm11_3_c4;
               bh537_wm10_2_c5 <= bh537_wm10_2_c4;
               bh537_wm9_2_c5 <= bh537_wm9_2_c4;
               bh537_wm8_1_c5 <= bh537_wm8_1_c4;
               bh537_wm42_5_c5 <= bh537_wm42_5_c4;
               bh537_wm33_12_c5 <= bh537_wm33_12_c4;
               bh537_wm32_11_c5 <= bh537_wm32_11_c4;
               bh537_wm31_10_c5 <= bh537_wm31_10_c4;
               bh537_wm30_11_c5 <= bh537_wm30_11_c4;
               bh537_wm28_10_c5 <= bh537_wm28_10_c4;
               bh537_wm27_10_c5 <= bh537_wm27_10_c4;
               bh537_wm26_10_c5 <= bh537_wm26_10_c4;
               bh537_wm24_10_c5 <= bh537_wm24_10_c4;
               bh537_wm23_10_c5 <= bh537_wm23_10_c4;
               bh537_wm22_10_c5 <= bh537_wm22_10_c4;
               bh537_wm21_11_c5 <= bh537_wm21_11_c4;
               bh537_wm18_10_c5 <= bh537_wm18_10_c4;
               bh537_wm10_3_c5 <= bh537_wm10_3_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c4;
               Compressor_23_3_Freq300_uid781_bh537_uid914_In1_c5 <= Compressor_23_3_Freq300_uid781_bh537_uid914_In1_c4;
               bh537_wm6_3_c5 <= bh537_wm6_3_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid994_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid994_In1_c4;
               bh537_wm4_5_c5 <= bh537_wm4_5_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid1054_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid1054_In1_c4;
               bh537_wm2_5_c5 <= bh537_wm2_5_c4;
               Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c5 <= Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c4;
            end if;
            if ce_6 = '1' then
               bh537_wm41_6_c6 <= bh537_wm41_6_c5;
               bh537_wm40_6_c6 <= bh537_wm40_6_c5;
               bh537_wm39_8_c6 <= bh537_wm39_8_c5;
               bh537_wm38_8_c6 <= bh537_wm38_8_c5;
               bh537_wm37_9_c6 <= bh537_wm37_9_c5;
               bh537_wm36_10_c6 <= bh537_wm36_10_c5;
               bh537_wm35_10_c6 <= bh537_wm35_10_c5;
               bh537_wm34_9_c6 <= bh537_wm34_9_c5;
               bh537_wm33_11_c6 <= bh537_wm33_11_c5;
               bh537_wm32_10_c6 <= bh537_wm32_10_c5;
               bh537_wm31_9_c6 <= bh537_wm31_9_c5;
               bh537_wm30_10_c6 <= bh537_wm30_10_c5;
               bh537_wm29_11_c6 <= bh537_wm29_11_c5;
               bh537_wm28_9_c6 <= bh537_wm28_9_c5;
               bh537_wm27_9_c6 <= bh537_wm27_9_c5;
               bh537_wm26_9_c6 <= bh537_wm26_9_c5;
               bh537_wm25_10_c6 <= bh537_wm25_10_c5;
               bh537_wm24_9_c6 <= bh537_wm24_9_c5;
               bh537_wm23_9_c6 <= bh537_wm23_9_c5;
               bh537_wm22_9_c6 <= bh537_wm22_9_c5;
               bh537_wm21_10_c6 <= bh537_wm21_10_c5;
               bh537_wm20_8_c6 <= bh537_wm20_8_c5;
               bh537_wm19_9_c6 <= bh537_wm19_9_c5;
               bh537_wm18_9_c6 <= bh537_wm18_9_c5;
               bh537_wm17_8_c6 <= bh537_wm17_8_c5;
               bh537_wm16_8_c6 <= bh537_wm16_8_c5;
               bh537_wm15_7_c6 <= bh537_wm15_7_c5;
               bh537_wm14_5_c6 <= bh537_wm14_5_c5;
               bh537_wm13_5_c6 <= bh537_wm13_5_c5;
               bh537_wm12_5_c6 <= bh537_wm12_5_c5;
               bh537_wm11_3_c6 <= bh537_wm11_3_c5;
               bh537_wm10_2_c6 <= bh537_wm10_2_c5;
               bh537_wm9_2_c6 <= bh537_wm9_2_c5;
               bh537_wm8_1_c6 <= bh537_wm8_1_c5;
               bh537_wm42_5_c6 <= bh537_wm42_5_c5;
               bh537_wm33_12_c6 <= bh537_wm33_12_c5;
               bh537_wm32_11_c6 <= bh537_wm32_11_c5;
               bh537_wm31_10_c6 <= bh537_wm31_10_c5;
               bh537_wm30_11_c6 <= bh537_wm30_11_c5;
               bh537_wm28_10_c6 <= bh537_wm28_10_c5;
               bh537_wm27_10_c6 <= bh537_wm27_10_c5;
               bh537_wm26_10_c6 <= bh537_wm26_10_c5;
               bh537_wm24_10_c6 <= bh537_wm24_10_c5;
               bh537_wm23_10_c6 <= bh537_wm23_10_c5;
               bh537_wm22_10_c6 <= bh537_wm22_10_c5;
               bh537_wm21_11_c6 <= bh537_wm21_11_c5;
               bh537_wm18_10_c6 <= bh537_wm18_10_c5;
               bh537_wm10_3_c6 <= bh537_wm10_3_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c5;
               Compressor_23_3_Freq300_uid781_bh537_uid914_In1_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid914_In1_c5;
               bh537_wm6_3_c6 <= bh537_wm6_3_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid994_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid994_In1_c5;
               bh537_wm4_5_c6 <= bh537_wm4_5_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid1054_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid1054_In1_c5;
               bh537_wm2_5_c6 <= bh537_wm2_5_c5;
               Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c5;
            end if;
            if ce_7 = '1' then
               bh537_wm21_1_c7 <= bh537_wm21_1_c6;
               bh537_wm21_2_c7 <= bh537_wm21_2_c6;
               bh537_wm29_2_c7 <= bh537_wm29_2_c6;
               bh537_wm28_1_c7 <= bh537_wm28_1_c6;
               bh537_wm33_2_c7 <= bh537_wm33_2_c6;
               bh537_wm32_2_c7 <= bh537_wm32_2_c6;
               bh537_wm31_2_c7 <= bh537_wm31_2_c6;
               bh537_wm30_2_c7 <= bh537_wm30_2_c6;
               bh537_wm29_3_c7 <= bh537_wm29_3_c6;
               bh537_wm37_2_c7 <= bh537_wm37_2_c6;
               bh537_wm36_2_c7 <= bh537_wm36_2_c6;
               bh537_wm35_2_c7 <= bh537_wm35_2_c6;
               bh537_wm34_2_c7 <= bh537_wm34_2_c6;
               bh537_wm33_3_c7 <= bh537_wm33_3_c6;
               bh537_wm21_3_c7 <= bh537_wm21_3_c6;
               bh537_wm30_3_c7 <= bh537_wm30_3_c6;
               bh537_wm29_4_c7 <= bh537_wm29_4_c6;
               bh537_wm28_2_c7 <= bh537_wm28_2_c6;
               bh537_wm33_4_c7 <= bh537_wm33_4_c6;
               bh537_wm32_3_c7 <= bh537_wm32_3_c6;
               bh537_wm31_3_c7 <= bh537_wm31_3_c6;
               bh537_wm30_4_c7 <= bh537_wm30_4_c6;
               bh537_wm29_5_c7 <= bh537_wm29_5_c6;
               bh537_wm36_3_c7 <= bh537_wm36_3_c6;
               bh537_wm35_3_c7 <= bh537_wm35_3_c6;
               bh537_wm34_3_c7 <= bh537_wm34_3_c6;
               bh537_wm33_5_c7 <= bh537_wm33_5_c6;
               bh537_wm32_4_c7 <= bh537_wm32_4_c6;
               bh537_wm39_2_c7 <= bh537_wm39_2_c6;
               bh537_wm37_3_c7 <= bh537_wm37_3_c6;
               bh537_wm36_4_c7 <= bh537_wm36_4_c6;
               bh537_wm35_4_c7 <= bh537_wm35_4_c6;
               bh537_wm28_3_c7 <= bh537_wm28_3_c6;
               bh537_wm32_5_c7 <= bh537_wm32_5_c6;
               bh537_wm31_4_c7 <= bh537_wm31_4_c6;
               bh537_wm30_5_c7 <= bh537_wm30_5_c6;
               bh537_wm28_4_c7 <= bh537_wm28_4_c6;
               bh537_wm35_5_c7 <= bh537_wm35_5_c6;
               bh537_wm34_4_c7 <= bh537_wm34_4_c6;
               bh537_wm33_6_c7 <= bh537_wm33_6_c6;
               bh537_wm31_5_c7 <= bh537_wm31_5_c6;
               bh537_wm37_4_c7 <= bh537_wm37_4_c6;
               bh537_wm36_5_c7 <= bh537_wm36_5_c6;
               bh537_wm35_6_c7 <= bh537_wm35_6_c6;
               bh537_wm34_5_c7 <= bh537_wm34_5_c6;
               bh537_wm41_2_c7 <= bh537_wm41_2_c6;
               bh537_wm40_2_c7 <= bh537_wm40_2_c6;
               bh537_wm39_3_c7 <= bh537_wm39_3_c6;
               bh537_wm37_5_c7 <= bh537_wm37_5_c6;
               bh537_wm28_5_c7 <= bh537_wm28_5_c6;
               bh537_wm34_6_c7 <= bh537_wm34_6_c6;
               bh537_wm33_7_c7 <= bh537_wm33_7_c6;
               bh537_wm36_6_c7 <= bh537_wm36_6_c6;
               bh537_wm33_8_c7 <= bh537_wm33_8_c6;
               bh537_wm40_3_c7 <= bh537_wm40_3_c6;
               bh537_wm39_4_c7 <= bh537_wm39_4_c6;
               bh537_wm43_2_c7 <= bh537_wm43_2_c6;
               bh537_wm42_2_c7 <= bh537_wm42_2_c6;
               bh537_wm41_3_c7 <= bh537_wm41_3_c6;
               bh537_wm40_4_c7 <= bh537_wm40_4_c6;
               bh537_wm39_5_c7 <= bh537_wm39_5_c6;
               bh537_wm33_9_c7 <= bh537_wm33_9_c6;
               bh537_wm33_10_c7 <= bh537_wm33_10_c6;
               bh537_wm42_3_c7 <= bh537_wm42_3_c6;
               bh537_wm41_4_c7 <= bh537_wm41_4_c6;
               bh537_wm40_5_c7 <= bh537_wm40_5_c6;
               bh537_wm45_2_c7 <= bh537_wm45_2_c6;
               bh537_wm44_2_c7 <= bh537_wm44_2_c6;
               bh537_wm43_3_c7 <= bh537_wm43_3_c6;
               bh537_wm42_4_c7 <= bh537_wm42_4_c6;
               bh537_wm41_5_c7 <= bh537_wm41_5_c6;
               bh537_wm20_1_c7 <= bh537_wm20_1_c6;
               bh537_wm19_1_c7 <= bh537_wm19_1_c6;
               bh537_wm17_1_c7 <= bh537_wm17_1_c6;
               bh537_wm19_2_c7 <= bh537_wm19_2_c6;
               bh537_wm17_2_c7 <= bh537_wm17_2_c6;
               bh537_wm21_4_c7 <= bh537_wm21_4_c6;
               bh537_wm20_2_c7 <= bh537_wm20_2_c6;
               bh537_wm19_3_c7 <= bh537_wm19_3_c6;
               bh537_wm17_3_c7 <= bh537_wm17_3_c6;
               bh537_wm21_5_c7 <= bh537_wm21_5_c6;
               bh537_wm20_3_c7 <= bh537_wm20_3_c6;
               bh537_wm19_4_c7 <= bh537_wm19_4_c6;
               bh537_wm17_4_c7 <= bh537_wm17_4_c6;
               bh537_wm20_4_c7 <= bh537_wm20_4_c6;
               bh537_wm17_5_c7 <= bh537_wm17_5_c6;
               bh537_wm20_5_c7 <= bh537_wm20_5_c6;
               bh537_wm19_5_c7 <= bh537_wm19_5_c6;
               bh537_wm41_6_c7 <= bh537_wm41_6_c6;
               bh537_wm40_6_c7 <= bh537_wm40_6_c6;
               bh537_wm38_8_c7 <= bh537_wm38_8_c6;
               bh537_wm33_11_c7 <= bh537_wm33_11_c6;
               bh537_wm42_5_c7 <= bh537_wm42_5_c6;
               bh537_wm33_12_c7 <= bh537_wm33_12_c6;
               bh537_wm28_10_c7 <= bh537_wm28_10_c6;
               bh537_wm22_10_c7 <= bh537_wm22_10_c6;
               Compressor_23_3_Freq300_uid781_bh537_uid806_In0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid806_In0_c6;
               bh537_wm38_12_c7 <= bh537_wm38_12_c6;
               bh537_wm37_12_c7 <= bh537_wm37_12_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid814_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid814_In0_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid818_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid818_In0_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid822_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid822_In0_c6;
               bh537_wm34_15_c7 <= bh537_wm34_15_c6;
               bh537_wm33_16_c7 <= bh537_wm33_16_c6;
               bh537_wm32_16_c7 <= bh537_wm32_16_c6;
               bh537_wm31_14_c7 <= bh537_wm31_14_c6;
               bh537_wm30_13_c7 <= bh537_wm30_13_c6;
               bh537_wm31_16_c7 <= bh537_wm31_16_c6;
               bh537_wm30_15_c7 <= bh537_wm30_15_c6;
               bh537_wm29_13_c7 <= bh537_wm29_13_c6;
               bh537_wm30_17_c7 <= bh537_wm30_17_c6;
               bh537_wm29_15_c7 <= bh537_wm29_15_c6;
               bh537_wm28_12_c7 <= bh537_wm28_12_c6;
               bh537_wm29_17_c7 <= bh537_wm29_17_c6;
               bh537_wm28_14_c7 <= bh537_wm28_14_c6;
               bh537_wm27_12_c7 <= bh537_wm27_12_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid852_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid852_In0_c6;
               bh537_wm27_15_c7 <= bh537_wm27_15_c6;
               bh537_wm26_13_c7 <= bh537_wm26_13_c6;
               bh537_wm25_11_c7 <= bh537_wm25_11_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid856_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid856_In0_c6;
               bh537_wm26_15_c7 <= bh537_wm26_15_c6;
               bh537_wm25_13_c7 <= bh537_wm25_13_c6;
               bh537_wm24_11_c7 <= bh537_wm24_11_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid860_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid860_In0_c6;
               bh537_wm25_15_c7 <= bh537_wm25_15_c6;
               bh537_wm24_13_c7 <= bh537_wm24_13_c6;
               bh537_wm23_11_c7 <= bh537_wm23_11_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid864_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid864_In0_c6;
               bh537_wm24_15_c7 <= bh537_wm24_15_c6;
               bh537_wm23_13_c7 <= bh537_wm23_13_c6;
               bh537_wm22_11_c7 <= bh537_wm22_11_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid868_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid868_In0_c6;
               bh537_wm23_15_c7 <= bh537_wm23_15_c6;
               bh537_wm22_13_c7 <= bh537_wm22_13_c6;
               bh537_wm21_12_c7 <= bh537_wm21_12_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid872_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid872_In0_c6;
               bh537_wm22_15_c7 <= bh537_wm22_15_c6;
               bh537_wm21_14_c7 <= bh537_wm21_14_c6;
               bh537_wm20_9_c7 <= bh537_wm20_9_c6;
               bh537_wm22_16_c7 <= bh537_wm22_16_c6;
               bh537_wm21_15_c7 <= bh537_wm21_15_c6;
               bh537_wm21_17_c7 <= bh537_wm21_17_c6;
               bh537_wm20_11_c7 <= bh537_wm20_11_c6;
               bh537_wm19_12_c7 <= bh537_wm19_12_c6;
               bh537_wm20_13_c7 <= bh537_wm20_13_c6;
               bh537_wm19_14_c7 <= bh537_wm19_14_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid888_In0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid888_In0_c6;
               bh537_wm18_14_c7 <= bh537_wm18_14_c6;
               bh537_wm17_11_c7 <= bh537_wm17_11_c6;
               bh537_wm16_9_c7 <= bh537_wm16_9_c6;
               bh537_wm18_15_c7 <= bh537_wm18_15_c6;
               bh537_wm17_12_c7 <= bh537_wm17_12_c6;
               bh537_wm16_10_c7 <= bh537_wm16_10_c6;
               bh537_wm17_14_c7 <= bh537_wm17_14_c6;
               bh537_wm16_12_c7 <= bh537_wm16_12_c6;
               bh537_wm16_13_c7 <= bh537_wm16_13_c6;
               bh537_wm15_9_c7 <= bh537_wm15_9_c6;
               bh537_wm16_14_c7 <= bh537_wm16_14_c6;
               bh537_wm15_10_c7 <= bh537_wm15_10_c6;
               bh537_wm15_11_c7 <= bh537_wm15_11_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid938_In1_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid938_In1_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c6;
               bh537_wm14_13_c7 <= bh537_wm14_13_c6;
               bh537_wm13_10_c7 <= bh537_wm13_10_c6;
               bh537_wm13_11_c7 <= bh537_wm13_11_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c6;
               Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_copy1047_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_copy1047_c6;
               Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_copy1049_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_copy1049_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_copy1051_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_copy1051_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_copy1053_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_copy1053_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_copy1055_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_copy1055_c6;
               bh537_wm2_5_c7 <= bh537_wm2_5_c6;
               Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c6;
            end if;
            if ce_8 = '1' then
               bh537_wm69_0_c8 <= bh537_wm69_0_c7;
               bh537_wm68_0_c8 <= bh537_wm68_0_c7;
               bh537_wm67_0_c8 <= bh537_wm67_0_c7;
               bh537_wm66_0_c8 <= bh537_wm66_0_c7;
               bh537_wm65_0_c8 <= bh537_wm65_0_c7;
               bh537_wm64_0_c8 <= bh537_wm64_0_c7;
               bh537_wm63_0_c8 <= bh537_wm63_0_c7;
               bh537_wm62_0_c8 <= bh537_wm62_0_c7;
               bh537_wm61_0_c8 <= bh537_wm61_0_c7;
               bh537_wm60_0_c8 <= bh537_wm60_0_c7;
               bh537_wm59_0_c8 <= bh537_wm59_0_c7;
               bh537_wm58_0_c8 <= bh537_wm58_0_c7;
               bh537_wm57_0_c8 <= bh537_wm57_0_c7;
               bh537_wm56_0_c8 <= bh537_wm56_0_c7;
               bh537_wm55_0_c8 <= bh537_wm55_0_c7;
               bh537_wm54_0_c8 <= bh537_wm54_0_c7;
               bh537_wm53_0_c8 <= bh537_wm53_0_c7;
               bh537_wm52_2_c8 <= bh537_wm52_2_c7;
               bh537_wm51_2_c8 <= bh537_wm51_2_c7;
               bh537_wm50_4_c8 <= bh537_wm50_4_c7;
               bh537_wm49_3_c8 <= bh537_wm49_3_c7;
               bh537_wm48_6_c8 <= bh537_wm48_6_c7;
               bh537_wm47_4_c8 <= bh537_wm47_4_c7;
               bh537_wm40_12_c8 <= bh537_wm40_12_c7;
               Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_copy1059_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_copy1059_c7;
               Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_copy1061_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_copy1061_c7;
               Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_copy1063_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_copy1063_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_copy1065_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_copy1065_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_copy1067_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_copy1067_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_copy1069_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_copy1069_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_copy1071_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_copy1071_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_copy1073_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_copy1073_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_copy1075_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_copy1075_c7;
               Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_copy1077_c8 <= Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_copy1077_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_copy1079_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_copy1079_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_copy1081_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_copy1081_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_copy1083_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_copy1083_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_copy1085_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_copy1085_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_copy1087_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_copy1087_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_copy1089_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_copy1089_c7;
               Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_copy1091_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_copy1091_c7;
               Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_copy1093_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_copy1093_c7;
               bh537_wm10_12_c8 <= bh537_wm10_12_c7;
               bh537_wm9_7_c8 <= bh537_wm9_7_c7;
               bh537_wm8_8_c8 <= bh537_wm8_8_c7;
               bh537_wm8_9_c8 <= bh537_wm8_9_c7;
               bh537_wm7_5_c8 <= bh537_wm7_5_c7;
               bh537_wm6_8_c8 <= bh537_wm6_8_c7;
               bh537_wm6_9_c8 <= bh537_wm6_9_c7;
               bh537_wm5_5_c8 <= bh537_wm5_5_c7;
               bh537_wm4_8_c8 <= bh537_wm4_8_c7;
               bh537_wm4_9_c8 <= bh537_wm4_9_c7;
               bh537_wm3_5_c8 <= bh537_wm3_5_c7;
               bh537_wm2_6_c8 <= bh537_wm2_6_c7;
               bh537_wm2_7_c8 <= bh537_wm2_7_c7;
               bh537_wm1_3_c8 <= bh537_wm1_3_c7;
            end if;
         end if;
      end process;
XX_c4 <= signed(X);
YY_c6 <= signed(Y);
AA_c4 <= signed(A);
   tile_0_X_c4 <= X(16 downto 0);
   tile_0_Y_c6 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid539
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 X => tile_0_X_c4,
                 Y => tile_0_Y_c6,
                 R => tile_0_output_c7);

   tile_0_filtered_output_c7 <= unsigned(tile_0_output_c7(40 downto 0));
   bh537_wm69_0_c7 <= tile_0_filtered_output_c7(0);
   bh537_wm68_0_c7 <= tile_0_filtered_output_c7(1);
   bh537_wm67_0_c7 <= tile_0_filtered_output_c7(2);
   bh537_wm66_0_c7 <= tile_0_filtered_output_c7(3);
   bh537_wm65_0_c7 <= tile_0_filtered_output_c7(4);
   bh537_wm64_0_c7 <= tile_0_filtered_output_c7(5);
   bh537_wm63_0_c7 <= tile_0_filtered_output_c7(6);
   bh537_wm62_0_c7 <= tile_0_filtered_output_c7(7);
   bh537_wm61_0_c7 <= tile_0_filtered_output_c7(8);
   bh537_wm60_0_c7 <= tile_0_filtered_output_c7(9);
   bh537_wm59_0_c7 <= tile_0_filtered_output_c7(10);
   bh537_wm58_0_c7 <= tile_0_filtered_output_c7(11);
   bh537_wm57_0_c7 <= tile_0_filtered_output_c7(12);
   bh537_wm56_0_c7 <= tile_0_filtered_output_c7(13);
   bh537_wm55_0_c7 <= tile_0_filtered_output_c7(14);
   bh537_wm54_0_c7 <= tile_0_filtered_output_c7(15);
   bh537_wm53_0_c7 <= tile_0_filtered_output_c7(16);
   bh537_wm52_0_c7 <= tile_0_filtered_output_c7(17);
   bh537_wm51_0_c7 <= tile_0_filtered_output_c7(18);
   bh537_wm50_0_c7 <= tile_0_filtered_output_c7(19);
   bh537_wm49_0_c7 <= tile_0_filtered_output_c7(20);
   bh537_wm48_0_c7 <= tile_0_filtered_output_c7(21);
   bh537_wm47_0_c7 <= tile_0_filtered_output_c7(22);
   bh537_wm46_0_c7 <= tile_0_filtered_output_c7(23);
   bh537_wm45_0_c7 <= tile_0_filtered_output_c7(24);
   bh537_wm44_0_c7 <= tile_0_filtered_output_c7(25);
   bh537_wm43_0_c7 <= tile_0_filtered_output_c7(26);
   bh537_wm42_0_c7 <= tile_0_filtered_output_c7(27);
   bh537_wm41_0_c7 <= tile_0_filtered_output_c7(28);
   bh537_wm40_0_c7 <= tile_0_filtered_output_c7(29);
   bh537_wm39_0_c7 <= tile_0_filtered_output_c7(30);
   bh537_wm38_0_c7 <= tile_0_filtered_output_c7(31);
   bh537_wm37_0_c7 <= tile_0_filtered_output_c7(32);
   bh537_wm36_0_c7 <= tile_0_filtered_output_c7(33);
   bh537_wm35_0_c7 <= tile_0_filtered_output_c7(34);
   bh537_wm34_0_c7 <= tile_0_filtered_output_c7(35);
   bh537_wm33_0_c7 <= tile_0_filtered_output_c7(36);
   bh537_wm32_0_c7 <= tile_0_filtered_output_c7(37);
   bh537_wm31_0_c7 <= tile_0_filtered_output_c7(38);
   bh537_wm30_0_c7 <= tile_0_filtered_output_c7(39);
   bh537_wm29_0_c7 <= tile_0_filtered_output_c7(40);
   tile_1_X_c4 <= X(28 downto 17);
   tile_1_Y_c6 <= Y(23 downto 0);
   tile_1_mult: DSPBlock_12x24_Freq300_uid541
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 X => tile_1_X_c4,
                 Y => tile_1_Y_c6,
                 R => tile_1_output_c7);

   tile_1_filtered_output_c7 <= signed(tile_1_output_c7(35 downto 0));
   bh537_wm52_1_c7 <= tile_1_filtered_output_c7(0);
   bh537_wm51_1_c7 <= tile_1_filtered_output_c7(1);
   bh537_wm50_1_c7 <= tile_1_filtered_output_c7(2);
   bh537_wm49_1_c7 <= tile_1_filtered_output_c7(3);
   bh537_wm48_1_c7 <= tile_1_filtered_output_c7(4);
   bh537_wm47_1_c7 <= tile_1_filtered_output_c7(5);
   bh537_wm46_1_c7 <= tile_1_filtered_output_c7(6);
   bh537_wm45_1_c7 <= tile_1_filtered_output_c7(7);
   bh537_wm44_1_c7 <= tile_1_filtered_output_c7(8);
   bh537_wm43_1_c7 <= tile_1_filtered_output_c7(9);
   bh537_wm42_1_c7 <= tile_1_filtered_output_c7(10);
   bh537_wm41_1_c7 <= tile_1_filtered_output_c7(11);
   bh537_wm40_1_c7 <= tile_1_filtered_output_c7(12);
   bh537_wm39_1_c7 <= tile_1_filtered_output_c7(13);
   bh537_wm38_1_c7 <= tile_1_filtered_output_c7(14);
   bh537_wm37_1_c7 <= tile_1_filtered_output_c7(15);
   bh537_wm36_1_c7 <= tile_1_filtered_output_c7(16);
   bh537_wm35_1_c7 <= tile_1_filtered_output_c7(17);
   bh537_wm34_1_c7 <= tile_1_filtered_output_c7(18);
   bh537_wm33_1_c7 <= tile_1_filtered_output_c7(19);
   bh537_wm32_1_c7 <= tile_1_filtered_output_c7(20);
   bh537_wm31_1_c7 <= tile_1_filtered_output_c7(21);
   bh537_wm30_1_c7 <= tile_1_filtered_output_c7(22);
   bh537_wm29_1_c7 <= tile_1_filtered_output_c7(23);
   bh537_wm28_0_c7 <= tile_1_filtered_output_c7(24);
   bh537_wm27_0_c7 <= tile_1_filtered_output_c7(25);
   bh537_wm26_0_c7 <= tile_1_filtered_output_c7(26);
   bh537_wm25_0_c7 <= tile_1_filtered_output_c7(27);
   bh537_wm24_0_c7 <= tile_1_filtered_output_c7(28);
   bh537_wm23_0_c7 <= tile_1_filtered_output_c7(29);
   bh537_wm22_0_c7 <= tile_1_filtered_output_c7(30);
   bh537_wm21_0_c7 <= tile_1_filtered_output_c7(31);
   bh537_wm20_0_c7 <= tile_1_filtered_output_c7(32);
   bh537_wm19_0_c7 <= tile_1_filtered_output_c7(33);
   bh537_wm18_0_c7 <= tile_1_filtered_output_c7(34);
   bh537_wm17_0_c7 <= not tile_1_filtered_output_c7(35);
   tile_2_X_c4 <= X(16 downto 16);
   tile_2_Y_c6 <= Y(32 downto 32);
   tile_2_mult: IntMultiplierLUT_1x1_signed_Freq300_uid543
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_2_X_c4,
                 Y => tile_2_Y_c6,
                 R => tile_2_output_c6);

   tile_2_filtered_output_c6 <= signed(tile_2_output_c6(0 downto 0));
   bh537_wm21_1_c6 <= not tile_2_filtered_output_c6(0);
   tile_3_X_c4 <= X(15 downto 12);
   tile_3_Y_c6 <= Y(32 downto 32);
   tile_3_mult: IntMultiplierLUT_4x1_signed_Freq300_uid545
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_3_X_c4,
                 Y => tile_3_Y_c6,
                 R => tile_3_output_c6);

   tile_3_filtered_output_c6 <= signed(tile_3_output_c6(4 downto 0));
   bh537_wm25_1_c6 <= tile_3_filtered_output_c6(0);
   bh537_wm24_1_c6 <= tile_3_filtered_output_c6(1);
   bh537_wm23_1_c6 <= tile_3_filtered_output_c6(2);
   bh537_wm22_1_c6 <= tile_3_filtered_output_c6(3);
   bh537_wm21_2_c6 <= not tile_3_filtered_output_c6(4);
   tile_4_X_c4 <= X(11 downto 8);
   tile_4_Y_c6 <= Y(32 downto 32);
   tile_4_mult: IntMultiplierLUT_4x1_signed_Freq300_uid550
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_4_X_c4,
                 Y => tile_4_Y_c6,
                 R => tile_4_output_c6);

   tile_4_filtered_output_c6 <= signed(tile_4_output_c6(4 downto 0));
   bh537_wm29_2_c6 <= tile_4_filtered_output_c6(0);
   bh537_wm28_1_c6 <= tile_4_filtered_output_c6(1);
   bh537_wm27_1_c6 <= tile_4_filtered_output_c6(2);
   bh537_wm26_1_c6 <= tile_4_filtered_output_c6(3);
   bh537_wm25_2_c6 <= not tile_4_filtered_output_c6(4);
   tile_5_X_c4 <= X(7 downto 4);
   tile_5_Y_c6 <= Y(32 downto 32);
   tile_5_mult: IntMultiplierLUT_4x1_signed_Freq300_uid555
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_5_X_c4,
                 Y => tile_5_Y_c6,
                 R => tile_5_output_c6);

   tile_5_filtered_output_c6 <= signed(tile_5_output_c6(4 downto 0));
   bh537_wm33_2_c6 <= tile_5_filtered_output_c6(0);
   bh537_wm32_2_c6 <= tile_5_filtered_output_c6(1);
   bh537_wm31_2_c6 <= tile_5_filtered_output_c6(2);
   bh537_wm30_2_c6 <= tile_5_filtered_output_c6(3);
   bh537_wm29_3_c6 <= not tile_5_filtered_output_c6(4);
   tile_6_X_c4 <= X(3 downto 0);
   tile_6_Y_c6 <= Y(32 downto 32);
   tile_6_mult: IntMultiplierLUT_4x1_signed_Freq300_uid560
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_6_X_c4,
                 Y => tile_6_Y_c6,
                 R => tile_6_output_c6);

   tile_6_filtered_output_c6 <= signed(tile_6_output_c6(4 downto 0));
   bh537_wm37_2_c6 <= tile_6_filtered_output_c6(0);
   bh537_wm36_2_c6 <= tile_6_filtered_output_c6(1);
   bh537_wm35_2_c6 <= tile_6_filtered_output_c6(2);
   bh537_wm34_2_c6 <= tile_6_filtered_output_c6(3);
   bh537_wm33_3_c6 <= not tile_6_filtered_output_c6(4);
   tile_7_X_c4 <= X(16 downto 15);
   tile_7_Y_c6 <= Y(31 downto 30);
   tile_7_mult: IntMultiplierLUT_2x2_Freq300_uid565
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_7_X_c4,
                 Y => tile_7_Y_c6,
                 R => tile_7_output_c6);

   tile_7_filtered_output_c6 <= unsigned(tile_7_output_c6(3 downto 0));
   bh537_wm24_2_c6 <= tile_7_filtered_output_c6(0);
   bh537_wm23_2_c6 <= tile_7_filtered_output_c6(1);
   bh537_wm22_2_c6 <= tile_7_filtered_output_c6(2);
   bh537_wm21_3_c6 <= tile_7_filtered_output_c6(3);
   tile_8_X_c4 <= X(14 downto 12);
   tile_8_Y_c6 <= Y(31 downto 30);
   tile_8_mult: IntMultiplierLUT_3x2_Freq300_uid570
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_8_X_c4,
                 Y => tile_8_Y_c6,
                 R => tile_8_output_c6);

   tile_8_filtered_output_c6 <= unsigned(tile_8_output_c6(4 downto 0));
   bh537_wm27_2_c6 <= tile_8_filtered_output_c6(0);
   bh537_wm26_2_c6 <= tile_8_filtered_output_c6(1);
   bh537_wm25_3_c6 <= tile_8_filtered_output_c6(2);
   bh537_wm24_3_c6 <= tile_8_filtered_output_c6(3);
   bh537_wm23_3_c6 <= tile_8_filtered_output_c6(4);
   tile_9_X_c4 <= X(11 downto 9);
   tile_9_Y_c6 <= Y(31 downto 30);
   tile_9_mult: IntMultiplierLUT_3x2_Freq300_uid575
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_9_X_c4,
                 Y => tile_9_Y_c6,
                 R => tile_9_output_c6);

   tile_9_filtered_output_c6 <= unsigned(tile_9_output_c6(4 downto 0));
   bh537_wm30_3_c6 <= tile_9_filtered_output_c6(0);
   bh537_wm29_4_c6 <= tile_9_filtered_output_c6(1);
   bh537_wm28_2_c6 <= tile_9_filtered_output_c6(2);
   bh537_wm27_3_c6 <= tile_9_filtered_output_c6(3);
   bh537_wm26_3_c6 <= tile_9_filtered_output_c6(4);
   tile_10_X_c4 <= X(8 downto 6);
   tile_10_Y_c6 <= Y(31 downto 30);
   tile_10_mult: IntMultiplierLUT_3x2_Freq300_uid580
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_10_X_c4,
                 Y => tile_10_Y_c6,
                 R => tile_10_output_c6);

   tile_10_filtered_output_c6 <= unsigned(tile_10_output_c6(4 downto 0));
   bh537_wm33_4_c6 <= tile_10_filtered_output_c6(0);
   bh537_wm32_3_c6 <= tile_10_filtered_output_c6(1);
   bh537_wm31_3_c6 <= tile_10_filtered_output_c6(2);
   bh537_wm30_4_c6 <= tile_10_filtered_output_c6(3);
   bh537_wm29_5_c6 <= tile_10_filtered_output_c6(4);
   tile_11_X_c4 <= X(5 downto 3);
   tile_11_Y_c6 <= Y(31 downto 30);
   tile_11_mult: IntMultiplierLUT_3x2_Freq300_uid585
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_11_X_c4,
                 Y => tile_11_Y_c6,
                 R => tile_11_output_c6);

   tile_11_filtered_output_c6 <= unsigned(tile_11_output_c6(4 downto 0));
   bh537_wm36_3_c6 <= tile_11_filtered_output_c6(0);
   bh537_wm35_3_c6 <= tile_11_filtered_output_c6(1);
   bh537_wm34_3_c6 <= tile_11_filtered_output_c6(2);
   bh537_wm33_5_c6 <= tile_11_filtered_output_c6(3);
   bh537_wm32_4_c6 <= tile_11_filtered_output_c6(4);
   tile_12_X_c4 <= X(2 downto 0);
   tile_12_Y_c6 <= Y(31 downto 30);
   tile_12_mult: IntMultiplierLUT_3x2_Freq300_uid590
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_12_X_c4,
                 Y => tile_12_Y_c6,
                 R => tile_12_output_c6);

   tile_12_filtered_output_c6 <= unsigned(tile_12_output_c6(4 downto 0));
   bh537_wm39_2_c6 <= tile_12_filtered_output_c6(0);
   bh537_wm38_2_c6 <= tile_12_filtered_output_c6(1);
   bh537_wm37_3_c6 <= tile_12_filtered_output_c6(2);
   bh537_wm36_4_c6 <= tile_12_filtered_output_c6(3);
   bh537_wm35_4_c6 <= tile_12_filtered_output_c6(4);
   tile_13_X_c4 <= X(16 downto 15);
   tile_13_Y_c6 <= Y(29 downto 28);
   tile_13_mult: IntMultiplierLUT_2x2_Freq300_uid595
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_13_X_c4,
                 Y => tile_13_Y_c6,
                 R => tile_13_output_c6);

   tile_13_filtered_output_c6 <= unsigned(tile_13_output_c6(3 downto 0));
   bh537_wm26_4_c6 <= tile_13_filtered_output_c6(0);
   bh537_wm25_4_c6 <= tile_13_filtered_output_c6(1);
   bh537_wm24_4_c6 <= tile_13_filtered_output_c6(2);
   bh537_wm23_4_c6 <= tile_13_filtered_output_c6(3);
   tile_14_X_c4 <= X(14 downto 12);
   tile_14_Y_c6 <= Y(29 downto 28);
   tile_14_mult: IntMultiplierLUT_3x2_Freq300_uid600
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_14_X_c4,
                 Y => tile_14_Y_c6,
                 R => tile_14_output_c6);

   tile_14_filtered_output_c6 <= unsigned(tile_14_output_c6(4 downto 0));
   bh537_wm29_6_c6 <= tile_14_filtered_output_c6(0);
   bh537_wm28_3_c6 <= tile_14_filtered_output_c6(1);
   bh537_wm27_4_c6 <= tile_14_filtered_output_c6(2);
   bh537_wm26_5_c6 <= tile_14_filtered_output_c6(3);
   bh537_wm25_5_c6 <= tile_14_filtered_output_c6(4);
   tile_15_X_c4 <= X(11 downto 9);
   tile_15_Y_c6 <= Y(29 downto 28);
   tile_15_mult: IntMultiplierLUT_3x2_Freq300_uid605
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_15_X_c4,
                 Y => tile_15_Y_c6,
                 R => tile_15_output_c6);

   tile_15_filtered_output_c6 <= unsigned(tile_15_output_c6(4 downto 0));
   bh537_wm32_5_c6 <= tile_15_filtered_output_c6(0);
   bh537_wm31_4_c6 <= tile_15_filtered_output_c6(1);
   bh537_wm30_5_c6 <= tile_15_filtered_output_c6(2);
   bh537_wm29_7_c6 <= tile_15_filtered_output_c6(3);
   bh537_wm28_4_c6 <= tile_15_filtered_output_c6(4);
   tile_16_X_c4 <= X(8 downto 6);
   tile_16_Y_c6 <= Y(29 downto 28);
   tile_16_mult: IntMultiplierLUT_3x2_Freq300_uid610
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_16_X_c4,
                 Y => tile_16_Y_c6,
                 R => tile_16_output_c6);

   tile_16_filtered_output_c6 <= unsigned(tile_16_output_c6(4 downto 0));
   bh537_wm35_5_c6 <= tile_16_filtered_output_c6(0);
   bh537_wm34_4_c6 <= tile_16_filtered_output_c6(1);
   bh537_wm33_6_c6 <= tile_16_filtered_output_c6(2);
   bh537_wm32_6_c6 <= tile_16_filtered_output_c6(3);
   bh537_wm31_5_c6 <= tile_16_filtered_output_c6(4);
   tile_17_X_c4 <= X(5 downto 3);
   tile_17_Y_c6 <= Y(29 downto 28);
   tile_17_mult: IntMultiplierLUT_3x2_Freq300_uid615
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_17_X_c4,
                 Y => tile_17_Y_c6,
                 R => tile_17_output_c6);

   tile_17_filtered_output_c6 <= unsigned(tile_17_output_c6(4 downto 0));
   bh537_wm38_3_c6 <= tile_17_filtered_output_c6(0);
   bh537_wm37_4_c6 <= tile_17_filtered_output_c6(1);
   bh537_wm36_5_c6 <= tile_17_filtered_output_c6(2);
   bh537_wm35_6_c6 <= tile_17_filtered_output_c6(3);
   bh537_wm34_5_c6 <= tile_17_filtered_output_c6(4);
   tile_18_X_c4 <= X(2 downto 0);
   tile_18_Y_c6 <= Y(29 downto 28);
   tile_18_mult: IntMultiplierLUT_3x2_Freq300_uid620
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_18_X_c4,
                 Y => tile_18_Y_c6,
                 R => tile_18_output_c6);

   tile_18_filtered_output_c6 <= unsigned(tile_18_output_c6(4 downto 0));
   bh537_wm41_2_c6 <= tile_18_filtered_output_c6(0);
   bh537_wm40_2_c6 <= tile_18_filtered_output_c6(1);
   bh537_wm39_3_c6 <= tile_18_filtered_output_c6(2);
   bh537_wm38_4_c6 <= tile_18_filtered_output_c6(3);
   bh537_wm37_5_c6 <= tile_18_filtered_output_c6(4);
   tile_19_X_c4 <= X(16 downto 15);
   tile_19_Y_c6 <= Y(27 downto 26);
   tile_19_mult: IntMultiplierLUT_2x2_Freq300_uid625
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_19_X_c4,
                 Y => tile_19_Y_c6,
                 R => tile_19_output_c6);

   tile_19_filtered_output_c6 <= unsigned(tile_19_output_c6(3 downto 0));
   bh537_wm28_5_c6 <= tile_19_filtered_output_c6(0);
   bh537_wm27_5_c6 <= tile_19_filtered_output_c6(1);
   bh537_wm26_6_c6 <= tile_19_filtered_output_c6(2);
   bh537_wm25_6_c6 <= tile_19_filtered_output_c6(3);
   tile_20_X_c4 <= X(14 downto 12);
   tile_20_Y_c6 <= Y(27 downto 26);
   tile_20_mult: IntMultiplierLUT_3x2_Freq300_uid630
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_20_X_c4,
                 Y => tile_20_Y_c6,
                 R => tile_20_output_c6);

   tile_20_filtered_output_c6 <= unsigned(tile_20_output_c6(4 downto 0));
   bh537_wm31_6_c6 <= tile_20_filtered_output_c6(0);
   bh537_wm30_6_c6 <= tile_20_filtered_output_c6(1);
   bh537_wm29_8_c6 <= tile_20_filtered_output_c6(2);
   bh537_wm28_6_c6 <= tile_20_filtered_output_c6(3);
   bh537_wm27_6_c6 <= tile_20_filtered_output_c6(4);
   tile_21_X_c4 <= X(11 downto 9);
   tile_21_Y_c6 <= Y(27 downto 26);
   tile_21_mult: IntMultiplierLUT_3x2_Freq300_uid635
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_21_X_c4,
                 Y => tile_21_Y_c6,
                 R => tile_21_output_c6);

   tile_21_filtered_output_c6 <= unsigned(tile_21_output_c6(4 downto 0));
   bh537_wm34_6_c6 <= tile_21_filtered_output_c6(0);
   bh537_wm33_7_c6 <= tile_21_filtered_output_c6(1);
   bh537_wm32_7_c6 <= tile_21_filtered_output_c6(2);
   bh537_wm31_7_c6 <= tile_21_filtered_output_c6(3);
   bh537_wm30_7_c6 <= tile_21_filtered_output_c6(4);
   tile_22_X_c4 <= X(8 downto 6);
   tile_22_Y_c6 <= Y(27 downto 26);
   tile_22_mult: IntMultiplierLUT_3x2_Freq300_uid640
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_22_X_c4,
                 Y => tile_22_Y_c6,
                 R => tile_22_output_c6);

   tile_22_filtered_output_c6 <= unsigned(tile_22_output_c6(4 downto 0));
   bh537_wm37_6_c6 <= tile_22_filtered_output_c6(0);
   bh537_wm36_6_c6 <= tile_22_filtered_output_c6(1);
   bh537_wm35_7_c6 <= tile_22_filtered_output_c6(2);
   bh537_wm34_7_c6 <= tile_22_filtered_output_c6(3);
   bh537_wm33_8_c6 <= tile_22_filtered_output_c6(4);
   tile_23_X_c4 <= X(5 downto 3);
   tile_23_Y_c6 <= Y(27 downto 26);
   tile_23_mult: IntMultiplierLUT_3x2_Freq300_uid645
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_23_X_c4,
                 Y => tile_23_Y_c6,
                 R => tile_23_output_c6);

   tile_23_filtered_output_c6 <= unsigned(tile_23_output_c6(4 downto 0));
   bh537_wm40_3_c6 <= tile_23_filtered_output_c6(0);
   bh537_wm39_4_c6 <= tile_23_filtered_output_c6(1);
   bh537_wm38_5_c6 <= tile_23_filtered_output_c6(2);
   bh537_wm37_7_c6 <= tile_23_filtered_output_c6(3);
   bh537_wm36_7_c6 <= tile_23_filtered_output_c6(4);
   tile_24_X_c4 <= X(2 downto 0);
   tile_24_Y_c6 <= Y(27 downto 26);
   tile_24_mult: IntMultiplierLUT_3x2_Freq300_uid650
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_24_X_c4,
                 Y => tile_24_Y_c6,
                 R => tile_24_output_c6);

   tile_24_filtered_output_c6 <= unsigned(tile_24_output_c6(4 downto 0));
   bh537_wm43_2_c6 <= tile_24_filtered_output_c6(0);
   bh537_wm42_2_c6 <= tile_24_filtered_output_c6(1);
   bh537_wm41_3_c6 <= tile_24_filtered_output_c6(2);
   bh537_wm40_4_c6 <= tile_24_filtered_output_c6(3);
   bh537_wm39_5_c6 <= tile_24_filtered_output_c6(4);
   tile_25_X_c4 <= X(16 downto 15);
   tile_25_Y_c6 <= Y(25 downto 24);
   tile_25_mult: IntMultiplierLUT_2x2_Freq300_uid655
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_25_X_c4,
                 Y => tile_25_Y_c6,
                 R => tile_25_output_c6);

   tile_25_filtered_output_c6 <= unsigned(tile_25_output_c6(3 downto 0));
   bh537_wm30_8_c6 <= tile_25_filtered_output_c6(0);
   bh537_wm29_9_c6 <= tile_25_filtered_output_c6(1);
   bh537_wm28_7_c6 <= tile_25_filtered_output_c6(2);
   bh537_wm27_7_c6 <= tile_25_filtered_output_c6(3);
   tile_26_X_c4 <= X(14 downto 12);
   tile_26_Y_c6 <= Y(25 downto 24);
   tile_26_mult: IntMultiplierLUT_3x2_Freq300_uid660
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_26_X_c4,
                 Y => tile_26_Y_c6,
                 R => tile_26_output_c6);

   tile_26_filtered_output_c6 <= unsigned(tile_26_output_c6(4 downto 0));
   bh537_wm33_9_c6 <= tile_26_filtered_output_c6(0);
   bh537_wm32_8_c6 <= tile_26_filtered_output_c6(1);
   bh537_wm31_8_c6 <= tile_26_filtered_output_c6(2);
   bh537_wm30_9_c6 <= tile_26_filtered_output_c6(3);
   bh537_wm29_10_c6 <= tile_26_filtered_output_c6(4);
   tile_27_X_c4 <= X(11 downto 9);
   tile_27_Y_c6 <= Y(25 downto 24);
   tile_27_mult: IntMultiplierLUT_3x2_Freq300_uid665
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_27_X_c4,
                 Y => tile_27_Y_c6,
                 R => tile_27_output_c6);

   tile_27_filtered_output_c6 <= unsigned(tile_27_output_c6(4 downto 0));
   bh537_wm36_8_c6 <= tile_27_filtered_output_c6(0);
   bh537_wm35_8_c6 <= tile_27_filtered_output_c6(1);
   bh537_wm34_8_c6 <= tile_27_filtered_output_c6(2);
   bh537_wm33_10_c6 <= tile_27_filtered_output_c6(3);
   bh537_wm32_9_c6 <= tile_27_filtered_output_c6(4);
   tile_28_X_c4 <= X(8 downto 6);
   tile_28_Y_c6 <= Y(25 downto 24);
   tile_28_mult: IntMultiplierLUT_3x2_Freq300_uid670
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_28_X_c4,
                 Y => tile_28_Y_c6,
                 R => tile_28_output_c6);

   tile_28_filtered_output_c6 <= unsigned(tile_28_output_c6(4 downto 0));
   bh537_wm39_6_c6 <= tile_28_filtered_output_c6(0);
   bh537_wm38_6_c6 <= tile_28_filtered_output_c6(1);
   bh537_wm37_8_c6 <= tile_28_filtered_output_c6(2);
   bh537_wm36_9_c6 <= tile_28_filtered_output_c6(3);
   bh537_wm35_9_c6 <= tile_28_filtered_output_c6(4);
   tile_29_X_c4 <= X(5 downto 3);
   tile_29_Y_c6 <= Y(25 downto 24);
   tile_29_mult: IntMultiplierLUT_3x2_Freq300_uid675
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_29_X_c4,
                 Y => tile_29_Y_c6,
                 R => tile_29_output_c6);

   tile_29_filtered_output_c6 <= unsigned(tile_29_output_c6(4 downto 0));
   bh537_wm42_3_c6 <= tile_29_filtered_output_c6(0);
   bh537_wm41_4_c6 <= tile_29_filtered_output_c6(1);
   bh537_wm40_5_c6 <= tile_29_filtered_output_c6(2);
   bh537_wm39_7_c6 <= tile_29_filtered_output_c6(3);
   bh537_wm38_7_c6 <= tile_29_filtered_output_c6(4);
   tile_30_X_c4 <= X(2 downto 0);
   tile_30_Y_c6 <= Y(25 downto 24);
   tile_30_mult: IntMultiplierLUT_3x2_Freq300_uid680
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_30_X_c4,
                 Y => tile_30_Y_c6,
                 R => tile_30_output_c6);

   tile_30_filtered_output_c6 <= unsigned(tile_30_output_c6(4 downto 0));
   bh537_wm45_2_c6 <= tile_30_filtered_output_c6(0);
   bh537_wm44_2_c6 <= tile_30_filtered_output_c6(1);
   bh537_wm43_3_c6 <= tile_30_filtered_output_c6(2);
   bh537_wm42_4_c6 <= tile_30_filtered_output_c6(3);
   bh537_wm41_5_c6 <= tile_30_filtered_output_c6(4);
   tile_31_X_c4 <= X(28 downto 25);
   tile_31_Y_c6 <= Y(32 downto 32);
   tile_31_mult: IntMultiplierLUT_4_signedx1_signed_Freq300_uid685
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_31_X_c4,
                 Y => tile_31_Y_c6,
                 R => tile_31_output_c6);

   tile_31_filtered_output_c6 <= signed(tile_31_output_c6(4 downto 0));
   bh537_wm12_0_c6 <= tile_31_filtered_output_c6(0);
   bh537_wm11_0_c6 <= tile_31_filtered_output_c6(1);
   bh537_wm10_0_c6 <= tile_31_filtered_output_c6(2);
   bh537_wm9_0_c6 <= tile_31_filtered_output_c6(3);
   bh537_wm8_0_c6 <= not tile_31_filtered_output_c6(4);
   tile_32_X_c4 <= X(24 downto 21);
   tile_32_Y_c6 <= Y(32 downto 32);
   tile_32_mult: IntMultiplierLUT_4x1_signed_Freq300_uid690
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_32_X_c4,
                 Y => tile_32_Y_c6,
                 R => tile_32_output_c6);

   tile_32_filtered_output_c6 <= signed(tile_32_output_c6(4 downto 0));
   bh537_wm16_0_c6 <= tile_32_filtered_output_c6(0);
   bh537_wm15_0_c6 <= tile_32_filtered_output_c6(1);
   bh537_wm14_0_c6 <= tile_32_filtered_output_c6(2);
   bh537_wm13_0_c6 <= tile_32_filtered_output_c6(3);
   bh537_wm12_1_c6 <= not tile_32_filtered_output_c6(4);
   tile_33_X_c4 <= X(20 downto 17);
   tile_33_Y_c6 <= Y(32 downto 32);
   tile_33_mult: IntMultiplierLUT_4x1_signed_Freq300_uid695
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_33_X_c4,
                 Y => tile_33_Y_c6,
                 R => tile_33_output_c6);

   tile_33_filtered_output_c6 <= signed(tile_33_output_c6(4 downto 0));
   bh537_wm20_1_c6 <= tile_33_filtered_output_c6(0);
   bh537_wm19_1_c6 <= tile_33_filtered_output_c6(1);
   bh537_wm18_1_c6 <= tile_33_filtered_output_c6(2);
   bh537_wm17_1_c6 <= tile_33_filtered_output_c6(3);
   bh537_wm16_1_c6 <= not tile_33_filtered_output_c6(4);
   tile_34_X_c4 <= X(28 downto 26);
   tile_34_Y_c6 <= Y(31 downto 30);
   tile_34_mult: IntMultiplierLUT_3_signedx2_Freq300_uid700
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_34_X_c4,
                 Y => tile_34_Y_c6,
                 R => tile_34_output_c6);

   tile_34_filtered_output_c6 <= signed(tile_34_output_c6(4 downto 0));
   bh537_wm13_1_c6 <= tile_34_filtered_output_c6(0);
   bh537_wm12_2_c6 <= tile_34_filtered_output_c6(1);
   bh537_wm11_1_c6 <= tile_34_filtered_output_c6(2);
   bh537_wm10_1_c6 <= tile_34_filtered_output_c6(3);
   bh537_wm9_1_c6 <= not tile_34_filtered_output_c6(4);
   tile_35_X_c4 <= X(25 downto 23);
   tile_35_Y_c6 <= Y(31 downto 30);
   tile_35_mult: IntMultiplierLUT_3x2_Freq300_uid705
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_35_X_c4,
                 Y => tile_35_Y_c6,
                 R => tile_35_output_c6);

   tile_35_filtered_output_c6 <= unsigned(tile_35_output_c6(4 downto 0));
   bh537_wm16_2_c6 <= tile_35_filtered_output_c6(0);
   bh537_wm15_1_c6 <= tile_35_filtered_output_c6(1);
   bh537_wm14_1_c6 <= tile_35_filtered_output_c6(2);
   bh537_wm13_2_c6 <= tile_35_filtered_output_c6(3);
   bh537_wm12_3_c6 <= tile_35_filtered_output_c6(4);
   tile_36_X_c4 <= X(22 downto 20);
   tile_36_Y_c6 <= Y(31 downto 30);
   tile_36_mult: IntMultiplierLUT_3x2_Freq300_uid710
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_36_X_c4,
                 Y => tile_36_Y_c6,
                 R => tile_36_output_c6);

   tile_36_filtered_output_c6 <= unsigned(tile_36_output_c6(4 downto 0));
   bh537_wm19_2_c6 <= tile_36_filtered_output_c6(0);
   bh537_wm18_2_c6 <= tile_36_filtered_output_c6(1);
   bh537_wm17_2_c6 <= tile_36_filtered_output_c6(2);
   bh537_wm16_3_c6 <= tile_36_filtered_output_c6(3);
   bh537_wm15_2_c6 <= tile_36_filtered_output_c6(4);
   tile_37_X_c4 <= X(19 downto 17);
   tile_37_Y_c6 <= Y(31 downto 30);
   tile_37_mult: IntMultiplierLUT_3x2_Freq300_uid715
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_37_X_c4,
                 Y => tile_37_Y_c6,
                 R => tile_37_output_c6);

   tile_37_filtered_output_c6 <= unsigned(tile_37_output_c6(4 downto 0));
   bh537_wm22_3_c6 <= tile_37_filtered_output_c6(0);
   bh537_wm21_4_c6 <= tile_37_filtered_output_c6(1);
   bh537_wm20_2_c6 <= tile_37_filtered_output_c6(2);
   bh537_wm19_3_c6 <= tile_37_filtered_output_c6(3);
   bh537_wm18_3_c6 <= tile_37_filtered_output_c6(4);
   tile_38_X_c4 <= X(28 downto 26);
   tile_38_Y_c6 <= Y(29 downto 28);
   tile_38_mult: IntMultiplierLUT_3_signedx2_Freq300_uid720
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_38_X_c4,
                 Y => tile_38_Y_c6,
                 R => tile_38_output_c6);

   tile_38_filtered_output_c6 <= signed(tile_38_output_c6(4 downto 0));
   bh537_wm15_3_c6 <= tile_38_filtered_output_c6(0);
   bh537_wm14_2_c6 <= tile_38_filtered_output_c6(1);
   bh537_wm13_3_c6 <= tile_38_filtered_output_c6(2);
   bh537_wm12_4_c6 <= tile_38_filtered_output_c6(3);
   bh537_wm11_2_c6 <= not tile_38_filtered_output_c6(4);
   tile_39_X_c4 <= X(25 downto 23);
   tile_39_Y_c6 <= Y(29 downto 28);
   tile_39_mult: IntMultiplierLUT_3x2_Freq300_uid725
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_39_X_c4,
                 Y => tile_39_Y_c6,
                 R => tile_39_output_c6);

   tile_39_filtered_output_c6 <= unsigned(tile_39_output_c6(4 downto 0));
   bh537_wm18_4_c6 <= tile_39_filtered_output_c6(0);
   bh537_wm17_3_c6 <= tile_39_filtered_output_c6(1);
   bh537_wm16_4_c6 <= tile_39_filtered_output_c6(2);
   bh537_wm15_4_c6 <= tile_39_filtered_output_c6(3);
   bh537_wm14_3_c6 <= tile_39_filtered_output_c6(4);
   tile_40_X_c4 <= X(22 downto 20);
   tile_40_Y_c6 <= Y(29 downto 28);
   tile_40_mult: IntMultiplierLUT_3x2_Freq300_uid730
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_40_X_c4,
                 Y => tile_40_Y_c6,
                 R => tile_40_output_c6);

   tile_40_filtered_output_c6 <= unsigned(tile_40_output_c6(4 downto 0));
   bh537_wm21_5_c6 <= tile_40_filtered_output_c6(0);
   bh537_wm20_3_c6 <= tile_40_filtered_output_c6(1);
   bh537_wm19_4_c6 <= tile_40_filtered_output_c6(2);
   bh537_wm18_5_c6 <= tile_40_filtered_output_c6(3);
   bh537_wm17_4_c6 <= tile_40_filtered_output_c6(4);
   tile_41_X_c4 <= X(19 downto 17);
   tile_41_Y_c6 <= Y(29 downto 28);
   tile_41_mult: IntMultiplierLUT_3x2_Freq300_uid735
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_41_X_c4,
                 Y => tile_41_Y_c6,
                 R => tile_41_output_c6);

   tile_41_filtered_output_c6 <= unsigned(tile_41_output_c6(4 downto 0));
   bh537_wm24_5_c6 <= tile_41_filtered_output_c6(0);
   bh537_wm23_5_c6 <= tile_41_filtered_output_c6(1);
   bh537_wm22_4_c6 <= tile_41_filtered_output_c6(2);
   bh537_wm21_6_c6 <= tile_41_filtered_output_c6(3);
   bh537_wm20_4_c6 <= tile_41_filtered_output_c6(4);
   tile_42_X_c4 <= X(28 downto 26);
   tile_42_Y_c6 <= Y(27 downto 26);
   tile_42_mult: IntMultiplierLUT_3_signedx2_Freq300_uid740
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_42_X_c4,
                 Y => tile_42_Y_c6,
                 R => tile_42_output_c6);

   tile_42_filtered_output_c6 <= signed(tile_42_output_c6(4 downto 0));
   bh537_wm17_5_c6 <= tile_42_filtered_output_c6(0);
   bh537_wm16_5_c6 <= tile_42_filtered_output_c6(1);
   bh537_wm15_5_c6 <= tile_42_filtered_output_c6(2);
   bh537_wm14_4_c6 <= tile_42_filtered_output_c6(3);
   bh537_wm13_4_c6 <= not tile_42_filtered_output_c6(4);
   tile_43_X_c4 <= X(25 downto 23);
   tile_43_Y_c6 <= Y(27 downto 26);
   tile_43_mult: IntMultiplierLUT_3x2_Freq300_uid745
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_43_X_c4,
                 Y => tile_43_Y_c6,
                 R => tile_43_output_c6);

   tile_43_filtered_output_c6 <= unsigned(tile_43_output_c6(4 downto 0));
   bh537_wm20_5_c6 <= tile_43_filtered_output_c6(0);
   bh537_wm19_5_c6 <= tile_43_filtered_output_c6(1);
   bh537_wm18_6_c6 <= tile_43_filtered_output_c6(2);
   bh537_wm17_6_c6 <= tile_43_filtered_output_c6(3);
   bh537_wm16_6_c6 <= tile_43_filtered_output_c6(4);
   tile_44_X_c4 <= X(22 downto 20);
   tile_44_Y_c6 <= Y(27 downto 26);
   tile_44_mult: IntMultiplierLUT_3x2_Freq300_uid750
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_44_X_c4,
                 Y => tile_44_Y_c6,
                 R => tile_44_output_c6);

   tile_44_filtered_output_c6 <= unsigned(tile_44_output_c6(4 downto 0));
   bh537_wm23_6_c6 <= tile_44_filtered_output_c6(0);
   bh537_wm22_5_c6 <= tile_44_filtered_output_c6(1);
   bh537_wm21_7_c6 <= tile_44_filtered_output_c6(2);
   bh537_wm20_6_c6 <= tile_44_filtered_output_c6(3);
   bh537_wm19_6_c6 <= tile_44_filtered_output_c6(4);
   tile_45_X_c4 <= X(19 downto 17);
   tile_45_Y_c6 <= Y(27 downto 26);
   tile_45_mult: IntMultiplierLUT_3x2_Freq300_uid755
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_45_X_c4,
                 Y => tile_45_Y_c6,
                 R => tile_45_output_c6);

   tile_45_filtered_output_c6 <= unsigned(tile_45_output_c6(4 downto 0));
   bh537_wm26_7_c6 <= tile_45_filtered_output_c6(0);
   bh537_wm25_7_c6 <= tile_45_filtered_output_c6(1);
   bh537_wm24_6_c6 <= tile_45_filtered_output_c6(2);
   bh537_wm23_7_c6 <= tile_45_filtered_output_c6(3);
   bh537_wm22_6_c6 <= tile_45_filtered_output_c6(4);
   tile_46_X_c4 <= X(28 downto 26);
   tile_46_Y_c6 <= Y(25 downto 24);
   tile_46_mult: IntMultiplierLUT_3_signedx2_Freq300_uid760
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_46_X_c4,
                 Y => tile_46_Y_c6,
                 R => tile_46_output_c6);

   tile_46_filtered_output_c6 <= signed(tile_46_output_c6(4 downto 0));
   bh537_wm19_7_c6 <= tile_46_filtered_output_c6(0);
   bh537_wm18_7_c6 <= tile_46_filtered_output_c6(1);
   bh537_wm17_7_c6 <= tile_46_filtered_output_c6(2);
   bh537_wm16_7_c6 <= tile_46_filtered_output_c6(3);
   bh537_wm15_6_c6 <= not tile_46_filtered_output_c6(4);
   tile_47_X_c4 <= X(25 downto 23);
   tile_47_Y_c6 <= Y(25 downto 24);
   tile_47_mult: IntMultiplierLUT_3x2_Freq300_uid765
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_47_X_c4,
                 Y => tile_47_Y_c6,
                 R => tile_47_output_c6);

   tile_47_filtered_output_c6 <= unsigned(tile_47_output_c6(4 downto 0));
   bh537_wm22_7_c6 <= tile_47_filtered_output_c6(0);
   bh537_wm21_8_c6 <= tile_47_filtered_output_c6(1);
   bh537_wm20_7_c6 <= tile_47_filtered_output_c6(2);
   bh537_wm19_8_c6 <= tile_47_filtered_output_c6(3);
   bh537_wm18_8_c6 <= tile_47_filtered_output_c6(4);
   tile_48_X_c4 <= X(22 downto 20);
   tile_48_Y_c6 <= Y(25 downto 24);
   tile_48_mult: IntMultiplierLUT_3x2_Freq300_uid770
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_48_X_c4,
                 Y => tile_48_Y_c6,
                 R => tile_48_output_c6);

   tile_48_filtered_output_c6 <= unsigned(tile_48_output_c6(4 downto 0));
   bh537_wm25_8_c6 <= tile_48_filtered_output_c6(0);
   bh537_wm24_7_c6 <= tile_48_filtered_output_c6(1);
   bh537_wm23_8_c6 <= tile_48_filtered_output_c6(2);
   bh537_wm22_8_c6 <= tile_48_filtered_output_c6(3);
   bh537_wm21_9_c6 <= tile_48_filtered_output_c6(4);
   tile_49_X_c4 <= X(19 downto 17);
   tile_49_Y_c6 <= Y(25 downto 24);
   tile_49_mult: IntMultiplierLUT_3x2_Freq300_uid775
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 X => tile_49_X_c4,
                 Y => tile_49_Y_c6,
                 R => tile_49_output_c6);

   tile_49_filtered_output_c6 <= unsigned(tile_49_output_c6(4 downto 0));
   bh537_wm28_8_c6 <= tile_49_filtered_output_c6(0);
   bh537_wm27_8_c6 <= tile_49_filtered_output_c6(1);
   bh537_wm26_8_c6 <= tile_49_filtered_output_c6(2);
   bh537_wm25_9_c6 <= tile_49_filtered_output_c6(3);
   bh537_wm24_8_c6 <= tile_49_filtered_output_c6(4);
   bh537_wm41_6_c4 <= AA_c4(0);
   bh537_wm40_6_c4 <= AA_c4(1);
   bh537_wm39_8_c4 <= AA_c4(2);
   bh537_wm38_8_c4 <= AA_c4(3);
   bh537_wm37_9_c4 <= AA_c4(4);
   bh537_wm36_10_c4 <= AA_c4(5);
   bh537_wm35_10_c4 <= AA_c4(6);
   bh537_wm34_9_c4 <= AA_c4(7);
   bh537_wm33_11_c4 <= AA_c4(8);
   bh537_wm32_10_c4 <= AA_c4(9);
   bh537_wm31_9_c4 <= AA_c4(10);
   bh537_wm30_10_c4 <= AA_c4(11);
   bh537_wm29_11_c4 <= AA_c4(12);
   bh537_wm28_9_c4 <= AA_c4(13);
   bh537_wm27_9_c4 <= AA_c4(14);
   bh537_wm26_9_c4 <= AA_c4(15);
   bh537_wm25_10_c4 <= AA_c4(16);
   bh537_wm24_9_c4 <= AA_c4(17);
   bh537_wm23_9_c4 <= AA_c4(18);
   bh537_wm22_9_c4 <= AA_c4(19);
   bh537_wm21_10_c4 <= AA_c4(20);
   bh537_wm20_8_c4 <= AA_c4(21);
   bh537_wm19_9_c4 <= AA_c4(22);
   bh537_wm18_9_c4 <= AA_c4(23);
   bh537_wm17_8_c4 <= AA_c4(24);
   bh537_wm16_8_c4 <= AA_c4(25);
   bh537_wm15_7_c4 <= AA_c4(26);
   bh537_wm14_5_c4 <= AA_c4(27);
   bh537_wm13_5_c4 <= AA_c4(28);
   bh537_wm12_5_c4 <= AA_c4(29);
   bh537_wm11_3_c4 <= AA_c4(30);
   bh537_wm10_2_c4 <= AA_c4(31);
   bh537_wm9_2_c4 <= AA_c4(32);
   bh537_wm8_1_c4 <= AA_c4(33);
   bh537_wm7_0_c4 <= AA_c4(34);
   bh537_wm6_0_c4 <= AA_c4(35);
   bh537_wm5_0_c4 <= AA_c4(36);
   bh537_wm4_0_c4 <= AA_c4(37);
   bh537_wm3_0_c4 <= AA_c4(38);
   bh537_wm2_0_c4 <= not AA_c4(39);

   -- Adding the constant bits 
   bh537_wm42_5_c0 <= '1';
   bh537_wm33_12_c0 <= '1';
   bh537_wm32_11_c0 <= '1';
   bh537_wm31_10_c0 <= '1';
   bh537_wm30_11_c0 <= '1';
   bh537_wm28_10_c0 <= '1';
   bh537_wm27_10_c0 <= '1';
   bh537_wm26_10_c0 <= '1';
   bh537_wm24_10_c0 <= '1';
   bh537_wm23_10_c0 <= '1';
   bh537_wm22_10_c0 <= '1';
   bh537_wm21_11_c0 <= '1';
   bh537_wm19_10_c0 <= '1';
   bh537_wm18_10_c0 <= '1';
   bh537_wm14_6_c0 <= '1';
   bh537_wm10_3_c0 <= '1';
   bh537_wm7_1_c0 <= '1';
   bh537_wm6_1_c0 <= '1';
   bh537_wm5_1_c0 <= '1';
   bh537_wm4_1_c0 <= '1';
   bh537_wm3_1_c0 <= '1';
   bh537_wm1_0_c0 <= '1';


   Compressor_23_3_Freq300_uid781_bh537_uid782_In0_c7 <= "" & bh537_wm52_0_c7 & bh537_wm52_1_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid782_In1_c7 <= "" & bh537_wm51_0_c7 & bh537_wm51_1_c7;
   bh537_wm52_2_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid782_Out0_c7(0);
   bh537_wm51_2_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid782_Out0_c7(1);
   bh537_wm50_2_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid782_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid782: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid782_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid782_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid782_Out0_copy783_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid782_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid782_Out0_copy783_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid784_In0_c7 <= "" & bh537_wm50_0_c7 & bh537_wm50_1_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid784_In1_c7 <= "" & bh537_wm49_0_c7 & bh537_wm49_1_c7;
   bh537_wm50_3_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid784_Out0_c7(0);
   bh537_wm49_2_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid784_Out0_c7(1);
   bh537_wm48_2_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid784_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid784: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid784_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid784_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid784_Out0_copy785_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid784_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid784_Out0_copy785_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid786_In0_c7 <= "" & bh537_wm48_0_c7 & bh537_wm48_1_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid786_In1_c7 <= "" & bh537_wm47_0_c7 & bh537_wm47_1_c7;
   bh537_wm48_3_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid786_Out0_c7(0);
   bh537_wm47_2_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid786_Out0_c7(1);
   bh537_wm46_2_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid786_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid786: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid786_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid786_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid786_Out0_copy787_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid786_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid786_Out0_copy787_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid790_In0_c7 <= "" & bh537_wm46_0_c7 & bh537_wm46_1_c7 & "0";
   bh537_wm46_3_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid790_Out0_c7(0);
   bh537_wm45_3_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid790_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid790: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid790_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid790_Out0_copy791_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid790_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid790_Out0_copy791_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid792_In0_c7 <= "" & bh537_wm45_0_c7 & bh537_wm45_1_c7 & bh537_wm45_2_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid792_In1_c7 <= "" & bh537_wm44_0_c7 & bh537_wm44_1_c7;
   bh537_wm45_4_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid792_Out0_c7(0);
   bh537_wm44_3_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid792_Out0_c7(1);
   bh537_wm43_4_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid792_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid792: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid792_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid792_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid792_Out0_copy793_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid792_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid792_Out0_copy793_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid794_In0_c7 <= "" & bh537_wm43_0_c7 & bh537_wm43_1_c7 & bh537_wm43_2_c7;
   bh537_wm43_5_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid794_Out0_c7(0);
   bh537_wm42_6_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid794_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid794: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid794_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid794_Out0_copy795_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid794_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid794_Out0_copy795_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid798_In0_c7 <= "" & bh537_wm42_0_c7 & bh537_wm42_1_c7 & bh537_wm42_2_c7 & bh537_wm42_3_c7 & bh537_wm42_4_c7 & bh537_wm42_5_c7;
   bh537_wm42_7_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid798_Out0_c7(0);
   bh537_wm41_7_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid798_Out0_c7(1);
   bh537_wm40_7_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid798_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid798: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid798_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid798_Out0_copy799_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid798_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid798_Out0_copy799_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid800_In0_c7 <= "" & bh537_wm41_0_c7 & bh537_wm41_1_c7 & bh537_wm41_2_c7 & bh537_wm41_3_c7 & bh537_wm41_4_c7 & bh537_wm41_5_c7;
   bh537_wm41_8_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid800_Out0_c7(0);
   bh537_wm40_8_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid800_Out0_c7(1);
   bh537_wm39_9_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid800_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid800: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid800_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid800_Out0_copy801_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid800_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid800_Out0_copy801_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid802_In0_c7 <= "" & bh537_wm40_0_c7 & bh537_wm40_1_c7 & bh537_wm40_2_c7 & bh537_wm40_3_c7 & bh537_wm40_4_c7 & bh537_wm40_5_c7;
   bh537_wm40_9_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid802_Out0_c7(0);
   bh537_wm39_10_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid802_Out0_c7(1);
   bh537_wm38_9_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid802_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid802: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid802_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid802_Out0_copy803_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid802_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid802_Out0_copy803_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid804_In0_c7 <= "" & bh537_wm39_0_c7 & bh537_wm39_1_c7 & bh537_wm39_2_c7 & bh537_wm39_3_c7 & bh537_wm39_4_c7 & bh537_wm39_5_c7;
   bh537_wm39_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid804_Out0_c7(0);
   bh537_wm38_10_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid804_Out0_c7(1);
   bh537_wm37_10_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid804_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid804: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid804_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid804_Out0_copy805_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid804_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid804_Out0_copy805_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid806_In0_c6 <= "" & bh537_wm39_6_c6 & bh537_wm39_7_c6 & bh537_wm39_8_c6;
   Compressor_23_3_Freq300_uid781_bh537_uid806_In1_c7 <= "" & bh537_wm38_0_c7 & bh537_wm38_1_c7;
   bh537_wm39_12_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid806_Out0_c7(0);
   bh537_wm38_11_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid806_Out0_c7(1);
   bh537_wm37_11_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid806_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid806: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid806_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid806_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid806_Out0_copy807_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid806_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid806_Out0_copy807_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid808_In0_c6 <= "" & bh537_wm38_2_c6 & bh537_wm38_3_c6 & bh537_wm38_4_c6 & bh537_wm38_5_c6 & bh537_wm38_6_c6 & bh537_wm38_7_c6;
   bh537_wm38_12_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid808_Out0_c6(0);
   bh537_wm37_12_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid808_Out0_c6(1);
   bh537_wm36_11_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid808_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid808: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid808_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid808_Out0_copy809_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid808_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid808_Out0_copy809_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid810_In0_c7 <= "" & bh537_wm37_0_c7 & bh537_wm37_1_c7 & bh537_wm37_2_c7 & bh537_wm37_3_c7 & bh537_wm37_4_c7 & bh537_wm37_5_c7;
   bh537_wm37_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid810_Out0_c7(0);
   bh537_wm36_12_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid810_Out0_c7(1);
   bh537_wm35_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid810_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid810: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid810_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid810_Out0_copy811_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid810_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid810_Out0_copy811_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid814_In0_c6 <= "" & bh537_wm37_6_c6 & bh537_wm37_7_c6 & bh537_wm37_8_c6 & bh537_wm37_9_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid814_In1_c7 <= "" & bh537_wm36_0_c7;
   bh537_wm37_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid814_Out0_c7(0);
   bh537_wm36_13_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid814_Out0_c7(1);
   bh537_wm35_12_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid814_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid814: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid814_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid814_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid814_Out0_copy815_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid814_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid814_Out0_copy815_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid816_In0_c7 <= "" & bh537_wm36_1_c7 & bh537_wm36_2_c7 & bh537_wm36_3_c7 & bh537_wm36_4_c7 & bh537_wm36_5_c7 & bh537_wm36_6_c7;
   bh537_wm36_14_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid816_Out0_c7(0);
   bh537_wm35_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid816_Out0_c7(1);
   bh537_wm34_10_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid816_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid816: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid816_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid816_Out0_copy817_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid816_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid816_Out0_copy817_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid818_In0_c6 <= "" & bh537_wm36_7_c6 & bh537_wm36_8_c6 & bh537_wm36_9_c6 & bh537_wm36_10_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid818_In1_c7 <= "" & bh537_wm35_0_c7;
   bh537_wm36_15_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid818_Out0_c7(0);
   bh537_wm35_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid818_Out0_c7(1);
   bh537_wm34_11_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid818_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid818: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid818_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid818_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid818_Out0_copy819_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid818_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid818_Out0_copy819_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid820_In0_c7 <= "" & bh537_wm35_1_c7 & bh537_wm35_2_c7 & bh537_wm35_3_c7 & bh537_wm35_4_c7 & bh537_wm35_5_c7 & bh537_wm35_6_c7;
   bh537_wm35_15_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid820_Out0_c7(0);
   bh537_wm34_12_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid820_Out0_c7(1);
   bh537_wm33_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid820_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid820: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid820_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid820_Out0_copy821_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid820_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid820_Out0_copy821_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid822_In0_c6 <= "" & bh537_wm35_7_c6 & bh537_wm35_8_c6 & bh537_wm35_9_c6 & bh537_wm35_10_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid822_In1_c7 <= "" & bh537_wm34_0_c7;
   bh537_wm35_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid822_Out0_c7(0);
   bh537_wm34_13_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid822_Out0_c7(1);
   bh537_wm33_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid822_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid822: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid822_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid822_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid822_Out0_copy823_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid822_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid822_Out0_copy823_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid824_In0_c7 <= "" & bh537_wm34_1_c7 & bh537_wm34_2_c7 & bh537_wm34_3_c7 & bh537_wm34_4_c7 & bh537_wm34_5_c7 & bh537_wm34_6_c7;
   bh537_wm34_14_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid824_Out0_c7(0);
   bh537_wm33_15_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid824_Out0_c7(1);
   bh537_wm32_12_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid824_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid824: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid824_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid824_Out0_copy825_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid824_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid824_Out0_copy825_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid826_In0_c6 <= "" & bh537_wm34_7_c6 & bh537_wm34_8_c6 & bh537_wm34_9_c6;
   bh537_wm34_15_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid826_Out0_c6(0);
   bh537_wm33_16_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid826_Out0_c6(1);
   Compressor_3_2_Freq300_uid789_uid826: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid826_In0_c6,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid826_Out0_copy827_c6);
   Compressor_3_2_Freq300_uid789_bh537_uid826_Out0_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid826_Out0_copy827_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid828_In0_c7 <= "" & bh537_wm33_8_c7 & bh537_wm33_12_c7 & bh537_wm33_11_c7 & bh537_wm33_10_c7 & bh537_wm33_9_c7 & bh537_wm33_0_c7;
   bh537_wm33_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid828_Out0_c7(0);
   bh537_wm32_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid828_Out0_c7(1);
   bh537_wm31_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid828_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid828: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid828_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid828_Out0_copy829_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid828_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid828_Out0_copy829_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid830_In0_c7 <= "" & bh537_wm33_1_c7 & bh537_wm33_2_c7 & bh537_wm33_3_c7 & bh537_wm33_4_c7 & bh537_wm33_5_c7 & bh537_wm33_6_c7;
   bh537_wm33_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid830_Out0_c7(0);
   bh537_wm32_14_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid830_Out0_c7(1);
   bh537_wm31_12_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid830_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid830: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid830_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid830_Out0_copy831_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid830_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid830_Out0_copy831_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid832_In0_c7 <= "" & bh537_wm32_0_c7 & bh537_wm32_1_c7 & bh537_wm32_2_c7 & bh537_wm32_3_c7 & bh537_wm32_4_c7 & bh537_wm32_5_c7;
   bh537_wm32_15_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid832_Out0_c7(0);
   bh537_wm31_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid832_Out0_c7(1);
   bh537_wm30_12_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid832_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid832: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid832_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid832_Out0_copy833_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid832_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid832_Out0_copy833_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid834_In0_c6 <= "" & bh537_wm32_6_c6 & bh537_wm32_7_c6 & bh537_wm32_8_c6 & bh537_wm32_9_c6 & bh537_wm32_10_c6 & bh537_wm32_11_c6;
   bh537_wm32_16_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid834_Out0_c6(0);
   bh537_wm31_14_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid834_Out0_c6(1);
   bh537_wm30_13_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid834_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid834: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid834_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid834_Out0_copy835_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid834_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid834_Out0_copy835_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid836_In0_c7 <= "" & bh537_wm31_0_c7 & bh537_wm31_1_c7 & bh537_wm31_2_c7 & bh537_wm31_3_c7 & bh537_wm31_4_c7 & bh537_wm31_5_c7;
   bh537_wm31_15_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid836_Out0_c7(0);
   bh537_wm30_14_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid836_Out0_c7(1);
   bh537_wm29_12_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid836_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid836: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid836_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid836_Out0_copy837_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid836_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid836_Out0_copy837_c7; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid839_bh537_uid840_In0_c6 <= "" & bh537_wm31_6_c6 & bh537_wm31_7_c6 & bh537_wm31_8_c6 & bh537_wm31_9_c6 & bh537_wm31_10_c6;
   bh537_wm31_16_c6 <= Compressor_5_3_Freq300_uid839_bh537_uid840_Out0_c6(0);
   bh537_wm30_15_c6 <= Compressor_5_3_Freq300_uid839_bh537_uid840_Out0_c6(1);
   bh537_wm29_13_c6 <= Compressor_5_3_Freq300_uid839_bh537_uid840_Out0_c6(2);
   Compressor_5_3_Freq300_uid839_uid840: Compressor_5_3_Freq300_uid839
      port map ( X0 => Compressor_5_3_Freq300_uid839_bh537_uid840_In0_c6,
                 R => Compressor_5_3_Freq300_uid839_bh537_uid840_Out0_copy841_c6);
   Compressor_5_3_Freq300_uid839_bh537_uid840_Out0_c6 <= Compressor_5_3_Freq300_uid839_bh537_uid840_Out0_copy841_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid842_In0_c7 <= "" & bh537_wm30_0_c7 & bh537_wm30_1_c7 & bh537_wm30_2_c7 & bh537_wm30_3_c7 & bh537_wm30_4_c7 & bh537_wm30_5_c7;
   bh537_wm30_16_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid842_Out0_c7(0);
   bh537_wm29_14_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid842_Out0_c7(1);
   bh537_wm28_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid842_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid842: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid842_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid842_Out0_copy843_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid842_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid842_Out0_copy843_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid844_In0_c6 <= "" & bh537_wm30_8_c6 & bh537_wm30_11_c6 & bh537_wm30_10_c6 & bh537_wm30_9_c6 & bh537_wm30_7_c6 & bh537_wm30_6_c6;
   bh537_wm30_17_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid844_Out0_c6(0);
   bh537_wm29_15_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid844_Out0_c6(1);
   bh537_wm28_12_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid844_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid844: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid844_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid844_Out0_copy845_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid844_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid844_Out0_copy845_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid846_In0_c7 <= "" & bh537_wm29_0_c7 & bh537_wm29_1_c7 & bh537_wm29_2_c7 & bh537_wm29_3_c7 & bh537_wm29_4_c7 & bh537_wm29_5_c7;
   bh537_wm29_16_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid846_Out0_c7(0);
   bh537_wm28_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid846_Out0_c7(1);
   bh537_wm27_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid846_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid846: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid846_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid846_Out0_copy847_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid846_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid846_Out0_copy847_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid848_In0_c6 <= "" & bh537_wm29_8_c6 & bh537_wm29_11_c6 & bh537_wm29_10_c6 & bh537_wm29_9_c6 & bh537_wm29_7_c6 & bh537_wm29_6_c6;
   bh537_wm29_17_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid848_Out0_c6(0);
   bh537_wm28_14_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid848_Out0_c6(1);
   bh537_wm27_12_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid848_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid848: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid848_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid848_Out0_copy849_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid848_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid848_Out0_copy849_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid850_In0_c7 <= "" & bh537_wm28_0_c7 & bh537_wm28_1_c7 & bh537_wm28_2_c7 & bh537_wm28_3_c7 & bh537_wm28_4_c7 & bh537_wm28_5_c7;
   bh537_wm28_15_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid850_Out0_c7(0);
   bh537_wm27_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid850_Out0_c7(1);
   bh537_wm26_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid850_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid850: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid850_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid850_Out0_copy851_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid850_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid850_Out0_copy851_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid852_In0_c6 <= "" & bh537_wm28_6_c6 & bh537_wm28_7_c6 & bh537_wm28_8_c6 & bh537_wm28_9_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid852_In1_c7 <= "" & bh537_wm27_0_c7;
   bh537_wm28_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid852_Out0_c7(0);
   bh537_wm27_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid852_Out0_c7(1);
   bh537_wm26_12_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid852_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid852: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid852_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid852_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid852_Out0_copy853_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid852_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid852_Out0_copy853_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid854_In0_c6 <= "" & bh537_wm27_1_c6 & bh537_wm27_2_c6 & bh537_wm27_3_c6 & bh537_wm27_4_c6 & bh537_wm27_5_c6 & bh537_wm27_6_c6;
   bh537_wm27_15_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid854_Out0_c6(0);
   bh537_wm26_13_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid854_Out0_c6(1);
   bh537_wm25_11_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid854_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid854: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid854_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid854_Out0_copy855_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid854_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid854_Out0_copy855_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid856_In0_c6 <= "" & bh537_wm27_7_c6 & bh537_wm27_8_c6 & bh537_wm27_9_c6 & bh537_wm27_10_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid856_In1_c7 <= "" & bh537_wm26_0_c7;
   bh537_wm27_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid856_Out0_c7(0);
   bh537_wm26_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid856_Out0_c7(1);
   bh537_wm25_12_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid856_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid856: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid856_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid856_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid856_Out0_copy857_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid856_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid856_Out0_copy857_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid858_In0_c6 <= "" & bh537_wm26_1_c6 & bh537_wm26_2_c6 & bh537_wm26_3_c6 & bh537_wm26_4_c6 & bh537_wm26_5_c6 & bh537_wm26_6_c6;
   bh537_wm26_15_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid858_Out0_c6(0);
   bh537_wm25_13_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid858_Out0_c6(1);
   bh537_wm24_11_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid858_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid858: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid858_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid858_Out0_copy859_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid858_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid858_Out0_copy859_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid860_In0_c6 <= "" & bh537_wm26_7_c6 & bh537_wm26_8_c6 & bh537_wm26_9_c6 & bh537_wm26_10_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid860_In1_c7 <= "" & bh537_wm25_0_c7;
   bh537_wm26_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid860_Out0_c7(0);
   bh537_wm25_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid860_Out0_c7(1);
   bh537_wm24_12_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid860_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid860: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid860_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid860_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid860_Out0_copy861_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid860_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid860_Out0_copy861_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid862_In0_c6 <= "" & bh537_wm25_1_c6 & bh537_wm25_2_c6 & bh537_wm25_3_c6 & bh537_wm25_4_c6 & bh537_wm25_5_c6 & bh537_wm25_6_c6;
   bh537_wm25_15_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid862_Out0_c6(0);
   bh537_wm24_13_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid862_Out0_c6(1);
   bh537_wm23_11_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid862_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid862: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid862_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid862_Out0_copy863_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid862_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid862_Out0_copy863_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid864_In0_c6 <= "" & bh537_wm25_7_c6 & bh537_wm25_8_c6 & bh537_wm25_9_c6 & bh537_wm25_10_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid864_In1_c7 <= "" & bh537_wm24_0_c7;
   bh537_wm25_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid864_Out0_c7(0);
   bh537_wm24_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid864_Out0_c7(1);
   bh537_wm23_12_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid864_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid864: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid864_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid864_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid864_Out0_copy865_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid864_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid864_Out0_copy865_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid866_In0_c6 <= "" & bh537_wm24_1_c6 & bh537_wm24_2_c6 & bh537_wm24_3_c6 & bh537_wm24_4_c6 & bh537_wm24_5_c6 & bh537_wm24_6_c6;
   bh537_wm24_15_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid866_Out0_c6(0);
   bh537_wm23_13_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid866_Out0_c6(1);
   bh537_wm22_11_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid866_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid866: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid866_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid866_Out0_copy867_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid866_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid866_Out0_copy867_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid868_In0_c6 <= "" & bh537_wm24_7_c6 & bh537_wm24_8_c6 & bh537_wm24_9_c6 & bh537_wm24_10_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid868_In1_c7 <= "" & bh537_wm23_0_c7;
   bh537_wm24_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid868_Out0_c7(0);
   bh537_wm23_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid868_Out0_c7(1);
   bh537_wm22_12_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid868_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid868: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid868_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid868_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid868_Out0_copy869_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid868_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid868_Out0_copy869_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid870_In0_c6 <= "" & bh537_wm23_1_c6 & bh537_wm23_2_c6 & bh537_wm23_3_c6 & bh537_wm23_4_c6 & bh537_wm23_5_c6 & bh537_wm23_6_c6;
   bh537_wm23_15_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid870_Out0_c6(0);
   bh537_wm22_13_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid870_Out0_c6(1);
   bh537_wm21_12_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid870_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid870: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid870_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid870_Out0_copy871_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid870_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid870_Out0_copy871_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid872_In0_c6 <= "" & bh537_wm23_7_c6 & bh537_wm23_8_c6 & bh537_wm23_9_c6 & bh537_wm23_10_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid872_In1_c7 <= "" & bh537_wm22_0_c7;
   bh537_wm23_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid872_Out0_c7(0);
   bh537_wm22_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid872_Out0_c7(1);
   bh537_wm21_13_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid872_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid872: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid872_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid872_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid872_Out0_copy873_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid872_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid872_Out0_copy873_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid874_In0_c6 <= "" & bh537_wm22_1_c6 & bh537_wm22_2_c6 & bh537_wm22_3_c6 & bh537_wm22_4_c6 & bh537_wm22_5_c6 & bh537_wm22_6_c6;
   bh537_wm22_15_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid874_Out0_c6(0);
   bh537_wm21_14_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid874_Out0_c6(1);
   bh537_wm20_9_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid874_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid874: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid874_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid874_Out0_copy875_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid874_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid874_Out0_copy875_c6; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid876_In0_c6 <= "" & bh537_wm22_7_c6 & bh537_wm22_8_c6 & bh537_wm22_9_c6;
   bh537_wm22_16_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid876_Out0_c6(0);
   bh537_wm21_15_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid876_Out0_c6(1);
   Compressor_3_2_Freq300_uid789_uid876: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid876_In0_c6,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid876_Out0_copy877_c6);
   Compressor_3_2_Freq300_uid789_bh537_uid876_Out0_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid876_Out0_copy877_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid878_In0_c7 <= "" & bh537_wm21_0_c7 & bh537_wm21_1_c7 & bh537_wm21_2_c7 & bh537_wm21_3_c7 & bh537_wm21_4_c7 & bh537_wm21_5_c7;
   bh537_wm21_16_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid878_Out0_c7(0);
   bh537_wm20_10_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid878_Out0_c7(1);
   bh537_wm19_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid878_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid878: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid878_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid878_Out0_copy879_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid878_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid878_Out0_copy879_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid880_In0_c6 <= "" & bh537_wm21_8_c6 & bh537_wm21_11_c6 & bh537_wm21_10_c6 & bh537_wm21_9_c6 & bh537_wm21_7_c6 & bh537_wm21_6_c6;
   bh537_wm21_17_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid880_Out0_c6(0);
   bh537_wm20_11_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid880_Out0_c6(1);
   bh537_wm19_12_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid880_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid880: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid880_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid880_Out0_copy881_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid880_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid880_Out0_copy881_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid882_In0_c7 <= "" & bh537_wm20_0_c7 & bh537_wm20_1_c7 & bh537_wm20_2_c7 & bh537_wm20_3_c7 & bh537_wm20_4_c7 & bh537_wm20_5_c7;
   bh537_wm20_12_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid882_Out0_c7(0);
   bh537_wm19_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid882_Out0_c7(1);
   bh537_wm18_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid882_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid882: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid882_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid882_Out0_copy883_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid882_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid882_Out0_copy883_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid884_In0_c6 <= "" & bh537_wm20_6_c6 & bh537_wm20_7_c6 & bh537_wm20_8_c6;
   bh537_wm20_13_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid884_Out0_c6(0);
   bh537_wm19_14_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid884_Out0_c6(1);
   Compressor_3_2_Freq300_uid789_uid884: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid884_In0_c6,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid884_Out0_copy885_c6);
   Compressor_3_2_Freq300_uid789_bh537_uid884_Out0_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid884_Out0_copy885_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid886_In0_c7 <= "" & bh537_wm19_0_c7 & bh537_wm19_1_c7 & bh537_wm19_2_c7 & bh537_wm19_3_c7 & bh537_wm19_4_c7 & bh537_wm19_5_c7;
   bh537_wm19_15_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid886_Out0_c7(0);
   bh537_wm18_12_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid886_Out0_c7(1);
   bh537_wm17_9_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid886_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid886: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid886_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid886_Out0_copy887_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid886_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid886_Out0_copy887_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid888_In0_c6 <= "" & bh537_wm19_6_c6 & bh537_wm19_7_c6 & bh537_wm19_8_c6 & bh537_wm19_9_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid888_In1_c7 <= "" & bh537_wm18_0_c7;
   bh537_wm19_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid888_Out0_c7(0);
   bh537_wm18_13_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid888_Out0_c7(1);
   bh537_wm17_10_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid888_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid888: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid888_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid888_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid888_Out0_copy889_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid888_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid888_Out0_copy889_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid890_In0_c6 <= "" & bh537_wm18_1_c6 & bh537_wm18_2_c6 & bh537_wm18_3_c6 & bh537_wm18_4_c6 & bh537_wm18_5_c6 & bh537_wm18_6_c6;
   bh537_wm18_14_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid890_Out0_c6(0);
   bh537_wm17_11_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid890_Out0_c6(1);
   bh537_wm16_9_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid890_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid890: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid890_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid890_Out0_copy891_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid890_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid890_Out0_copy891_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid892_In0_c6 <= "" & bh537_wm18_7_c6 & bh537_wm18_8_c6 & bh537_wm18_9_c6 & bh537_wm18_10_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c0 <= "" & "0";
   bh537_wm18_15_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid892_Out0_c6(0);
   bh537_wm17_12_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid892_Out0_c6(1);
   bh537_wm16_10_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid892_Out0_c6(2);
   Compressor_14_3_Freq300_uid813_uid892: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid892_In0_c6,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid892_In1_c6,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid892_Out0_copy893_c6);
   Compressor_14_3_Freq300_uid813_bh537_uid892_Out0_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid892_Out0_copy893_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid894_In0_c7 <= "" & bh537_wm17_0_c7 & bh537_wm17_1_c7 & bh537_wm17_2_c7 & bh537_wm17_3_c7 & bh537_wm17_4_c7 & bh537_wm17_5_c7;
   bh537_wm17_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid894_Out0_c7(0);
   bh537_wm16_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid894_Out0_c7(1);
   bh537_wm15_8_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid894_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid894: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid894_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid894_Out0_copy895_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid894_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid894_Out0_copy895_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid896_In0_c6 <= "" & bh537_wm17_6_c6 & bh537_wm17_7_c6 & bh537_wm17_8_c6;
   bh537_wm17_14_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid896_Out0_c6(0);
   bh537_wm16_12_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid896_Out0_c6(1);
   Compressor_3_2_Freq300_uid789_uid896: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid896_In0_c6,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid896_Out0_copy897_c6);
   Compressor_3_2_Freq300_uid789_bh537_uid896_Out0_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid896_Out0_copy897_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid898_In0_c6 <= "" & bh537_wm16_0_c6 & bh537_wm16_1_c6 & bh537_wm16_2_c6 & bh537_wm16_3_c6 & bh537_wm16_4_c6 & bh537_wm16_5_c6;
   bh537_wm16_13_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid898_Out0_c6(0);
   bh537_wm15_9_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid898_Out0_c6(1);
   bh537_wm14_7_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid898_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid898: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid898_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid898_Out0_copy899_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid898_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid898_Out0_copy899_c6; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid900_In0_c6 <= "" & bh537_wm16_6_c6 & bh537_wm16_7_c6 & bh537_wm16_8_c6;
   Compressor_23_3_Freq300_uid781_bh537_uid900_In1_c6 <= "" & bh537_wm15_0_c6 & bh537_wm15_1_c6;
   bh537_wm16_14_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid900_Out0_c6(0);
   bh537_wm15_10_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid900_Out0_c6(1);
   bh537_wm14_8_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid900_Out0_c6(2);
   Compressor_23_3_Freq300_uid781_uid900: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid900_In0_c6,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid900_In1_c6,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid900_Out0_copy901_c6);
   Compressor_23_3_Freq300_uid781_bh537_uid900_Out0_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid900_Out0_copy901_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid902_In0_c6 <= "" & bh537_wm15_2_c6 & bh537_wm15_3_c6 & bh537_wm15_4_c6 & bh537_wm15_5_c6 & bh537_wm15_6_c6 & bh537_wm15_7_c6;
   bh537_wm15_11_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid902_Out0_c6(0);
   bh537_wm14_9_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid902_Out0_c6(1);
   bh537_wm13_6_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid902_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid902: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid902_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid902_Out0_copy903_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid902_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid902_Out0_copy903_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid904_In0_c6 <= "" & bh537_wm14_0_c6 & bh537_wm14_1_c6 & bh537_wm14_2_c6 & bh537_wm14_3_c6 & bh537_wm14_4_c6 & bh537_wm14_5_c6;
   bh537_wm14_10_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid904_Out0_c6(0);
   bh537_wm13_7_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid904_Out0_c6(1);
   bh537_wm12_6_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid904_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid904: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid904_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid904_Out0_copy905_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid904_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid904_Out0_copy905_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid906_In0_c6 <= "" & bh537_wm13_0_c6 & bh537_wm13_1_c6 & bh537_wm13_2_c6 & bh537_wm13_3_c6 & bh537_wm13_4_c6 & bh537_wm13_5_c6;
   bh537_wm13_8_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid906_Out0_c6(0);
   bh537_wm12_7_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid906_Out0_c6(1);
   bh537_wm11_4_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid906_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid906: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid906_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid906_Out0_copy907_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid906_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid906_Out0_copy907_c6; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid908_In0_c6 <= "" & bh537_wm12_0_c6 & bh537_wm12_1_c6 & bh537_wm12_2_c6 & bh537_wm12_3_c6 & bh537_wm12_4_c6 & bh537_wm12_5_c6;
   bh537_wm12_8_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid908_Out0_c6(0);
   bh537_wm11_5_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid908_Out0_c6(1);
   bh537_wm10_4_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid908_Out0_c6(2);
   Compressor_6_3_Freq300_uid797_uid908: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid908_In0_c6,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid908_Out0_copy909_c6);
   Compressor_6_3_Freq300_uid797_bh537_uid908_Out0_c6 <= Compressor_6_3_Freq300_uid797_bh537_uid908_Out0_copy909_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid910_In0_c6 <= "" & bh537_wm11_0_c6 & bh537_wm11_1_c6 & bh537_wm11_2_c6 & bh537_wm11_3_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid910_In1_c6 <= "" & bh537_wm10_0_c6;
   bh537_wm11_6_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid910_Out0_c6(0);
   bh537_wm10_5_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid910_Out0_c6(1);
   bh537_wm9_3_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid910_Out0_c6(2);
   Compressor_14_3_Freq300_uid813_uid910: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid910_In0_c6,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid910_In1_c6,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid910_Out0_copy911_c6);
   Compressor_14_3_Freq300_uid813_bh537_uid910_Out0_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid910_Out0_copy911_c6; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid912_In0_c6 <= "" & bh537_wm10_1_c6 & bh537_wm10_2_c6 & bh537_wm10_3_c6;
   Compressor_23_3_Freq300_uid781_bh537_uid912_In1_c6 <= "" & bh537_wm9_0_c6 & bh537_wm9_1_c6;
   bh537_wm10_6_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid912_Out0_c6(0);
   bh537_wm9_4_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid912_Out0_c6(1);
   bh537_wm8_2_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid912_Out0_c6(2);
   Compressor_23_3_Freq300_uid781_uid912: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid912_In0_c6,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid912_In1_c6,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid912_Out0_copy913_c6);
   Compressor_23_3_Freq300_uid781_bh537_uid912_Out0_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid912_Out0_copy913_c6; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid914_In0_c6 <= "" & bh537_wm8_0_c6 & bh537_wm8_1_c6 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid914_In1_c4 <= "" & bh537_wm7_0_c4 & bh537_wm7_1_c4;
   bh537_wm8_3_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid914_Out0_c6(0);
   bh537_wm7_2_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid914_Out0_c6(1);
   bh537_wm6_2_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid914_Out0_c6(2);
   Compressor_23_3_Freq300_uid781_uid914: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid914_In0_c6,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid914_In1_c6,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid914_Out0_copy915_c6);
   Compressor_23_3_Freq300_uid781_bh537_uid914_Out0_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid914_Out0_copy915_c6; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid916_In0_c4 <= "" & bh537_wm6_0_c4 & bh537_wm6_1_c4 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid916_In1_c4 <= "" & bh537_wm5_0_c4 & bh537_wm5_1_c4;
   bh537_wm6_3_c4 <= Compressor_23_3_Freq300_uid781_bh537_uid916_Out0_c4(0);
   bh537_wm5_2_c4 <= Compressor_23_3_Freq300_uid781_bh537_uid916_Out0_c4(1);
   bh537_wm4_2_c4 <= Compressor_23_3_Freq300_uid781_bh537_uid916_Out0_c4(2);
   Compressor_23_3_Freq300_uid781_uid916: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid916_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid916_In1_c4,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid916_Out0_copy917_c4);
   Compressor_23_3_Freq300_uid781_bh537_uid916_Out0_c4 <= Compressor_23_3_Freq300_uid781_bh537_uid916_Out0_copy917_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid918_In0_c4 <= "" & bh537_wm4_0_c4 & bh537_wm4_1_c4 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid918_In1_c4 <= "" & bh537_wm3_0_c4 & bh537_wm3_1_c4;
   bh537_wm4_3_c4 <= Compressor_23_3_Freq300_uid781_bh537_uid918_Out0_c4(0);
   bh537_wm3_2_c4 <= Compressor_23_3_Freq300_uid781_bh537_uid918_Out0_c4(1);
   bh537_wm2_1_c4 <= Compressor_23_3_Freq300_uid781_bh537_uid918_Out0_c4(2);
   Compressor_23_3_Freq300_uid781_uid918: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid918_In0_c4,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid918_In1_c4,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid918_Out0_copy919_c4);
   Compressor_23_3_Freq300_uid781_bh537_uid918_Out0_c4 <= Compressor_23_3_Freq300_uid781_bh537_uid918_Out0_copy919_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid920_In0_c7 <= "" & bh537_wm50_2_c7 & bh537_wm50_3_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid920_In1_c7 <= "" & bh537_wm49_2_c7;
   bh537_wm50_4_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid920_Out0_c7(0);
   bh537_wm49_3_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid920_Out0_c7(1);
   bh537_wm48_4_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid920_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid920: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid920_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid920_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid920_Out0_copy921_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid920_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid920_Out0_copy921_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid922_In0_c7 <= "" & bh537_wm48_2_c7 & bh537_wm48_3_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid922_In1_c7 <= "" & bh537_wm47_2_c7;
   bh537_wm48_5_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid922_Out0_c7(0);
   bh537_wm47_3_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid922_Out0_c7(1);
   bh537_wm46_4_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid922_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid922: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid922_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid922_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid922_Out0_copy923_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid922_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid922_Out0_copy923_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid924_In0_c7 <= "" & bh537_wm46_2_c7 & bh537_wm46_3_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid924_In1_c7 <= "" & bh537_wm45_3_c7 & bh537_wm45_4_c7;
   bh537_wm46_5_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid924_Out0_c7(0);
   bh537_wm45_5_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid924_Out0_c7(1);
   bh537_wm44_4_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid924_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid924: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid924_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid924_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid924_Out0_copy925_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid924_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid924_Out0_copy925_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid926_In0_c7 <= "" & bh537_wm44_2_c7 & bh537_wm44_3_c7 & "0";
   bh537_wm44_5_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid926_Out0_c7(0);
   bh537_wm43_6_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid926_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid926: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid926_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid926_Out0_copy927_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid926_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid926_Out0_copy927_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid928_In0_c7 <= "" & bh537_wm43_3_c7 & bh537_wm43_4_c7 & bh537_wm43_5_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid928_In1_c7 <= "" & bh537_wm42_6_c7 & bh537_wm42_7_c7;
   bh537_wm43_7_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid928_Out0_c7(0);
   bh537_wm42_8_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid928_Out0_c7(1);
   bh537_wm41_9_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid928_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid928: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid928_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid928_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid928_Out0_copy929_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid928_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid928_Out0_copy929_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid930_In0_c7 <= "" & bh537_wm41_6_c7 & bh537_wm41_7_c7 & bh537_wm41_8_c7;
   bh537_wm41_10_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid930_Out0_c7(0);
   bh537_wm40_10_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid930_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid930: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid930_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid930_Out0_copy931_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid930_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid930_Out0_copy931_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid932_In0_c7 <= "" & bh537_wm40_6_c7 & bh537_wm40_7_c7 & bh537_wm40_8_c7 & bh537_wm40_9_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid932_In1_c7 <= "" & bh537_wm39_9_c7;
   bh537_wm40_11_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid932_Out0_c7(0);
   bh537_wm39_13_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid932_Out0_c7(1);
   bh537_wm38_13_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid932_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid932: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid932_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid932_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid932_Out0_copy933_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid932_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid932_Out0_copy933_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid934_In0_c7 <= "" & bh537_wm39_10_c7 & bh537_wm39_11_c7 & bh537_wm39_12_c7;
   bh537_wm39_14_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid934_Out0_c7(0);
   bh537_wm38_14_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid934_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid934: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid934_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid934_Out0_copy935_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid934_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid934_Out0_copy935_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid936_In0_c7 <= "" & bh537_wm38_8_c7 & bh537_wm38_9_c7 & bh537_wm38_10_c7 & bh537_wm38_11_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid936_In1_c7 <= "" & bh537_wm37_10_c7;
   bh537_wm38_15_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid936_Out0_c7(0);
   bh537_wm37_15_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid936_Out0_c7(1);
   bh537_wm36_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid936_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid936: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid936_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid936_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid936_Out0_copy937_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid936_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid936_Out0_copy937_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid938_In0_c7 <= "" & bh537_wm37_11_c7 & bh537_wm37_12_c7 & bh537_wm37_13_c7 & bh537_wm37_14_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid938_In1_c6 <= "" & bh537_wm36_11_c6;
   bh537_wm37_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid938_Out0_c7(0);
   bh537_wm36_17_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid938_Out0_c7(1);
   bh537_wm35_17_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid938_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid938: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid938_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid938_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid938_Out0_copy939_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid938_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid938_Out0_copy939_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid940_In0_c7 <= "" & bh537_wm36_12_c7 & bh537_wm36_13_c7 & bh537_wm36_14_c7;
   bh537_wm36_18_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid940_Out0_c7(0);
   bh537_wm35_18_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid940_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid940: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid940_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid940_Out0_copy941_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid940_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid940_Out0_copy941_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid942_In0_c7 <= "" & bh537_wm35_11_c7 & bh537_wm35_12_c7 & bh537_wm35_13_c7 & bh537_wm35_14_c7 & bh537_wm35_15_c7 & bh537_wm35_16_c7;
   bh537_wm35_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid942_Out0_c7(0);
   bh537_wm34_16_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid942_Out0_c7(1);
   bh537_wm33_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid942_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid942: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid942_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid942_Out0_copy943_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid942_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid942_Out0_copy943_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid944_In0_c7 <= "" & bh537_wm34_10_c7 & bh537_wm34_11_c7 & bh537_wm34_12_c7 & bh537_wm34_13_c7 & bh537_wm34_14_c7 & bh537_wm34_15_c7;
   bh537_wm34_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid944_Out0_c7(0);
   bh537_wm33_20_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid944_Out0_c7(1);
   bh537_wm32_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid944_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid944: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid944_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid944_Out0_copy945_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid944_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid944_Out0_copy945_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid946_In0_c7 <= "" & bh537_wm33_17_c7 & bh537_wm33_7_c7 & bh537_wm33_13_c7 & bh537_wm33_14_c7 & bh537_wm33_15_c7 & bh537_wm33_16_c7;
   bh537_wm33_21_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid946_Out0_c7(0);
   bh537_wm32_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid946_Out0_c7(1);
   bh537_wm31_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid946_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid946: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid946_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid946_Out0_copy947_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid946_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid946_Out0_copy947_c7; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid839_bh537_uid948_In0_c7 <= "" & bh537_wm32_12_c7 & bh537_wm32_13_c7 & bh537_wm32_14_c7 & bh537_wm32_15_c7 & bh537_wm32_16_c7;
   bh537_wm32_19_c7 <= Compressor_5_3_Freq300_uid839_bh537_uid948_Out0_c7(0);
   bh537_wm31_18_c7 <= Compressor_5_3_Freq300_uid839_bh537_uid948_Out0_c7(1);
   bh537_wm30_18_c7 <= Compressor_5_3_Freq300_uid839_bh537_uid948_Out0_c7(2);
   Compressor_5_3_Freq300_uid839_uid948: Compressor_5_3_Freq300_uid839
      port map ( X0 => Compressor_5_3_Freq300_uid839_bh537_uid948_In0_c7,
                 R => Compressor_5_3_Freq300_uid839_bh537_uid948_Out0_copy949_c7);
   Compressor_5_3_Freq300_uid839_bh537_uid948_Out0_c7 <= Compressor_5_3_Freq300_uid839_bh537_uid948_Out0_copy949_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid950_In0_c7 <= "" & bh537_wm31_11_c7 & bh537_wm31_12_c7 & bh537_wm31_13_c7 & bh537_wm31_14_c7 & bh537_wm31_15_c7 & bh537_wm31_16_c7;
   bh537_wm31_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid950_Out0_c7(0);
   bh537_wm30_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid950_Out0_c7(1);
   bh537_wm29_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid950_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid950: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid950_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid950_Out0_copy951_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid950_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid950_Out0_copy951_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid952_In0_c7 <= "" & bh537_wm30_16_c7 & bh537_wm30_15_c7 & bh537_wm30_14_c7 & bh537_wm30_13_c7 & bh537_wm30_12_c7 & bh537_wm30_17_c7;
   bh537_wm30_20_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid952_Out0_c7(0);
   bh537_wm29_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid952_Out0_c7(1);
   bh537_wm28_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid952_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid952: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid952_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid952_Out0_copy953_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid952_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid952_Out0_copy953_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid954_In0_c7 <= "" & bh537_wm29_16_c7 & bh537_wm29_15_c7 & bh537_wm29_14_c7 & bh537_wm29_13_c7 & bh537_wm29_12_c7 & bh537_wm29_17_c7;
   bh537_wm29_20_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid954_Out0_c7(0);
   bh537_wm28_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid954_Out0_c7(1);
   bh537_wm27_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid954_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid954: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid954_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid954_Out0_copy955_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid954_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid954_Out0_copy955_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid956_In0_c7 <= "" & bh537_wm28_10_c7 & bh537_wm28_11_c7 & bh537_wm28_12_c7 & bh537_wm28_13_c7 & bh537_wm28_14_c7 & bh537_wm28_15_c7;
   bh537_wm28_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid956_Out0_c7(0);
   bh537_wm27_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid956_Out0_c7(1);
   bh537_wm26_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid956_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid956: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid956_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid956_Out0_copy957_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid956_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid956_Out0_copy957_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid958_In0_c7 <= "" & bh537_wm27_11_c7 & bh537_wm27_12_c7 & bh537_wm27_13_c7 & bh537_wm27_14_c7 & bh537_wm27_15_c7 & bh537_wm27_16_c7;
   bh537_wm27_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid958_Out0_c7(0);
   bh537_wm26_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid958_Out0_c7(1);
   bh537_wm25_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid958_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid958: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid958_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid958_Out0_copy959_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid958_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid958_Out0_copy959_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid960_In0_c7 <= "" & bh537_wm26_11_c7 & bh537_wm26_12_c7 & bh537_wm26_13_c7 & bh537_wm26_14_c7 & bh537_wm26_15_c7 & bh537_wm26_16_c7;
   bh537_wm26_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid960_Out0_c7(0);
   bh537_wm25_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid960_Out0_c7(1);
   bh537_wm24_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid960_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid960: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid960_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid960_Out0_copy961_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid960_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid960_Out0_copy961_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid962_In0_c7 <= "" & bh537_wm25_11_c7 & bh537_wm25_12_c7 & bh537_wm25_13_c7 & bh537_wm25_14_c7 & bh537_wm25_15_c7 & bh537_wm25_16_c7;
   bh537_wm25_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid962_Out0_c7(0);
   bh537_wm24_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid962_Out0_c7(1);
   bh537_wm23_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid962_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid962: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid962_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid962_Out0_copy963_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid962_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid962_Out0_copy963_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid964_In0_c7 <= "" & bh537_wm24_11_c7 & bh537_wm24_12_c7 & bh537_wm24_13_c7 & bh537_wm24_14_c7 & bh537_wm24_15_c7 & bh537_wm24_16_c7;
   bh537_wm24_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid964_Out0_c7(0);
   bh537_wm23_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid964_Out0_c7(1);
   bh537_wm22_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid964_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid964: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid964_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid964_Out0_copy965_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid964_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid964_Out0_copy965_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid966_In0_c7 <= "" & bh537_wm23_11_c7 & bh537_wm23_12_c7 & bh537_wm23_13_c7 & bh537_wm23_14_c7 & bh537_wm23_15_c7 & bh537_wm23_16_c7;
   bh537_wm23_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid966_Out0_c7(0);
   bh537_wm22_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid966_Out0_c7(1);
   bh537_wm21_18_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid966_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid966: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid966_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid966_Out0_copy967_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid966_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid966_Out0_copy967_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid968_In0_c7 <= "" & bh537_wm22_10_c7 & bh537_wm22_11_c7 & bh537_wm22_12_c7 & bh537_wm22_13_c7 & bh537_wm22_14_c7 & bh537_wm22_15_c7;
   bh537_wm22_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid968_Out0_c7(0);
   bh537_wm21_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid968_Out0_c7(1);
   bh537_wm20_14_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid968_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid968: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid968_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid968_Out0_copy969_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid968_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid968_Out0_copy969_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid970_In0_c7 <= "" & bh537_wm21_16_c7 & bh537_wm21_15_c7 & bh537_wm21_14_c7 & bh537_wm21_13_c7 & bh537_wm21_12_c7 & bh537_wm21_17_c7;
   bh537_wm21_20_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid970_Out0_c7(0);
   bh537_wm20_15_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid970_Out0_c7(1);
   bh537_wm19_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid970_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid970: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid970_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid970_Out0_copy971_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid970_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid970_Out0_copy971_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid972_In0_c7 <= "" & bh537_wm20_9_c7 & bh537_wm20_10_c7 & bh537_wm20_11_c7 & bh537_wm20_12_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c0 <= "" & bh537_wm19_10_c0;
   bh537_wm20_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid972_Out0_c7(0);
   bh537_wm19_18_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid972_Out0_c7(1);
   bh537_wm18_16_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid972_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid972: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid972_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid972_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid972_Out0_copy973_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid972_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid972_Out0_copy973_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid974_In0_c7 <= "" & bh537_wm19_11_c7 & bh537_wm19_12_c7 & bh537_wm19_13_c7 & bh537_wm19_14_c7 & bh537_wm19_15_c7 & bh537_wm19_16_c7;
   bh537_wm19_19_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid974_Out0_c7(0);
   bh537_wm18_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid974_Out0_c7(1);
   bh537_wm17_15_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid974_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid974: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid974_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid974_Out0_copy975_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid974_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid974_Out0_copy975_c7; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid839_bh537_uid976_In0_c7 <= "" & bh537_wm18_11_c7 & bh537_wm18_12_c7 & bh537_wm18_13_c7 & bh537_wm18_14_c7 & bh537_wm18_15_c7;
   bh537_wm18_18_c7 <= Compressor_5_3_Freq300_uid839_bh537_uid976_Out0_c7(0);
   bh537_wm17_16_c7 <= Compressor_5_3_Freq300_uid839_bh537_uid976_Out0_c7(1);
   bh537_wm16_15_c7 <= Compressor_5_3_Freq300_uid839_bh537_uid976_Out0_c7(2);
   Compressor_5_3_Freq300_uid839_uid976: Compressor_5_3_Freq300_uid839
      port map ( X0 => Compressor_5_3_Freq300_uid839_bh537_uid976_In0_c7,
                 R => Compressor_5_3_Freq300_uid839_bh537_uid976_Out0_copy977_c7);
   Compressor_5_3_Freq300_uid839_bh537_uid976_Out0_c7 <= Compressor_5_3_Freq300_uid839_bh537_uid976_Out0_copy977_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid978_In0_c7 <= "" & bh537_wm17_9_c7 & bh537_wm17_10_c7 & bh537_wm17_11_c7 & bh537_wm17_12_c7 & bh537_wm17_13_c7 & bh537_wm17_14_c7;
   bh537_wm17_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid978_Out0_c7(0);
   bh537_wm16_16_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid978_Out0_c7(1);
   bh537_wm15_12_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid978_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid978: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid978_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid978_Out0_copy979_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid978_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid978_Out0_copy979_c7; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid797_bh537_uid980_In0_c7 <= "" & bh537_wm16_9_c7 & bh537_wm16_10_c7 & bh537_wm16_11_c7 & bh537_wm16_12_c7 & bh537_wm16_13_c7 & bh537_wm16_14_c7;
   bh537_wm16_17_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid980_Out0_c7(0);
   bh537_wm15_13_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid980_Out0_c7(1);
   bh537_wm14_11_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid980_Out0_c7(2);
   Compressor_6_3_Freq300_uid797_uid980: Compressor_6_3_Freq300_uid797
      port map ( X0 => Compressor_6_3_Freq300_uid797_bh537_uid980_In0_c7,
                 R => Compressor_6_3_Freq300_uid797_bh537_uid980_Out0_copy981_c7);
   Compressor_6_3_Freq300_uid797_bh537_uid980_Out0_c7 <= Compressor_6_3_Freq300_uid797_bh537_uid980_Out0_copy981_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid982_In0_c7 <= "" & bh537_wm15_8_c7 & bh537_wm15_9_c7 & bh537_wm15_10_c7 & bh537_wm15_11_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c0 <= "" & bh537_wm14_6_c0;
   bh537_wm15_14_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid982_Out0_c7(0);
   bh537_wm14_12_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid982_Out0_c7(1);
   bh537_wm13_9_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid982_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid982: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid982_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid982_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid982_Out0_copy983_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid982_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid982_Out0_copy983_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid984_In0_c6 <= "" & bh537_wm14_7_c6 & bh537_wm14_8_c6 & bh537_wm14_9_c6 & bh537_wm14_10_c6;
   Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c0 <= "" & "0";
   bh537_wm14_13_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid984_Out0_c6(0);
   bh537_wm13_10_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid984_Out0_c6(1);
   bh537_wm12_9_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid984_Out0_c6(2);
   Compressor_14_3_Freq300_uid813_uid984: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid984_In0_c6,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid984_In1_c6,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid984_Out0_copy985_c6);
   Compressor_14_3_Freq300_uid813_bh537_uid984_Out0_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid984_Out0_copy985_c6; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid986_In0_c6 <= "" & bh537_wm13_6_c6 & bh537_wm13_7_c6 & bh537_wm13_8_c6;
   bh537_wm13_11_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid986_Out0_c6(0);
   bh537_wm12_10_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid986_Out0_c6(1);
   Compressor_3_2_Freq300_uid789_uid986: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid986_In0_c6,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid986_Out0_copy987_c6);
   Compressor_3_2_Freq300_uid789_bh537_uid986_Out0_c6 <= Compressor_3_2_Freq300_uid789_bh537_uid986_Out0_copy987_c6; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid988_In0_c6 <= "" & bh537_wm12_6_c6 & bh537_wm12_7_c6 & bh537_wm12_8_c6;
   Compressor_23_3_Freq300_uid781_bh537_uid988_In1_c6 <= "" & bh537_wm11_4_c6 & bh537_wm11_5_c6;
   bh537_wm12_11_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid988_Out0_c6(0);
   bh537_wm11_7_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid988_Out0_c6(1);
   bh537_wm10_7_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid988_Out0_c6(2);
   Compressor_23_3_Freq300_uid781_uid988: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid988_In0_c6,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid988_In1_c6,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid988_Out0_copy989_c6);
   Compressor_23_3_Freq300_uid781_bh537_uid988_Out0_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid988_Out0_copy989_c6; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid990_In0_c6 <= "" & bh537_wm10_4_c6 & bh537_wm10_5_c6 & bh537_wm10_6_c6;
   Compressor_23_3_Freq300_uid781_bh537_uid990_In1_c6 <= "" & bh537_wm9_2_c6 & bh537_wm9_3_c6;
   bh537_wm10_8_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid990_Out0_c6(0);
   bh537_wm9_5_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid990_Out0_c6(1);
   bh537_wm8_4_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid990_Out0_c6(2);
   Compressor_23_3_Freq300_uid781_uid990: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid990_In0_c6,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid990_In1_c6,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid990_Out0_copy991_c6);
   Compressor_23_3_Freq300_uid781_bh537_uid990_Out0_c6 <= Compressor_23_3_Freq300_uid781_bh537_uid990_Out0_copy991_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid992_In0_c6 <= "" & bh537_wm8_2_c6 & bh537_wm8_3_c6 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid992_In1_c6 <= "" & bh537_wm7_2_c6;
   bh537_wm8_5_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid992_Out0_c6(0);
   bh537_wm7_3_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid992_Out0_c6(1);
   bh537_wm6_4_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid992_Out0_c6(2);
   Compressor_14_3_Freq300_uid813_uid992: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid992_In0_c6,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid992_In1_c6,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid992_Out0_copy993_c6);
   Compressor_14_3_Freq300_uid813_bh537_uid992_Out0_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid992_Out0_copy993_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid994_In0_c6 <= "" & bh537_wm6_2_c6 & bh537_wm6_3_c6 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid994_In1_c4 <= "" & bh537_wm5_2_c4;
   bh537_wm6_5_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid994_Out0_c6(0);
   bh537_wm5_3_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid994_Out0_c6(1);
   bh537_wm4_4_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid994_Out0_c6(2);
   Compressor_14_3_Freq300_uid813_uid994: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid994_In0_c6,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid994_In1_c6,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid994_Out0_copy995_c6);
   Compressor_14_3_Freq300_uid813_bh537_uid994_Out0_c6 <= Compressor_14_3_Freq300_uid813_bh537_uid994_Out0_copy995_c6; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid996_In0_c4 <= "" & bh537_wm4_2_c4 & bh537_wm4_3_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid996_In1_c4 <= "" & bh537_wm3_2_c4;
   bh537_wm4_5_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid996_Out0_c4(0);
   bh537_wm3_3_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid996_Out0_c4(1);
   bh537_wm2_2_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid996_Out0_c4(2);
   Compressor_14_3_Freq300_uid813_uid996: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid996_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid996_In1_c4,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid996_Out0_copy997_c4);
   Compressor_14_3_Freq300_uid813_bh537_uid996_Out0_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid996_Out0_copy997_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid998_In0_c4 <= "" & bh537_wm2_0_c4 & bh537_wm2_1_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid998_In1_c0 <= "" & bh537_wm1_0_c0;
   bh537_wm2_3_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid998_Out0_c4(0);
   bh537_wm1_1_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid998_Out0_c4(1);
   Compressor_14_3_Freq300_uid813_uid998: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid998_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid998_In1_c4,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid998_Out0_copy999_c4);
   Compressor_14_3_Freq300_uid813_bh537_uid998_Out0_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid998_Out0_copy999_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1000_In0_c7 <= "" & bh537_wm48_4_c7 & bh537_wm48_5_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1000_In1_c7 <= "" & bh537_wm47_3_c7;
   bh537_wm48_6_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1000_Out0_c7(0);
   bh537_wm47_4_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1000_Out0_c7(1);
   bh537_wm46_6_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1000_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1000: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1000_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1000_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1000_Out0_copy1001_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1000_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1000_Out0_copy1001_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1002_In0_c7 <= "" & bh537_wm46_4_c7 & bh537_wm46_5_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1002_In1_c7 <= "" & bh537_wm45_5_c7;
   bh537_wm46_7_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1002_Out0_c7(0);
   bh537_wm45_6_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1002_Out0_c7(1);
   bh537_wm44_6_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1002_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1002: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1002_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1002_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1002_Out0_copy1003_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1002_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1002_Out0_copy1003_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1004_In0_c7 <= "" & bh537_wm44_4_c7 & bh537_wm44_5_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1004_In1_c7 <= "" & bh537_wm43_6_c7 & bh537_wm43_7_c7;
   bh537_wm44_7_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1004_Out0_c7(0);
   bh537_wm43_8_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1004_Out0_c7(1);
   bh537_wm42_9_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1004_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1004: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1004_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1004_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1004_Out0_copy1005_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1004_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1004_Out0_copy1005_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1006_In0_c7 <= "" & bh537_wm41_9_c7 & bh537_wm41_10_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1006_In1_c7 <= "" & bh537_wm40_10_c7 & bh537_wm40_11_c7;
   bh537_wm41_11_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1006_Out0_c7(0);
   bh537_wm40_12_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1006_Out0_c7(1);
   bh537_wm39_15_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1006_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1006: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1006_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1006_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1006_Out0_copy1007_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1006_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1006_Out0_copy1007_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid1008_In0_c7 <= "" & bh537_wm39_13_c7 & bh537_wm39_14_c7 & "0";
   bh537_wm39_16_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1008_Out0_c7(0);
   bh537_wm38_16_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1008_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid1008: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid1008_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid1008_Out0_copy1009_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid1008_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1008_Out0_copy1009_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1010_In0_c7 <= "" & bh537_wm38_12_c7 & bh537_wm38_13_c7 & bh537_wm38_14_c7 & bh537_wm38_15_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid1010_In1_c7 <= "" & bh537_wm37_15_c7;
   bh537_wm38_17_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1010_Out0_c7(0);
   bh537_wm37_17_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1010_Out0_c7(1);
   bh537_wm36_19_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1010_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1010: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1010_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1010_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1010_Out0_copy1011_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1010_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1010_Out0_copy1011_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1012_In0_c7 <= "" & bh537_wm36_15_c7 & bh537_wm36_16_c7 & bh537_wm36_17_c7 & bh537_wm36_18_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c0 <= "" & "0";
   bh537_wm36_20_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1012_Out0_c7(0);
   bh537_wm35_20_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1012_Out0_c7(1);
   bh537_wm34_18_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1012_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1012: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1012_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1012_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1012_Out0_copy1013_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1012_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1012_Out0_copy1013_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1014_In0_c7 <= "" & bh537_wm35_17_c7 & bh537_wm35_18_c7 & bh537_wm35_19_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1014_In1_c7 <= "" & bh537_wm34_16_c7 & bh537_wm34_17_c7;
   bh537_wm35_21_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1014_Out0_c7(0);
   bh537_wm34_19_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1014_Out0_c7(1);
   bh537_wm33_22_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1014_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1014: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1014_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1014_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1014_Out0_copy1015_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1014_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1014_Out0_copy1015_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1016_In0_c7 <= "" & bh537_wm33_18_c7 & bh537_wm33_19_c7 & bh537_wm33_20_c7 & bh537_wm33_21_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c0 <= "" & "0";
   bh537_wm33_23_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1016_Out0_c7(0);
   bh537_wm32_20_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1016_Out0_c7(1);
   bh537_wm31_20_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1016_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1016: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1016_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1016_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1016_Out0_copy1017_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1016_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1016_Out0_copy1017_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid1018_In0_c7 <= "" & bh537_wm32_17_c7 & bh537_wm32_18_c7 & bh537_wm32_19_c7;
   bh537_wm32_21_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1018_Out0_c7(0);
   bh537_wm31_21_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1018_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid1018: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid1018_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid1018_Out0_copy1019_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid1018_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1018_Out0_copy1019_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1020_In0_c7 <= "" & bh537_wm31_17_c7 & bh537_wm31_18_c7 & bh537_wm31_19_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1020_In1_c7 <= "" & bh537_wm30_18_c7 & bh537_wm30_19_c7;
   bh537_wm31_22_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1020_Out0_c7(0);
   bh537_wm30_21_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1020_Out0_c7(1);
   bh537_wm29_21_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1020_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1020: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1020_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1020_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1020_Out0_copy1021_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1020_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1020_Out0_copy1021_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid1022_In0_c7 <= "" & bh537_wm29_18_c7 & bh537_wm29_19_c7 & bh537_wm29_20_c7;
   bh537_wm29_22_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1022_Out0_c7(0);
   bh537_wm28_20_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1022_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid1022: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid1022_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid1022_Out0_copy1023_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid1022_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1022_Out0_copy1023_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1024_In0_c7 <= "" & bh537_wm28_16_c7 & bh537_wm28_17_c7 & bh537_wm28_18_c7 & bh537_wm28_19_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c0 <= "" & "0";
   bh537_wm28_21_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1024_Out0_c7(0);
   bh537_wm27_20_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1024_Out0_c7(1);
   bh537_wm26_20_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1024_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1024: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1024_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1024_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1024_Out0_copy1025_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1024_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1024_Out0_copy1025_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid1026_In0_c7 <= "" & bh537_wm27_17_c7 & bh537_wm27_18_c7 & bh537_wm27_19_c7;
   bh537_wm27_21_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1026_Out0_c7(0);
   bh537_wm26_21_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1026_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid1026: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid1026_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid1026_Out0_copy1027_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid1026_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1026_Out0_copy1027_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1028_In0_c7 <= "" & bh537_wm26_17_c7 & bh537_wm26_18_c7 & bh537_wm26_19_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1028_In1_c7 <= "" & bh537_wm25_17_c7 & bh537_wm25_18_c7;
   bh537_wm26_22_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1028_Out0_c7(0);
   bh537_wm25_20_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1028_Out0_c7(1);
   bh537_wm24_20_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1028_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1028: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1028_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1028_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1028_Out0_copy1029_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1028_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1028_Out0_copy1029_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1030_In0_c7 <= "" & bh537_wm24_17_c7 & bh537_wm24_18_c7 & bh537_wm24_19_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1030_In1_c7 <= "" & bh537_wm23_17_c7 & bh537_wm23_18_c7;
   bh537_wm24_21_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1030_Out0_c7(0);
   bh537_wm23_20_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1030_Out0_c7(1);
   bh537_wm22_20_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1030_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1030: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1030_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1030_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1030_Out0_copy1031_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1030_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1030_Out0_copy1031_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1032_In0_c7 <= "" & bh537_wm22_16_c7 & bh537_wm22_17_c7 & bh537_wm22_18_c7 & bh537_wm22_19_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c0 <= "" & "0";
   bh537_wm22_21_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1032_Out0_c7(0);
   bh537_wm21_21_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1032_Out0_c7(1);
   bh537_wm20_17_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1032_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1032: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1032_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1032_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1032_Out0_copy1033_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1032_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1032_Out0_copy1033_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid1034_In0_c7 <= "" & bh537_wm21_18_c7 & bh537_wm21_19_c7 & bh537_wm21_20_c7;
   bh537_wm21_22_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1034_Out0_c7(0);
   bh537_wm20_18_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1034_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid1034: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid1034_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid1034_Out0_copy1035_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid1034_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1034_Out0_copy1035_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1036_In0_c7 <= "" & bh537_wm20_13_c7 & bh537_wm20_14_c7 & bh537_wm20_15_c7 & bh537_wm20_16_c7;
   Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c0 <= "" & "0";
   bh537_wm20_19_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1036_Out0_c7(0);
   bh537_wm19_20_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1036_Out0_c7(1);
   bh537_wm18_19_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1036_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1036: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1036_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1036_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1036_Out0_copy1037_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1036_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1036_Out0_copy1037_c7; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid1038_In0_c7 <= "" & bh537_wm19_17_c7 & bh537_wm19_18_c7 & bh537_wm19_19_c7;
   bh537_wm19_21_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1038_Out0_c7(0);
   bh537_wm18_20_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1038_Out0_c7(1);
   Compressor_3_2_Freq300_uid789_uid1038: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid1038_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid1038_Out0_copy1039_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid1038_Out0_c7 <= Compressor_3_2_Freq300_uid789_bh537_uid1038_Out0_copy1039_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1040_In0_c7 <= "" & bh537_wm18_16_c7 & bh537_wm18_17_c7 & bh537_wm18_18_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1040_In1_c7 <= "" & bh537_wm17_15_c7 & bh537_wm17_16_c7;
   bh537_wm18_21_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1040_Out0_c7(0);
   bh537_wm17_18_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1040_Out0_c7(1);
   bh537_wm16_18_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1040_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1040: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1040_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1040_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1040_Out0_copy1041_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1040_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1040_Out0_copy1041_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1042_In0_c7 <= "" & bh537_wm16_15_c7 & bh537_wm16_16_c7 & bh537_wm16_17_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1042_In1_c7 <= "" & bh537_wm15_12_c7 & bh537_wm15_13_c7;
   bh537_wm16_19_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1042_Out0_c7(0);
   bh537_wm15_15_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1042_Out0_c7(1);
   bh537_wm14_14_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1042_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1042: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1042_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1042_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1042_Out0_copy1043_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1042_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1042_Out0_copy1043_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1044_In0_c7 <= "" & bh537_wm14_11_c7 & bh537_wm14_12_c7 & bh537_wm14_13_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1044_In1_c7 <= "" & bh537_wm13_9_c7 & bh537_wm13_10_c7;
   bh537_wm14_15_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1044_Out0_c7(0);
   bh537_wm13_12_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1044_Out0_c7(1);
   bh537_wm12_12_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1044_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1044: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1044_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1044_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1044_Out0_copy1045_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1044_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1044_Out0_copy1045_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1046_In0_c6 <= "" & bh537_wm12_9_c6 & bh537_wm12_10_c6 & bh537_wm12_11_c6;
   Compressor_23_3_Freq300_uid781_bh537_uid1046_In1_c6 <= "" & bh537_wm11_6_c6 & bh537_wm11_7_c6;
   bh537_wm12_13_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_c7(0);
   bh537_wm11_8_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_c7(1);
   bh537_wm10_9_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1046: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1046_In0_c6,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1046_In1_c6,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_copy1047_c6);
   Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1046_Out0_copy1047_c7; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1048_In0_c6 <= "" & bh537_wm10_7_c6 & bh537_wm10_8_c6 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1048_In1_c6 <= "" & bh537_wm9_4_c6 & bh537_wm9_5_c6;
   bh537_wm10_10_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_c7(0);
   bh537_wm9_6_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_c7(1);
   bh537_wm8_6_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_c7(2);
   Compressor_23_3_Freq300_uid781_uid1048: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1048_In0_c6,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1048_In1_c6,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_copy1049_c6);
   Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_c7 <= Compressor_23_3_Freq300_uid781_bh537_uid1048_Out0_copy1049_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1050_In0_c6 <= "" & bh537_wm8_4_c6 & bh537_wm8_5_c6 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1050_In1_c6 <= "" & bh537_wm7_3_c6;
   bh537_wm8_7_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_c7(0);
   bh537_wm7_4_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_c7(1);
   bh537_wm6_6_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1050: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1050_In0_c6,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1050_In1_c6,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_copy1051_c6);
   Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1050_Out0_copy1051_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1052_In0_c6 <= "" & bh537_wm6_4_c6 & bh537_wm6_5_c6 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1052_In1_c6 <= "" & bh537_wm5_3_c6;
   bh537_wm6_7_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_c7(0);
   bh537_wm5_4_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_c7(1);
   bh537_wm4_6_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1052: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1052_In0_c6,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1052_In1_c6,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_copy1053_c6);
   Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1052_Out0_copy1053_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1054_In0_c6 <= "" & bh537_wm4_4_c6 & bh537_wm4_5_c6 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1054_In1_c4 <= "" & bh537_wm3_3_c4;
   bh537_wm4_7_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_c7(0);
   bh537_wm3_4_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_c7(1);
   bh537_wm2_4_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1054: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1054_In0_c6,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1054_In1_c6,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_copy1055_c6);
   Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1054_Out0_copy1055_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1056_In0_c4 <= "" & bh537_wm2_2_c4 & bh537_wm2_3_c4 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1056_In1_c4 <= "" & bh537_wm1_1_c4;
   bh537_wm2_5_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid1056_Out0_c4(0);
   bh537_wm1_2_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid1056_Out0_c4(1);
   Compressor_14_3_Freq300_uid813_uid1056: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1056_In0_c4,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1056_In1_c4,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1056_Out0_copy1057_c4);
   Compressor_14_3_Freq300_uid813_bh537_uid1056_Out0_c4 <= Compressor_14_3_Freq300_uid813_bh537_uid1056_Out0_copy1057_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1058_In0_c7 <= "" & bh537_wm46_6_c7 & bh537_wm46_7_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1058_In1_c7 <= "" & bh537_wm45_6_c7;
   bh537_wm46_8_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_c8(0);
   bh537_wm45_7_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_c8(1);
   bh537_wm44_8_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_c8(2);
   Compressor_14_3_Freq300_uid813_uid1058: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1058_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1058_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_copy1059_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1058_Out0_copy1059_c8; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1060_In0_c7 <= "" & bh537_wm44_6_c7 & bh537_wm44_7_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1060_In1_c7 <= "" & bh537_wm43_8_c7;
   bh537_wm44_9_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_c8(0);
   bh537_wm43_9_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_c8(1);
   bh537_wm42_10_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_c8(2);
   Compressor_14_3_Freq300_uid813_uid1060: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1060_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1060_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_copy1061_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1060_Out0_copy1061_c8; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1062_In0_c7 <= "" & bh537_wm42_8_c7 & bh537_wm42_9_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1062_In1_c7 <= "" & bh537_wm41_11_c7;
   bh537_wm42_11_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_c8(0);
   bh537_wm41_12_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_c8(1);
   bh537_wm40_13_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_c8(2);
   Compressor_14_3_Freq300_uid813_uid1062: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1062_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1062_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_copy1063_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1062_Out0_copy1063_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1064_In0_c7 <= "" & bh537_wm39_15_c7 & bh537_wm39_16_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1064_In1_c7 <= "" & bh537_wm38_16_c7 & bh537_wm38_17_c7;
   bh537_wm39_17_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_c8(0);
   bh537_wm38_18_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_c8(1);
   bh537_wm37_18_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1064: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1064_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1064_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_copy1065_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1064_Out0_copy1065_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1066_In0_c7 <= "" & bh537_wm37_16_c7 & bh537_wm37_17_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1066_In1_c7 <= "" & bh537_wm36_19_c7 & bh537_wm36_20_c7;
   bh537_wm37_19_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_c8(0);
   bh537_wm36_21_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_c8(1);
   bh537_wm35_22_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1066: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1066_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1066_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_copy1067_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1066_Out0_copy1067_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1068_In0_c7 <= "" & bh537_wm35_20_c7 & bh537_wm35_21_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1068_In1_c7 <= "" & bh537_wm34_18_c7 & bh537_wm34_19_c7;
   bh537_wm35_23_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_c8(0);
   bh537_wm34_20_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_c8(1);
   bh537_wm33_24_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1068: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1068_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1068_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_copy1069_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1068_Out0_copy1069_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1070_In0_c7 <= "" & bh537_wm33_22_c7 & bh537_wm33_23_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1070_In1_c7 <= "" & bh537_wm32_20_c7 & bh537_wm32_21_c7;
   bh537_wm33_25_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_c8(0);
   bh537_wm32_22_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_c8(1);
   bh537_wm31_23_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1070: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1070_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1070_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_copy1071_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1070_Out0_copy1071_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1072_In0_c7 <= "" & bh537_wm31_20_c7 & bh537_wm31_21_c7 & bh537_wm31_22_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1072_In1_c7 <= "" & bh537_wm30_20_c7 & bh537_wm30_21_c7;
   bh537_wm31_24_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_c8(0);
   bh537_wm30_22_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_c8(1);
   bh537_wm29_23_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1072: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1072_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1072_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_copy1073_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1072_Out0_copy1073_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1074_In0_c7 <= "" & bh537_wm29_21_c7 & bh537_wm29_22_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1074_In1_c7 <= "" & bh537_wm28_20_c7 & bh537_wm28_21_c7;
   bh537_wm29_24_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_c8(0);
   bh537_wm28_22_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_c8(1);
   bh537_wm27_22_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1074: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1074_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1074_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_copy1075_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1074_Out0_copy1075_c8; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid789_bh537_uid1076_In0_c7 <= "" & bh537_wm27_20_c7 & bh537_wm27_21_c7 & "0";
   bh537_wm27_23_c8 <= Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_c8(0);
   bh537_wm26_23_c8 <= Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_c8(1);
   Compressor_3_2_Freq300_uid789_uid1076: Compressor_3_2_Freq300_uid789
      port map ( X0 => Compressor_3_2_Freq300_uid789_bh537_uid1076_In0_c7,
                 R => Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_copy1077_c7);
   Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_c8 <= Compressor_3_2_Freq300_uid789_bh537_uid1076_Out0_copy1077_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1078_In0_c7 <= "" & bh537_wm26_20_c7 & bh537_wm26_21_c7 & bh537_wm26_22_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1078_In1_c7 <= "" & bh537_wm25_19_c7 & bh537_wm25_20_c7;
   bh537_wm26_24_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_c8(0);
   bh537_wm25_21_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_c8(1);
   bh537_wm24_22_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1078: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1078_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1078_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_copy1079_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1078_Out0_copy1079_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1080_In0_c7 <= "" & bh537_wm24_20_c7 & bh537_wm24_21_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1080_In1_c7 <= "" & bh537_wm23_19_c7 & bh537_wm23_20_c7;
   bh537_wm24_23_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_c8(0);
   bh537_wm23_21_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_c8(1);
   bh537_wm22_22_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1080: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1080_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1080_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_copy1081_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1080_Out0_copy1081_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1082_In0_c7 <= "" & bh537_wm22_20_c7 & bh537_wm22_21_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1082_In1_c7 <= "" & bh537_wm21_21_c7 & bh537_wm21_22_c7;
   bh537_wm22_23_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_c8(0);
   bh537_wm21_23_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_c8(1);
   bh537_wm20_20_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1082: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1082_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1082_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_copy1083_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1082_Out0_copy1083_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1084_In0_c7 <= "" & bh537_wm20_17_c7 & bh537_wm20_18_c7 & bh537_wm20_19_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1084_In1_c7 <= "" & bh537_wm19_20_c7 & bh537_wm19_21_c7;
   bh537_wm20_21_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_c8(0);
   bh537_wm19_22_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_c8(1);
   bh537_wm18_22_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1084: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1084_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1084_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_copy1085_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1084_Out0_copy1085_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1086_In0_c7 <= "" & bh537_wm18_19_c7 & bh537_wm18_20_c7 & bh537_wm18_21_c7;
   Compressor_23_3_Freq300_uid781_bh537_uid1086_In1_c7 <= "" & bh537_wm17_17_c7 & bh537_wm17_18_c7;
   bh537_wm18_23_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_c8(0);
   bh537_wm17_19_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_c8(1);
   bh537_wm16_20_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1086: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1086_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1086_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_copy1087_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1086_Out0_copy1087_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1088_In0_c7 <= "" & bh537_wm16_18_c7 & bh537_wm16_19_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1088_In1_c7 <= "" & bh537_wm15_14_c7 & bh537_wm15_15_c7;
   bh537_wm16_21_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_c8(0);
   bh537_wm15_16_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_c8(1);
   bh537_wm14_16_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1088: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1088_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1088_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_copy1089_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1088_Out0_copy1089_c8; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid781_bh537_uid1090_In0_c7 <= "" & bh537_wm14_14_c7 & bh537_wm14_15_c7 & "0";
   Compressor_23_3_Freq300_uid781_bh537_uid1090_In1_c7 <= "" & bh537_wm13_11_c7 & bh537_wm13_12_c7;
   bh537_wm14_17_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_c8(0);
   bh537_wm13_13_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_c8(1);
   bh537_wm12_14_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_c8(2);
   Compressor_23_3_Freq300_uid781_uid1090: Compressor_23_3_Freq300_uid781
      port map ( X0 => Compressor_23_3_Freq300_uid781_bh537_uid1090_In0_c7,
                 X1 => Compressor_23_3_Freq300_uid781_bh537_uid1090_In1_c7,
                 R => Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_copy1091_c7);
   Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_c8 <= Compressor_23_3_Freq300_uid781_bh537_uid1090_Out0_copy1091_c8; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1092_In0_c7 <= "" & bh537_wm12_12_c7 & bh537_wm12_13_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1092_In1_c7 <= "" & bh537_wm11_8_c7;
   bh537_wm12_15_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_c8(0);
   bh537_wm11_9_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_c8(1);
   bh537_wm10_11_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_c8(2);
   Compressor_14_3_Freq300_uid813_uid1092: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1092_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1092_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_copy1093_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_c8 <= Compressor_14_3_Freq300_uid813_bh537_uid1092_Out0_copy1093_c8; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1094_In0_c7 <= "" & bh537_wm10_9_c7 & bh537_wm10_10_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1094_In1_c7 <= "" & bh537_wm9_6_c7;
   bh537_wm10_12_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1094_Out0_c7(0);
   bh537_wm9_7_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1094_Out0_c7(1);
   bh537_wm8_8_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1094_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1094: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1094_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1094_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1094_Out0_copy1095_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1094_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1094_Out0_copy1095_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1096_In0_c7 <= "" & bh537_wm8_6_c7 & bh537_wm8_7_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1096_In1_c7 <= "" & bh537_wm7_4_c7;
   bh537_wm8_9_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1096_Out0_c7(0);
   bh537_wm7_5_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1096_Out0_c7(1);
   bh537_wm6_8_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1096_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1096: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1096_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1096_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1096_Out0_copy1097_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1096_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1096_Out0_copy1097_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1098_In0_c7 <= "" & bh537_wm6_6_c7 & bh537_wm6_7_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1098_In1_c7 <= "" & bh537_wm5_4_c7;
   bh537_wm6_9_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1098_Out0_c7(0);
   bh537_wm5_5_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1098_Out0_c7(1);
   bh537_wm4_8_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1098_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1098: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1098_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1098_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1098_Out0_copy1099_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1098_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1098_Out0_copy1099_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1100_In0_c7 <= "" & bh537_wm4_6_c7 & bh537_wm4_7_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1100_In1_c7 <= "" & bh537_wm3_4_c7;
   bh537_wm4_9_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1100_Out0_c7(0);
   bh537_wm3_5_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1100_Out0_c7(1);
   bh537_wm2_6_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1100_Out0_c7(2);
   Compressor_14_3_Freq300_uid813_uid1100: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1100_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1100_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1100_Out0_copy1101_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1100_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1100_Out0_copy1101_c7; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid813_bh537_uid1102_In0_c7 <= "" & bh537_wm2_4_c7 & bh537_wm2_5_c7 & "0" & "0";
   Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c4 <= "" & bh537_wm1_2_c4;
   bh537_wm2_7_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1102_Out0_c7(0);
   bh537_wm1_3_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1102_Out0_c7(1);
   Compressor_14_3_Freq300_uid813_uid1102: Compressor_14_3_Freq300_uid813
      port map ( X0 => Compressor_14_3_Freq300_uid813_bh537_uid1102_In0_c7,
                 X1 => Compressor_14_3_Freq300_uid813_bh537_uid1102_In1_c7,
                 R => Compressor_14_3_Freq300_uid813_bh537_uid1102_Out0_copy1103_c7);
   Compressor_14_3_Freq300_uid813_bh537_uid1102_Out0_c7 <= Compressor_14_3_Freq300_uid813_bh537_uid1102_Out0_copy1103_c7; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh537_24_c8 <= bh537_wm45_7_c8 & bh537_wm46_8_c8 & bh537_wm47_4_c8 & bh537_wm48_6_c8 & bh537_wm49_3_c8 & bh537_wm50_4_c8 & bh537_wm51_2_c8 & bh537_wm52_2_c8 & bh537_wm53_0_c8 & bh537_wm54_0_c8 & bh537_wm55_0_c8 & bh537_wm56_0_c8 & bh537_wm57_0_c8 & bh537_wm58_0_c8 & bh537_wm59_0_c8 & bh537_wm60_0_c8 & bh537_wm61_0_c8 & bh537_wm62_0_c8 & bh537_wm63_0_c8 & bh537_wm64_0_c8 & bh537_wm65_0_c8 & bh537_wm66_0_c8 & bh537_wm67_0_c8 & bh537_wm68_0_c8 & bh537_wm69_0_c8;

   bitheapFinalAdd_bh537_In0_c8 <= "0" & bh537_wm1_3_c8 & bh537_wm2_6_c8 & bh537_wm3_5_c8 & bh537_wm4_8_c8 & bh537_wm5_5_c8 & bh537_wm6_8_c8 & bh537_wm7_5_c8 & bh537_wm8_8_c8 & bh537_wm9_7_c8 & bh537_wm10_11_c8 & bh537_wm11_9_c8 & bh537_wm12_14_c8 & bh537_wm13_13_c8 & bh537_wm14_16_c8 & bh537_wm15_16_c8 & bh537_wm16_20_c8 & bh537_wm17_19_c8 & bh537_wm18_22_c8 & bh537_wm19_22_c8 & bh537_wm20_20_c8 & bh537_wm21_23_c8 & bh537_wm22_22_c8 & bh537_wm23_21_c8 & bh537_wm24_22_c8 & bh537_wm25_21_c8 & bh537_wm26_23_c8 & bh537_wm27_22_c8 & bh537_wm28_22_c8 & bh537_wm29_23_c8 & bh537_wm30_22_c8 & bh537_wm31_23_c8 & bh537_wm32_22_c8 & bh537_wm33_24_c8 & bh537_wm34_20_c8 & bh537_wm35_22_c8 & bh537_wm36_21_c8 & bh537_wm37_18_c8 & bh537_wm38_18_c8 & bh537_wm39_17_c8 & bh537_wm40_12_c8 & bh537_wm41_12_c8 & bh537_wm42_10_c8 & bh537_wm43_9_c8 & bh537_wm44_8_c8;
   bitheapFinalAdd_bh537_In1_c8 <= "0" & "0" & bh537_wm2_7_c8 & "0" & bh537_wm4_9_c8 & "0" & bh537_wm6_9_c8 & "0" & bh537_wm8_9_c8 & "0" & bh537_wm10_12_c8 & "0" & bh537_wm12_15_c8 & "0" & bh537_wm14_17_c8 & "0" & bh537_wm16_21_c8 & "0" & bh537_wm18_23_c8 & "0" & bh537_wm20_21_c8 & "0" & bh537_wm22_23_c8 & "0" & bh537_wm24_23_c8 & "0" & bh537_wm26_24_c8 & bh537_wm27_23_c8 & "0" & bh537_wm29_24_c8 & "0" & bh537_wm31_24_c8 & "0" & bh537_wm33_25_c8 & "0" & bh537_wm35_23_c8 & "0" & bh537_wm37_19_c8 & "0" & "0" & bh537_wm40_13_c8 & "0" & bh537_wm42_11_c8 & "0" & bh537_wm44_9_c8;
   bitheapFinalAdd_bh537_Cin_c0 <= '0';

   bitheapFinalAdd_bh537: IntAdder_45_Freq300_uid1105
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 Cin => bitheapFinalAdd_bh537_Cin_c0,
                 X => bitheapFinalAdd_bh537_In0_c8,
                 Y => bitheapFinalAdd_bh537_In1_c8,
                 R => bitheapFinalAdd_bh537_Out_c8);
   bitheapResult_bh537_c8 <= bitheapFinalAdd_bh537_Out_c8(43 downto 0) & tmp_bitheapResult_bh537_24_c8;
   RR_c8 <= signed(bitheapResult_bh537_c8(68 downto 28));
R <= std_logic_vector(RR_c8);  
end architecture;

--------------------------------------------------------------------------------
--                      FixHornerEvaluator_Freq300_uid64
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin (2014-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: Y A0 A1 A2
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixHornerEvaluator_Freq300_uid64 is
    port (clk, ce_5, ce_6, ce_7, ce_8 : in std_logic;
          Y : in  std_logic_vector(28 downto 0);
          A0 : in  std_logic_vector(39 downto 0);
          A1 : in  std_logic_vector(32 downto 0);
          A2 : in  std_logic_vector(24 downto 0);
          R : out  std_logic_vector(35 downto 0)   );
end entity;

architecture arch of FixHornerEvaluator_Freq300_uid64 is
   component FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid66 is
      port ( clk, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(24 downto 0);
             Y : in  std_logic_vector(24 downto 0);
             A : in  std_logic_vector(32 downto 0);
             R : out  std_logic_vector(32 downto 0)   );
   end component;

   component FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid536 is
      port ( clk, ce_5, ce_6, ce_7, ce_8 : in std_logic;
             X : in  std_logic_vector(28 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             A : in  std_logic_vector(39 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

signal Ys_c4 :  signed(0+28 downto 0);
signal As0_c4 :  signed(-2+41 downto 0);
signal As1_c4 :  signed(-9+41 downto 0);
signal As2_c4 :  signed(-17+41 downto 0);
signal S2_c4 :  signed(-17+41 downto 0);
signal YsTrunc1_c4 :  signed(0+24 downto 0);
signal SS1_c6 :  std_logic_vector(32 downto 0);
signal S1_c6 :  signed(-9+41 downto 0);
signal YsTrunc0_c4 :  signed(0+28 downto 0);
signal SS0_c8 :  std_logic_vector(40 downto 0);
signal S0_c8 :  signed(-1+41 downto 0);
signal Rs_c8 :  signed(-2+37 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
            end if;
            if ce_6 = '1' then
            end if;
            if ce_7 = '1' then
            end if;
            if ce_8 = '1' then
            end if;
         end if;
      end process;
   Ys_c4 <= signed(Y);
   As0_c4 <= signed(A0);
   As1_c4 <= signed(A1);
   As2_c4 <= signed(A2);
   S2_c4 <= As2_c4(24 downto 0); -- fix resize from (-17, -41) to (-17, -41)
   YsTrunc1_c4 <= Ys_c4(28 downto 4); -- fix resize from (0, -28) to (0, -24)
   FixHornerEvaluator_Freq300_uid64_step_1: FixMultAdd_signed_x_0_M24_y_M17_M41_a_M9_M41_r_M9_M41_Freq300_uid66
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 A => std_logic_vector(As1_c4),
                 X => std_logic_vector(YsTrunc1_c4),
                 Y => std_logic_vector(S2_c4),
                 R => SS1_c6);
S1_c6 <= signed(SS1_c6);
   YsTrunc0_c4 <= Ys_c4(28 downto 0); -- fix resize from (0, -28) to (0, -28)
   FixHornerEvaluator_Freq300_uid64_step_0: FixMultAdd_signed_x_0_M28_y_M9_M41_a_M2_M41_r_M1_M41_Freq300_uid536
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 A => std_logic_vector(As0_c4),
                 X => std_logic_vector(YsTrunc0_c4),
                 Y => std_logic_vector(S1_c6),
                 R => SS0_c8);
S0_c8 <= signed(SS0_c8);
   Rs_c8 <= S0_c8(39 downto 4); -- fix resize from (-1, -41) to (-2, -37)
   R <= std_logic_vector(Rs_c8);
end architecture;

--------------------------------------------------------------------------------
--                  FixFunctionByPiecewisePoly_Freq300_uid59
-- Evaluator for 1b19*(exp(x*1b-10)-x*1b-10-1) on [0,1) for lsbIn=-36 (wIn=36), msbout=-2, lsbOut=-37 (wOut=36). Out interval: [0; 0.250081]. Output is unsigned

-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2014-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByPiecewisePoly_Freq300_uid59 is
    port (clk, ce_5, ce_6, ce_7, ce_8 : in std_logic;
          X : in  std_logic_vector(35 downto 0);
          Y : out  std_logic_vector(35 downto 0)   );
end entity;

architecture arch of FixFunctionByPiecewisePoly_Freq300_uid59 is
   component coeffTable_Freq300_uid61 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(94 downto 0)   );
   end component;

   component FixHornerEvaluator_Freq300_uid64 is
      port ( clk, ce_5, ce_6, ce_7, ce_8 : in std_logic;
             Y : in  std_logic_vector(28 downto 0);
             A0 : in  std_logic_vector(39 downto 0);
             A1 : in  std_logic_vector(32 downto 0);
             A2 : in  std_logic_vector(24 downto 0);
             R : out  std_logic_vector(35 downto 0)   );
   end component;

signal A_c4 :  std_logic_vector(6 downto 0);
signal Z_c4 :  std_logic_vector(28 downto 0);
signal Zs_c4 :  std_logic_vector(28 downto 0);
signal Coeffs_c4 :  std_logic_vector(94 downto 0);
signal Coeffs_copy62_c4 :  std_logic_vector(94 downto 0);
signal A2_c4 :  std_logic_vector(24 downto 0);
signal A1_c4 :  std_logic_vector(32 downto 0);
signal A0_c4 :  std_logic_vector(39 downto 0);
signal HornerOutput_c8 :  std_logic_vector(35 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
            end if;
            if ce_6 = '1' then
            end if;
            if ce_7 = '1' then
            end if;
            if ce_8 = '1' then
            end if;
         end if;
      end process;
   A_c4 <= X(35 downto 29);
   Z_c4 <= X(28 downto 0);
   Zs_c4 <= (not Z_c4(28)) & Z_c4(27 downto 0); -- centering the interval
   coeffTable: coeffTable_Freq300_uid61
      port map ( X => A_c4,
                 Y => Coeffs_copy62_c4);
   Coeffs_c4 <= Coeffs_copy62_c4; -- output copy to hold a pipeline register if needed
   --  Split the table output into each coefficient, adding back the constant signs if any
   A2_c4 <= "0" & Coeffs_c4(23 downto 0);
   A1_c4 <= "0" & Coeffs_c4(55 downto 24);
   A0_c4 <= "0" & Coeffs_c4(94 downto 56);
   Horner: FixHornerEvaluator_Freq300_uid64
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 A0 => A0_c4,
                 A1 => A1_c4,
                 A2 => A2_c4,
                 Y => Zs_c4,
                 R => HornerOutput_c8);
   Y <= std_logic_vector(HornerOutput_c8);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_47_Freq300_uid1108
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_47_Freq300_uid1108 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(46 downto 0);
          Y : in  std_logic_vector(46 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(46 downto 0)   );
end entity;

architecture arch of IntAdder_47_Freq300_uid1108 is
signal Rtmp_c9 :  std_logic_vector(46 downto 0);
signal X_c5, X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(46 downto 0);
signal Y_c9 :  std_logic_vector(46 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               X_c5 <= X;
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               X_c6 <= X_c5;
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
               Y_c9 <= Y;
               Cin_c9 <= Cin_c8;
            end if;
         end if;
      end process;
   Rtmp_c9 <= X_c9 + Y_c9 + Cin_c9;
   R <= Rtmp_c9;
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x24_Freq300_uid1114
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid1114 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid1114 is
signal Mfull_c9 :  std_logic_vector(40 downto 0);
signal M_c9 :  std_logic_vector(40 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(16 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
   Mfull_c9 <= std_logic_vector(unsigned(X_c9) * unsigned(Y)); -- multiplier
   M_c9 <= Mfull_c9(40 downto 0);
   R <= M_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1116
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1116 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1116 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1118
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1118 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1118 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid1120
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid1120 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid1120 is
   component MultTable_Freq300_uid1122 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(3 downto 0);
signal Y1_c9 :  std_logic_vector(3 downto 0);
signal Y1_copy1123_c9 :  std_logic_vector(3 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1122
      port map ( X => Xtable_c9,
                 Y => Y1_copy1123_c9);
   Y1_c9 <= Y1_copy1123_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1125
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1125 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1125 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid1127
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid1127 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid1127 is
signal replicated_c9 :  std_logic_vector(1 downto 0);
signal prod_c9 :  std_logic_vector(1 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
   replicated_c9 <= (1 downto 0 => Y(0));
   prod_c9 <= X_c9 and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1129
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1129 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1129 is
   component MultTable_Freq300_uid1131 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1132_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1131
      port map ( X => Xtable_c9,
                 Y => Y1_copy1132_c9);
   Y1_c9 <= Y1_copy1132_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1134
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1134 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1134 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1136
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1136 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1136 is
   component MultTable_Freq300_uid1138 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1139_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1138
      port map ( X => Xtable_c9,
                 Y => Y1_copy1139_c9);
   Y1_c9 <= Y1_copy1139_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1141
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1141 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1141 is
   component MultTable_Freq300_uid1143 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1144_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1143
      port map ( X => Xtable_c9,
                 Y => Y1_copy1144_c9);
   Y1_c9 <= Y1_copy1144_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1146
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1146 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1146 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid1148
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid1148 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid1148 is
   component MultTable_Freq300_uid1150 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(3 downto 0);
signal Y1_c9 :  std_logic_vector(3 downto 0);
signal Y1_copy1151_c9 :  std_logic_vector(3 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1150
      port map ( X => Xtable_c9,
                 Y => Y1_copy1151_c9);
   Y1_c9 <= Y1_copy1151_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1153
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1153 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1153 is
   component MultTable_Freq300_uid1155 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1156_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1155
      port map ( X => Xtable_c9,
                 Y => Y1_copy1156_c9);
   Y1_c9 <= Y1_copy1156_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1158
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1158 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1158 is
   component MultTable_Freq300_uid1160 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1161_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1160
      port map ( X => Xtable_c9,
                 Y => Y1_copy1161_c9);
   Y1_c9 <= Y1_copy1161_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1163
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1163 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1163 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid1165
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid1165 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid1165 is
signal replicated_c9 :  std_logic_vector(1 downto 0);
signal prod_c9 :  std_logic_vector(1 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
   replicated_c9 <= (1 downto 0 => Y(0));
   prod_c9 <= X_c9 and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1167
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1167 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1167 is
   component MultTable_Freq300_uid1169 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1170_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1169
      port map ( X => Xtable_c9,
                 Y => Y1_copy1170_c9);
   Y1_c9 <= Y1_copy1170_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1172
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1172 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1172 is
   component MultTable_Freq300_uid1174 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1175_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1174
      port map ( X => Xtable_c9,
                 Y => Y1_copy1175_c9);
   Y1_c9 <= Y1_copy1175_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1177
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1177 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1177 is
   component MultTable_Freq300_uid1179 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1180_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1179
      port map ( X => Xtable_c9,
                 Y => Y1_copy1180_c9);
   Y1_c9 <= Y1_copy1180_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1182
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1182 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1182 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1184
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1184 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1184 is
   component MultTable_Freq300_uid1186 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1187_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1186
      port map ( X => Xtable_c9,
                 Y => Y1_copy1187_c9);
   Y1_c9 <= Y1_copy1187_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1189
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1189 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1189 is
   component MultTable_Freq300_uid1191 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1192_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1191
      port map ( X => Xtable_c9,
                 Y => Y1_copy1192_c9);
   Y1_c9 <= Y1_copy1192_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1194
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1194 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1194 is
   component MultTable_Freq300_uid1196 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1197_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1196
      port map ( X => Xtable_c9,
                 Y => Y1_copy1197_c9);
   Y1_c9 <= Y1_copy1197_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1199
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1199 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1199 is
   component MultTable_Freq300_uid1201 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1202_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1201
      port map ( X => Xtable_c9,
                 Y => Y1_copy1202_c9);
   Y1_c9 <= Y1_copy1202_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x23_Freq300_uid1204
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x23_Freq300_uid1204 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(22 downto 0);
          R : out  std_logic_vector(39 downto 0)   );
end entity;

architecture arch of DSPBlock_17x23_Freq300_uid1204 is
signal Mfull_c9 :  std_logic_vector(39 downto 0);
signal M_c9 :  std_logic_vector(39 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(16 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
   Mfull_c9 <= std_logic_vector(unsigned(X_c9) * unsigned(Y)); -- multiplier
   M_c9 <= Mfull_c9(39 downto 0);
   R <= M_c9;
end architecture;

--------------------------------------------------------------------------------
--                       DSPBlock_17x23_Freq300_uid1206
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x23_Freq300_uid1206 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(22 downto 0);
          R : out  std_logic_vector(39 downto 0)   );
end entity;

architecture arch of DSPBlock_17x23_Freq300_uid1206 is
signal Mfull_c9 :  std_logic_vector(39 downto 0);
signal M_c9 :  std_logic_vector(39 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(16 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
   Mfull_c9 <= std_logic_vector(unsigned(X_c9) * unsigned(Y)); -- multiplier
   M_c9 <= Mfull_c9(39 downto 0);
   R <= M_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1208
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1208 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1208 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1210
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1210 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1210 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid1212
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid1212 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid1212 is
   component MultTable_Freq300_uid1214 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(3 downto 0);
signal Y1_c9 :  std_logic_vector(3 downto 0);
signal Y1_copy1215_c9 :  std_logic_vector(3 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1214
      port map ( X => Xtable_c9,
                 Y => Y1_copy1215_c9);
   Y1_c9 <= Y1_copy1215_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1217
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1217 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1217 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid1219
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid1219 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid1219 is
signal replicated_c9 :  std_logic_vector(1 downto 0);
signal prod_c9 :  std_logic_vector(1 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
   replicated_c9 <= (1 downto 0 => Y(0));
   prod_c9 <= X_c9 and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1221
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1221 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1221 is
   component MultTable_Freq300_uid1223 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1224_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1223
      port map ( X => Xtable_c9,
                 Y => Y1_copy1224_c9);
   Y1_c9 <= Y1_copy1224_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1226
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1226 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1226 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1228
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1228 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1228 is
   component MultTable_Freq300_uid1230 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1231_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1230
      port map ( X => Xtable_c9,
                 Y => Y1_copy1231_c9);
   Y1_c9 <= Y1_copy1231_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1233
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1233 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1233 is
   component MultTable_Freq300_uid1235 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1236_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1235
      port map ( X => Xtable_c9,
                 Y => Y1_copy1236_c9);
   Y1_c9 <= Y1_copy1236_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1238
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1238 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1238 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid1240
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid1240 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid1240 is
   component MultTable_Freq300_uid1242 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(3 downto 0);
signal Y1_c9 :  std_logic_vector(3 downto 0);
signal Y1_copy1243_c9 :  std_logic_vector(3 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1242
      port map ( X => Xtable_c9,
                 Y => Y1_copy1243_c9);
   Y1_c9 <= Y1_copy1243_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1245
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1245 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1245 is
   component MultTable_Freq300_uid1247 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1248_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1247
      port map ( X => Xtable_c9,
                 Y => Y1_copy1248_c9);
   Y1_c9 <= Y1_copy1248_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1250
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1250 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1250 is
   component MultTable_Freq300_uid1252 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1253_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1252
      port map ( X => Xtable_c9,
                 Y => Y1_copy1253_c9);
   Y1_c9 <= Y1_copy1253_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid1255
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid1255 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid1255 is
signal replicated_c5, replicated_c6, replicated_c7, replicated_c8, replicated_c9 :  std_logic_vector(0 downto 0);
signal prod_c9 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               replicated_c6 <= replicated_c5;
            end if;
            if ce_7 = '1' then
               replicated_c7 <= replicated_c6;
            end if;
            if ce_8 = '1' then
               replicated_c8 <= replicated_c7;
            end if;
            if ce_9 = '1' then
               replicated_c9 <= replicated_c8;
            end if;
         end if;
      end process;
   replicated_c5 <= (0 downto 0 => X(0));
   prod_c9 <= Y and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq300_uid1257
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq300_uid1257 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq300_uid1257 is
signal replicated_c9 :  std_logic_vector(1 downto 0);
signal prod_c9 :  std_logic_vector(1 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
   replicated_c9 <= (1 downto 0 => Y(0));
   prod_c9 <= X_c9 and replicated_c9;
   R <= prod_c9;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1259
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1259 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1259 is
   component MultTable_Freq300_uid1261 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1262_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1261
      port map ( X => Xtable_c9,
                 Y => Y1_copy1262_c9);
   Y1_c9 <= Y1_copy1262_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1264
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1264 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1264 is
   component MultTable_Freq300_uid1266 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1267_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1266
      port map ( X => Xtable_c9,
                 Y => Y1_copy1267_c9);
   Y1_c9 <= Y1_copy1267_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1269
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1269 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1269 is
   component MultTable_Freq300_uid1271 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1272_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1271
      port map ( X => Xtable_c9,
                 Y => Y1_copy1272_c9);
   Y1_c9 <= Y1_copy1272_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1274
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1274 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1274 is
   component MultTable_Freq300_uid1276 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1277_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1276
      port map ( X => Xtable_c9,
                 Y => Y1_copy1277_c9);
   Y1_c9 <= Y1_copy1277_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1279
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1279 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1279 is
   component MultTable_Freq300_uid1281 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1282_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1281
      port map ( X => Xtable_c9,
                 Y => Y1_copy1282_c9);
   Y1_c9 <= Y1_copy1282_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1284
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1284 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1284 is
   component MultTable_Freq300_uid1286 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1287_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1286
      port map ( X => Xtable_c9,
                 Y => Y1_copy1287_c9);
   Y1_c9 <= Y1_copy1287_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1289
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1289 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1289 is
   component MultTable_Freq300_uid1291 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1292_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1291
      port map ( X => Xtable_c9,
                 Y => Y1_copy1292_c9);
   Y1_c9 <= Y1_copy1292_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1294
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1294 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1294 is
   component MultTable_Freq300_uid1296 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1297_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1296
      port map ( X => Xtable_c9,
                 Y => Y1_copy1297_c9);
   Y1_c9 <= Y1_copy1297_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1299
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1299 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1299 is
   component MultTable_Freq300_uid1301 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1302_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1301
      port map ( X => Xtable_c9,
                 Y => Y1_copy1302_c9);
   Y1_c9 <= Y1_copy1302_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1304
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1304 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1304 is
   component MultTable_Freq300_uid1306 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1307_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1306
      port map ( X => Xtable_c9,
                 Y => Y1_copy1307_c9);
   Y1_c9 <= Y1_copy1307_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1309
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1309 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1309 is
   component MultTable_Freq300_uid1311 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1312_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1311
      port map ( X => Xtable_c9,
                 Y => Y1_copy1312_c9);
   Y1_c9 <= Y1_copy1312_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1314
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1314 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1314 is
   component MultTable_Freq300_uid1316 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1317_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1316
      port map ( X => Xtable_c9,
                 Y => Y1_copy1317_c9);
   Y1_c9 <= Y1_copy1317_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1319
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1319 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1319 is
   component MultTable_Freq300_uid1321 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1322_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1321
      port map ( X => Xtable_c9,
                 Y => Y1_copy1322_c9);
   Y1_c9 <= Y1_copy1322_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1324
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1324 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1324 is
   component MultTable_Freq300_uid1326 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1327_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1326
      port map ( X => Xtable_c9,
                 Y => Y1_copy1327_c9);
   Y1_c9 <= Y1_copy1327_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1329
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1329 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1329 is
   component MultTable_Freq300_uid1331 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1332_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1331
      port map ( X => Xtable_c9,
                 Y => Y1_copy1332_c9);
   Y1_c9 <= Y1_copy1332_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1334
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1334 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1334 is
   component MultTable_Freq300_uid1336 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1337_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1336
      port map ( X => Xtable_c9,
                 Y => Y1_copy1337_c9);
   Y1_c9 <= Y1_copy1337_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1339
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1339 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1339 is
   component MultTable_Freq300_uid1341 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1342_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1341
      port map ( X => Xtable_c9,
                 Y => Y1_copy1342_c9);
   Y1_c9 <= Y1_copy1342_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1344
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1344 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1344 is
   component MultTable_Freq300_uid1346 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1347_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1346
      port map ( X => Xtable_c9,
                 Y => Y1_copy1347_c9);
   Y1_c9 <= Y1_copy1347_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid1349
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid1349 is
    port (clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid1349 is
   component MultTable_Freq300_uid1351 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c9 :  std_logic_vector(4 downto 0);
signal Y1_c9 :  std_logic_vector(4 downto 0);
signal Y1_copy1352_c9 :  std_logic_vector(4 downto 0);
signal X_c6, X_c7, X_c8, X_c9 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               X_c6 <= X;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
            end if;
         end if;
      end process;
Xtable_c9 <= Y & X_c9;
   R <= Y1_c9;
   TableMult: MultTable_Freq300_uid1351
      port map ( X => Xtable_c9,
                 Y => Y1_copy1352_c9);
   Y1_c9 <= Y1_copy1352_c9; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_50_Freq300_uid1699
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_50_Freq300_uid1699 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(49 downto 0);
          Y : in  std_logic_vector(49 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(49 downto 0)   );
end entity;

architecture arch of IntAdder_50_Freq300_uid1699 is
signal Rtmp_c11 :  std_logic_vector(49 downto 0);
signal X_c11 :  std_logic_vector(49 downto 0);
signal Y_c11 :  std_logic_vector(49 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               X_c11 <= X;
               Y_c11 <= Y;
               Cin_c11 <= Cin_c10;
            end if;
         end if;
      end process;
   Rtmp_c11 <= X_c11 + Y_c11 + Cin_c11;
   R <= Rtmp_c11;
end architecture;

--------------------------------------------------------------------------------
--                   IntMultiplier_46x47_48_Freq300_uid1110
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_46x47_48_Freq300_uid1110 is
    port (clk, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(45 downto 0);
          Y : in  std_logic_vector(46 downto 0);
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_46x47_48_Freq300_uid1110 is
   component DSPBlock_17x24_Freq300_uid1114 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1116 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1118 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid1120 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1125 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid1127 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1129 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1134 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1136 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1141 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1146 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid1148 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1153 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1158 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1163 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid1165 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1167 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1172 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1177 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1182 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1184 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1189 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1194 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1199 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_17x23_Freq300_uid1204 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(22 downto 0);
             R : out  std_logic_vector(39 downto 0)   );
   end component;

   component DSPBlock_17x23_Freq300_uid1206 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(22 downto 0);
             R : out  std_logic_vector(39 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1208 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1210 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid1212 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1217 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid1219 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1221 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1226 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1228 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1233 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1238 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid1240 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1245 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1250 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid1255 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq300_uid1257 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1259 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1264 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1269 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1274 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1279 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1284 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1289 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1294 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1299 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1304 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1309 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1314 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1319 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1324 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1329 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1334 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1339 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1344 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid1349 is
      port ( clk, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid1355 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid1359 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid1363 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid1373 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq300_uid1557 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_50_Freq300_uid1699 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(49 downto 0);
             Y : in  std_logic_vector(49 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(49 downto 0)   );
   end component;

signal XX_m1111_c5 :  std_logic_vector(45 downto 0);
signal YY_m1111_c9 :  std_logic_vector(46 downto 0);
signal tile_0_X_c5 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c9 :  std_logic_vector(23 downto 0);
signal tile_0_output_c9 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c9 :  unsigned(40-0 downto 0);
signal bh1112_w29_0_c9, bh1112_w29_0_c10 :  std_logic;
signal bh1112_w30_0_c9, bh1112_w30_0_c10 :  std_logic;
signal bh1112_w31_0_c9, bh1112_w31_0_c10 :  std_logic;
signal bh1112_w32_0_c9, bh1112_w32_0_c10 :  std_logic;
signal bh1112_w33_0_c9, bh1112_w33_0_c10 :  std_logic;
signal bh1112_w34_0_c9, bh1112_w34_0_c10 :  std_logic;
signal bh1112_w35_0_c9, bh1112_w35_0_c10 :  std_logic;
signal bh1112_w36_0_c9 :  std_logic;
signal bh1112_w37_0_c9 :  std_logic;
signal bh1112_w38_0_c9 :  std_logic;
signal bh1112_w39_0_c9 :  std_logic;
signal bh1112_w40_0_c9 :  std_logic;
signal bh1112_w41_0_c9 :  std_logic;
signal bh1112_w42_0_c9 :  std_logic;
signal bh1112_w43_0_c9 :  std_logic;
signal bh1112_w44_0_c9 :  std_logic;
signal bh1112_w45_0_c9 :  std_logic;
signal bh1112_w46_0_c9 :  std_logic;
signal bh1112_w47_0_c9 :  std_logic;
signal bh1112_w48_0_c9 :  std_logic;
signal bh1112_w49_0_c9 :  std_logic;
signal bh1112_w50_0_c9 :  std_logic;
signal bh1112_w51_0_c9 :  std_logic;
signal bh1112_w52_0_c9 :  std_logic;
signal bh1112_w53_0_c9 :  std_logic;
signal bh1112_w54_0_c9 :  std_logic;
signal bh1112_w55_0_c9 :  std_logic;
signal bh1112_w56_0_c9 :  std_logic;
signal bh1112_w57_0_c9 :  std_logic;
signal bh1112_w58_0_c9 :  std_logic;
signal bh1112_w59_0_c9 :  std_logic;
signal bh1112_w60_0_c9 :  std_logic;
signal bh1112_w61_0_c9 :  std_logic;
signal bh1112_w62_0_c9 :  std_logic;
signal bh1112_w63_0_c9 :  std_logic;
signal bh1112_w64_0_c9 :  std_logic;
signal bh1112_w65_0_c9 :  std_logic;
signal bh1112_w66_0_c9 :  std_logic;
signal bh1112_w67_0_c9 :  std_logic;
signal bh1112_w68_0_c9 :  std_logic;
signal bh1112_w69_0_c9 :  std_logic;
signal tile_1_X_c5 :  std_logic_vector(0 downto 0);
signal tile_1_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_1_output_c9 :  std_logic_vector(0 downto 0);
signal tile_1_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_1_c9 :  std_logic;
signal tile_2_X_c5 :  std_logic_vector(0 downto 0);
signal tile_2_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_2_output_c9 :  std_logic_vector(0 downto 0);
signal tile_2_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_2_c9 :  std_logic;
signal tile_3_X_c5 :  std_logic_vector(1 downto 0);
signal tile_3_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_3_output_c9 :  std_logic_vector(3 downto 0);
signal tile_3_filtered_output_c9 :  unsigned(3-0 downto 0);
signal bh1112_w39_3_c9 :  std_logic;
signal bh1112_w40_1_c9 :  std_logic;
signal bh1112_w41_1_c9 :  std_logic;
signal bh1112_w42_1_c9 :  std_logic;
signal tile_4_X_c5 :  std_logic_vector(0 downto 0);
signal tile_4_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_4_output_c9 :  std_logic_vector(0 downto 0);
signal tile_4_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_4_c9 :  std_logic;
signal tile_5_X_c5 :  std_logic_vector(1 downto 0);
signal tile_5_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_5_output_c9 :  std_logic_vector(1 downto 0);
signal tile_5_filtered_output_c9 :  unsigned(1-0 downto 0);
signal bh1112_w39_5_c9 :  std_logic;
signal bh1112_w40_2_c9 :  std_logic;
signal tile_6_X_c5 :  std_logic_vector(2 downto 0);
signal tile_6_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_6_output_c9 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w40_3_c9 :  std_logic;
signal bh1112_w41_2_c9 :  std_logic;
signal bh1112_w42_2_c9 :  std_logic;
signal bh1112_w43_1_c9 :  std_logic;
signal bh1112_w44_1_c9 :  std_logic;
signal tile_7_X_c5 :  std_logic_vector(0 downto 0);
signal tile_7_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_7_output_c9 :  std_logic_vector(0 downto 0);
signal tile_7_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_6_c9 :  std_logic;
signal tile_8_X_c5 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_8_output_c9 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w39_7_c9 :  std_logic;
signal bh1112_w40_4_c9 :  std_logic;
signal bh1112_w41_3_c9 :  std_logic;
signal bh1112_w42_3_c9 :  std_logic;
signal bh1112_w43_2_c9 :  std_logic;
signal tile_9_X_c5 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_9_output_c9 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w42_4_c9 :  std_logic;
signal bh1112_w43_3_c9 :  std_logic;
signal bh1112_w44_2_c9 :  std_logic;
signal bh1112_w45_1_c9 :  std_logic;
signal bh1112_w46_1_c9 :  std_logic;
signal tile_10_X_c5 :  std_logic_vector(0 downto 0);
signal tile_10_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_10_output_c9 :  std_logic_vector(0 downto 0);
signal tile_10_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_8_c9 :  std_logic;
signal tile_11_X_c5 :  std_logic_vector(1 downto 0);
signal tile_11_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_11_output_c9 :  std_logic_vector(3 downto 0);
signal tile_11_filtered_output_c9 :  unsigned(3-0 downto 0);
signal bh1112_w39_9_c9 :  std_logic;
signal bh1112_w40_5_c9 :  std_logic;
signal bh1112_w41_4_c9 :  std_logic;
signal bh1112_w42_5_c9 :  std_logic;
signal tile_12_X_c5 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_12_output_c9 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w41_5_c9 :  std_logic;
signal bh1112_w42_6_c9 :  std_logic;
signal bh1112_w43_4_c9 :  std_logic;
signal bh1112_w44_3_c9 :  std_logic;
signal bh1112_w45_2_c9 :  std_logic;
signal tile_13_X_c5 :  std_logic_vector(2 downto 0);
signal tile_13_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_13_output_c9 :  std_logic_vector(4 downto 0);
signal tile_13_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w44_4_c9 :  std_logic;
signal bh1112_w45_3_c9 :  std_logic;
signal bh1112_w46_2_c9 :  std_logic;
signal bh1112_w47_1_c9 :  std_logic;
signal bh1112_w48_1_c9 :  std_logic;
signal tile_14_X_c5 :  std_logic_vector(0 downto 0);
signal tile_14_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_14_output_c9 :  std_logic_vector(0 downto 0);
signal tile_14_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_10_c9 :  std_logic;
signal tile_15_X_c5 :  std_logic_vector(1 downto 0);
signal tile_15_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_15_output_c9 :  std_logic_vector(1 downto 0);
signal tile_15_filtered_output_c9 :  unsigned(1-0 downto 0);
signal bh1112_w39_11_c9 :  std_logic;
signal bh1112_w40_6_c9 :  std_logic;
signal tile_16_X_c5 :  std_logic_vector(2 downto 0);
signal tile_16_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_16_output_c9 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w40_7_c9 :  std_logic;
signal bh1112_w41_6_c9 :  std_logic;
signal bh1112_w42_7_c9 :  std_logic;
signal bh1112_w43_5_c9 :  std_logic;
signal bh1112_w44_5_c9 :  std_logic;
signal tile_17_X_c5 :  std_logic_vector(2 downto 0);
signal tile_17_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_17_output_c9 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w43_6_c9 :  std_logic;
signal bh1112_w44_6_c9 :  std_logic;
signal bh1112_w45_4_c9 :  std_logic;
signal bh1112_w46_3_c9 :  std_logic;
signal bh1112_w47_2_c9 :  std_logic;
signal tile_18_X_c5 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_18_output_c9 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w46_4_c9 :  std_logic;
signal bh1112_w47_3_c9 :  std_logic;
signal bh1112_w48_2_c9 :  std_logic;
signal bh1112_w49_1_c9 :  std_logic;
signal bh1112_w50_1_c9 :  std_logic;
signal tile_19_X_c5 :  std_logic_vector(0 downto 0);
signal tile_19_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_19_output_c9 :  std_logic_vector(0 downto 0);
signal tile_19_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_12_c9 :  std_logic;
signal tile_20_X_c5 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_20_output_c9 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w39_13_c9 :  std_logic;
signal bh1112_w40_8_c9 :  std_logic;
signal bh1112_w41_7_c9 :  std_logic;
signal bh1112_w42_8_c9 :  std_logic;
signal bh1112_w43_7_c9 :  std_logic;
signal tile_21_X_c5 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_21_output_c9 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w42_9_c9 :  std_logic;
signal bh1112_w43_8_c9 :  std_logic;
signal bh1112_w44_7_c9 :  std_logic;
signal bh1112_w45_5_c9 :  std_logic;
signal bh1112_w46_5_c9 :  std_logic;
signal tile_22_X_c5 :  std_logic_vector(2 downto 0);
signal tile_22_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_22_output_c9 :  std_logic_vector(4 downto 0);
signal tile_22_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w45_6_c9 :  std_logic;
signal bh1112_w46_6_c9 :  std_logic;
signal bh1112_w47_4_c9 :  std_logic;
signal bh1112_w48_3_c9 :  std_logic;
signal bh1112_w49_2_c9 :  std_logic;
signal tile_23_X_c5 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_23_output_c9 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w48_4_c9 :  std_logic;
signal bh1112_w49_3_c9 :  std_logic;
signal bh1112_w50_2_c9 :  std_logic;
signal bh1112_w51_1_c9 :  std_logic;
signal bh1112_w52_1_c9 :  std_logic;
signal tile_24_X_c5 :  std_logic_vector(16 downto 0);
signal tile_24_Y_c9 :  std_logic_vector(22 downto 0);
signal tile_24_output_c9 :  std_logic_vector(39 downto 0);
signal tile_24_filtered_output_c9 :  unsigned(39-0 downto 0);
signal bh1112_w53_1_c9 :  std_logic;
signal bh1112_w54_1_c9 :  std_logic;
signal bh1112_w55_1_c9 :  std_logic;
signal bh1112_w56_1_c9 :  std_logic;
signal bh1112_w57_1_c9 :  std_logic;
signal bh1112_w58_1_c9 :  std_logic;
signal bh1112_w59_1_c9 :  std_logic;
signal bh1112_w60_1_c9 :  std_logic;
signal bh1112_w61_1_c9 :  std_logic;
signal bh1112_w62_1_c9 :  std_logic;
signal bh1112_w63_1_c9 :  std_logic;
signal bh1112_w64_1_c9 :  std_logic;
signal bh1112_w65_1_c9 :  std_logic;
signal bh1112_w66_1_c9 :  std_logic;
signal bh1112_w67_1_c9 :  std_logic;
signal bh1112_w68_1_c9 :  std_logic;
signal bh1112_w69_1_c9 :  std_logic;
signal bh1112_w70_0_c9 :  std_logic;
signal bh1112_w71_0_c9 :  std_logic;
signal bh1112_w72_0_c9 :  std_logic;
signal bh1112_w73_0_c9 :  std_logic;
signal bh1112_w74_0_c9 :  std_logic;
signal bh1112_w75_0_c9 :  std_logic;
signal bh1112_w76_0_c9, bh1112_w76_0_c10 :  std_logic;
signal bh1112_w77_0_c9 :  std_logic;
signal bh1112_w78_0_c9, bh1112_w78_0_c10 :  std_logic;
signal bh1112_w79_0_c9 :  std_logic;
signal bh1112_w80_0_c9, bh1112_w80_0_c10 :  std_logic;
signal bh1112_w81_0_c9 :  std_logic;
signal bh1112_w82_0_c9, bh1112_w82_0_c10 :  std_logic;
signal bh1112_w83_0_c9 :  std_logic;
signal bh1112_w84_0_c9, bh1112_w84_0_c10 :  std_logic;
signal bh1112_w85_0_c9, bh1112_w85_0_c10 :  std_logic;
signal bh1112_w86_0_c9, bh1112_w86_0_c10 :  std_logic;
signal bh1112_w87_0_c9, bh1112_w87_0_c10 :  std_logic;
signal bh1112_w88_0_c9, bh1112_w88_0_c10 :  std_logic;
signal bh1112_w89_0_c9, bh1112_w89_0_c10 :  std_logic;
signal bh1112_w90_0_c9, bh1112_w90_0_c10 :  std_logic;
signal bh1112_w91_0_c9, bh1112_w91_0_c10 :  std_logic;
signal bh1112_w92_0_c9, bh1112_w92_0_c10 :  std_logic;
signal tile_25_X_c5 :  std_logic_vector(16 downto 0);
signal tile_25_Y_c9 :  std_logic_vector(22 downto 0);
signal tile_25_output_c9 :  std_logic_vector(39 downto 0);
signal tile_25_filtered_output_c9 :  unsigned(39-0 downto 0);
signal bh1112_w36_1_c9 :  std_logic;
signal bh1112_w37_1_c9 :  std_logic;
signal bh1112_w38_1_c9 :  std_logic;
signal bh1112_w39_14_c9 :  std_logic;
signal bh1112_w40_9_c9 :  std_logic;
signal bh1112_w41_8_c9 :  std_logic;
signal bh1112_w42_10_c9 :  std_logic;
signal bh1112_w43_9_c9 :  std_logic;
signal bh1112_w44_8_c9 :  std_logic;
signal bh1112_w45_7_c9 :  std_logic;
signal bh1112_w46_7_c9 :  std_logic;
signal bh1112_w47_5_c9 :  std_logic;
signal bh1112_w48_5_c9 :  std_logic;
signal bh1112_w49_4_c9 :  std_logic;
signal bh1112_w50_3_c9 :  std_logic;
signal bh1112_w51_2_c9 :  std_logic;
signal bh1112_w52_2_c9 :  std_logic;
signal bh1112_w53_2_c9 :  std_logic;
signal bh1112_w54_2_c9 :  std_logic;
signal bh1112_w55_2_c9 :  std_logic;
signal bh1112_w56_2_c9 :  std_logic;
signal bh1112_w57_2_c9 :  std_logic;
signal bh1112_w58_2_c9 :  std_logic;
signal bh1112_w59_2_c9 :  std_logic;
signal bh1112_w60_2_c9 :  std_logic;
signal bh1112_w61_2_c9, bh1112_w61_2_c10 :  std_logic;
signal bh1112_w62_2_c9 :  std_logic;
signal bh1112_w63_2_c9, bh1112_w63_2_c10 :  std_logic;
signal bh1112_w64_2_c9 :  std_logic;
signal bh1112_w65_2_c9, bh1112_w65_2_c10 :  std_logic;
signal bh1112_w66_2_c9 :  std_logic;
signal bh1112_w67_2_c9, bh1112_w67_2_c10 :  std_logic;
signal bh1112_w68_2_c9 :  std_logic;
signal bh1112_w69_2_c9, bh1112_w69_2_c10 :  std_logic;
signal bh1112_w70_1_c9 :  std_logic;
signal bh1112_w71_1_c9 :  std_logic;
signal bh1112_w72_1_c9 :  std_logic;
signal bh1112_w73_1_c9 :  std_logic;
signal bh1112_w74_1_c9 :  std_logic;
signal bh1112_w75_1_c9 :  std_logic;
signal tile_26_X_c5 :  std_logic_vector(0 downto 0);
signal tile_26_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_26_output_c9 :  std_logic_vector(0 downto 0);
signal tile_26_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_15_c9 :  std_logic;
signal tile_27_X_c5 :  std_logic_vector(0 downto 0);
signal tile_27_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_27_output_c9 :  std_logic_vector(0 downto 0);
signal tile_27_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_16_c9 :  std_logic;
signal tile_28_X_c5 :  std_logic_vector(1 downto 0);
signal tile_28_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_28_output_c9 :  std_logic_vector(3 downto 0);
signal tile_28_filtered_output_c9 :  unsigned(3-0 downto 0);
signal bh1112_w39_17_c9 :  std_logic;
signal bh1112_w40_10_c9 :  std_logic;
signal bh1112_w41_9_c9 :  std_logic;
signal bh1112_w42_11_c9 :  std_logic;
signal tile_29_X_c5 :  std_logic_vector(0 downto 0);
signal tile_29_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_29_output_c9 :  std_logic_vector(0 downto 0);
signal tile_29_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_18_c9 :  std_logic;
signal tile_30_X_c5 :  std_logic_vector(1 downto 0);
signal tile_30_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_30_output_c9 :  std_logic_vector(1 downto 0);
signal tile_30_filtered_output_c9 :  unsigned(1-0 downto 0);
signal bh1112_w39_19_c9 :  std_logic;
signal bh1112_w40_11_c9 :  std_logic;
signal tile_31_X_c5 :  std_logic_vector(2 downto 0);
signal tile_31_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_31_output_c9 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w40_12_c9 :  std_logic;
signal bh1112_w41_10_c9 :  std_logic;
signal bh1112_w42_12_c9 :  std_logic;
signal bh1112_w43_10_c9 :  std_logic;
signal bh1112_w44_9_c9 :  std_logic;
signal tile_32_X_c5 :  std_logic_vector(0 downto 0);
signal tile_32_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_32_output_c9 :  std_logic_vector(0 downto 0);
signal tile_32_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_20_c9 :  std_logic;
signal tile_33_X_c5 :  std_logic_vector(2 downto 0);
signal tile_33_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_33_output_c9 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w39_21_c9 :  std_logic;
signal bh1112_w40_13_c9 :  std_logic;
signal bh1112_w41_11_c9 :  std_logic;
signal bh1112_w42_13_c9 :  std_logic;
signal bh1112_w43_11_c9 :  std_logic;
signal tile_34_X_c5 :  std_logic_vector(2 downto 0);
signal tile_34_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_34_output_c9 :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w42_14_c9 :  std_logic;
signal bh1112_w43_12_c9 :  std_logic;
signal bh1112_w44_10_c9 :  std_logic;
signal bh1112_w45_8_c9 :  std_logic;
signal bh1112_w46_8_c9 :  std_logic;
signal tile_35_X_c5 :  std_logic_vector(0 downto 0);
signal tile_35_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_35_output_c9 :  std_logic_vector(0 downto 0);
signal tile_35_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_22_c9 :  std_logic;
signal tile_36_X_c5 :  std_logic_vector(1 downto 0);
signal tile_36_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_36_output_c9 :  std_logic_vector(3 downto 0);
signal tile_36_filtered_output_c9 :  unsigned(3-0 downto 0);
signal bh1112_w39_23_c9 :  std_logic;
signal bh1112_w40_14_c9 :  std_logic;
signal bh1112_w41_12_c9 :  std_logic;
signal bh1112_w42_15_c9 :  std_logic;
signal tile_37_X_c5 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_37_output_c9 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w41_13_c9 :  std_logic;
signal bh1112_w42_16_c9 :  std_logic;
signal bh1112_w43_13_c9 :  std_logic;
signal bh1112_w44_11_c9 :  std_logic;
signal bh1112_w45_9_c9 :  std_logic;
signal tile_38_X_c5 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_38_output_c9 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w44_12_c9 :  std_logic;
signal bh1112_w45_10_c9 :  std_logic;
signal bh1112_w46_9_c9 :  std_logic;
signal bh1112_w47_6_c9 :  std_logic;
signal bh1112_w48_6_c9 :  std_logic;
signal tile_39_X_c5 :  std_logic_vector(0 downto 0);
signal tile_39_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_39_output_c9 :  std_logic_vector(0 downto 0);
signal tile_39_filtered_output_c9 :  unsigned(0-0 downto 0);
signal bh1112_w39_24_c9 :  std_logic;
signal tile_40_X_c5 :  std_logic_vector(1 downto 0);
signal tile_40_Y_c9 :  std_logic_vector(0 downto 0);
signal tile_40_output_c9 :  std_logic_vector(1 downto 0);
signal tile_40_filtered_output_c9 :  unsigned(1-0 downto 0);
signal bh1112_w39_25_c9 :  std_logic;
signal bh1112_w40_15_c9 :  std_logic;
signal tile_41_X_c5 :  std_logic_vector(2 downto 0);
signal tile_41_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_41_output_c9 :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w40_16_c9 :  std_logic;
signal bh1112_w41_14_c9 :  std_logic;
signal bh1112_w42_17_c9 :  std_logic;
signal bh1112_w43_14_c9 :  std_logic;
signal bh1112_w44_13_c9 :  std_logic;
signal tile_42_X_c5 :  std_logic_vector(2 downto 0);
signal tile_42_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_42_output_c9 :  std_logic_vector(4 downto 0);
signal tile_42_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w43_15_c9 :  std_logic;
signal bh1112_w44_14_c9 :  std_logic;
signal bh1112_w45_11_c9 :  std_logic;
signal bh1112_w46_10_c9 :  std_logic;
signal bh1112_w47_7_c9 :  std_logic;
signal tile_43_X_c5 :  std_logic_vector(2 downto 0);
signal tile_43_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_43_output_c9 :  std_logic_vector(4 downto 0);
signal tile_43_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w46_11_c9 :  std_logic;
signal bh1112_w47_8_c9 :  std_logic;
signal bh1112_w48_7_c9 :  std_logic;
signal bh1112_w49_5_c9 :  std_logic;
signal bh1112_w50_4_c9 :  std_logic;
signal tile_44_X_c5 :  std_logic_vector(2 downto 0);
signal tile_44_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_44_output_c9 :  std_logic_vector(4 downto 0);
signal tile_44_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w39_26_c9 :  std_logic;
signal bh1112_w40_17_c9 :  std_logic;
signal bh1112_w41_15_c9 :  std_logic;
signal bh1112_w42_18_c9 :  std_logic;
signal bh1112_w43_16_c9 :  std_logic;
signal tile_45_X_c5 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_45_output_c9 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w42_19_c9 :  std_logic;
signal bh1112_w43_17_c9 :  std_logic;
signal bh1112_w44_15_c9 :  std_logic;
signal bh1112_w45_12_c9 :  std_logic;
signal bh1112_w46_12_c9 :  std_logic;
signal tile_46_X_c5 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_46_output_c9 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w45_13_c9 :  std_logic;
signal bh1112_w46_13_c9 :  std_logic;
signal bh1112_w47_9_c9 :  std_logic;
signal bh1112_w48_8_c9 :  std_logic;
signal bh1112_w49_6_c9, bh1112_w49_6_c10 :  std_logic;
signal tile_47_X_c5 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_47_output_c9 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w48_9_c9, bh1112_w48_9_c10 :  std_logic;
signal bh1112_w49_7_c9 :  std_logic;
signal bh1112_w50_5_c9 :  std_logic;
signal bh1112_w51_3_c9 :  std_logic;
signal bh1112_w52_3_c9 :  std_logic;
signal tile_48_X_c5 :  std_logic_vector(2 downto 0);
signal tile_48_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_48_output_c9 :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w41_16_c9 :  std_logic;
signal bh1112_w42_20_c9 :  std_logic;
signal bh1112_w43_18_c9 :  std_logic;
signal bh1112_w44_16_c9 :  std_logic;
signal bh1112_w45_14_c9 :  std_logic;
signal tile_49_X_c5 :  std_logic_vector(2 downto 0);
signal tile_49_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_49_output_c9 :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w44_17_c9 :  std_logic;
signal bh1112_w45_15_c9 :  std_logic;
signal bh1112_w46_14_c9 :  std_logic;
signal bh1112_w47_10_c9 :  std_logic;
signal bh1112_w48_10_c9 :  std_logic;
signal tile_50_X_c5 :  std_logic_vector(2 downto 0);
signal tile_50_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_50_output_c9 :  std_logic_vector(4 downto 0);
signal tile_50_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w47_11_c9 :  std_logic;
signal bh1112_w48_11_c9 :  std_logic;
signal bh1112_w49_8_c9 :  std_logic;
signal bh1112_w50_6_c9 :  std_logic;
signal bh1112_w51_4_c9 :  std_logic;
signal tile_51_X_c5 :  std_logic_vector(2 downto 0);
signal tile_51_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_51_output_c9 :  std_logic_vector(4 downto 0);
signal tile_51_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w50_7_c9 :  std_logic;
signal bh1112_w51_5_c9 :  std_logic;
signal bh1112_w52_4_c9 :  std_logic;
signal bh1112_w53_3_c9 :  std_logic;
signal bh1112_w54_3_c9 :  std_logic;
signal tile_52_X_c5 :  std_logic_vector(2 downto 0);
signal tile_52_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_52_output_c9 :  std_logic_vector(4 downto 0);
signal tile_52_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w43_19_c9 :  std_logic;
signal bh1112_w44_18_c9 :  std_logic;
signal bh1112_w45_16_c9 :  std_logic;
signal bh1112_w46_15_c9 :  std_logic;
signal bh1112_w47_12_c9 :  std_logic;
signal tile_53_X_c5 :  std_logic_vector(2 downto 0);
signal tile_53_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_53_output_c9 :  std_logic_vector(4 downto 0);
signal tile_53_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w46_16_c9 :  std_logic;
signal bh1112_w47_13_c9 :  std_logic;
signal bh1112_w48_12_c9 :  std_logic;
signal bh1112_w49_9_c9 :  std_logic;
signal bh1112_w50_8_c9 :  std_logic;
signal tile_54_X_c5 :  std_logic_vector(2 downto 0);
signal tile_54_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_54_output_c9 :  std_logic_vector(4 downto 0);
signal tile_54_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w49_10_c9 :  std_logic;
signal bh1112_w50_9_c9 :  std_logic;
signal bh1112_w51_6_c9 :  std_logic;
signal bh1112_w52_5_c9 :  std_logic;
signal bh1112_w53_4_c9 :  std_logic;
signal tile_55_X_c5 :  std_logic_vector(2 downto 0);
signal tile_55_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_55_output_c9 :  std_logic_vector(4 downto 0);
signal tile_55_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w52_6_c9 :  std_logic;
signal bh1112_w53_5_c9 :  std_logic;
signal bh1112_w54_4_c9 :  std_logic;
signal bh1112_w55_3_c9 :  std_logic;
signal bh1112_w56_3_c9 :  std_logic;
signal tile_56_X_c5 :  std_logic_vector(2 downto 0);
signal tile_56_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_56_output_c9 :  std_logic_vector(4 downto 0);
signal tile_56_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w45_17_c9 :  std_logic;
signal bh1112_w46_17_c9 :  std_logic;
signal bh1112_w47_14_c9 :  std_logic;
signal bh1112_w48_13_c9 :  std_logic;
signal bh1112_w49_11_c9 :  std_logic;
signal tile_57_X_c5 :  std_logic_vector(2 downto 0);
signal tile_57_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_57_output_c9 :  std_logic_vector(4 downto 0);
signal tile_57_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w48_14_c9 :  std_logic;
signal bh1112_w49_12_c9 :  std_logic;
signal bh1112_w50_10_c9 :  std_logic;
signal bh1112_w51_7_c9 :  std_logic;
signal bh1112_w52_7_c9 :  std_logic;
signal tile_58_X_c5 :  std_logic_vector(2 downto 0);
signal tile_58_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_58_output_c9 :  std_logic_vector(4 downto 0);
signal tile_58_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w51_8_c9 :  std_logic;
signal bh1112_w52_8_c9 :  std_logic;
signal bh1112_w53_6_c9, bh1112_w53_6_c10 :  std_logic;
signal bh1112_w54_5_c9 :  std_logic;
signal bh1112_w55_4_c9 :  std_logic;
signal tile_59_X_c5 :  std_logic_vector(2 downto 0);
signal tile_59_Y_c9 :  std_logic_vector(1 downto 0);
signal tile_59_output_c9 :  std_logic_vector(4 downto 0);
signal tile_59_filtered_output_c9 :  unsigned(4-0 downto 0);
signal bh1112_w54_6_c9 :  std_logic;
signal bh1112_w55_5_c9 :  std_logic;
signal bh1112_w56_4_c9, bh1112_w56_4_c10 :  std_logic;
signal bh1112_w57_3_c9 :  std_logic;
signal bh1112_w58_3_c9 :  std_logic;
signal bh1112_w39_27_c0, bh1112_w39_27_c1, bh1112_w39_27_c2, bh1112_w39_27_c3, bh1112_w39_27_c4, bh1112_w39_27_c5, bh1112_w39_27_c6, bh1112_w39_27_c7, bh1112_w39_27_c8, bh1112_w39_27_c9 :  std_logic;
signal bh1112_w40_18_c0, bh1112_w40_18_c1, bh1112_w40_18_c2, bh1112_w40_18_c3, bh1112_w40_18_c4, bh1112_w40_18_c5, bh1112_w40_18_c6, bh1112_w40_18_c7, bh1112_w40_18_c8, bh1112_w40_18_c9 :  std_logic;
signal bh1112_w41_17_c0, bh1112_w41_17_c1, bh1112_w41_17_c2, bh1112_w41_17_c3, bh1112_w41_17_c4, bh1112_w41_17_c5, bh1112_w41_17_c6, bh1112_w41_17_c7, bh1112_w41_17_c8, bh1112_w41_17_c9 :  std_logic;
signal bh1112_w42_21_c0, bh1112_w42_21_c1, bh1112_w42_21_c2, bh1112_w42_21_c3, bh1112_w42_21_c4, bh1112_w42_21_c5, bh1112_w42_21_c6, bh1112_w42_21_c7, bh1112_w42_21_c8, bh1112_w42_21_c9 :  std_logic;
signal bh1112_w43_20_c0, bh1112_w43_20_c1, bh1112_w43_20_c2, bh1112_w43_20_c3, bh1112_w43_20_c4, bh1112_w43_20_c5, bh1112_w43_20_c6, bh1112_w43_20_c7, bh1112_w43_20_c8, bh1112_w43_20_c9 :  std_logic;
signal bh1112_w44_19_c0, bh1112_w44_19_c1, bh1112_w44_19_c2, bh1112_w44_19_c3, bh1112_w44_19_c4, bh1112_w44_19_c5, bh1112_w44_19_c6, bh1112_w44_19_c7, bh1112_w44_19_c8, bh1112_w44_19_c9 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1356_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1356_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w36_2_c10 :  std_logic;
signal bh1112_w37_2_c10 :  std_logic;
signal bh1112_w38_2_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_copy1357_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_copy1357_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1360_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w38_3_c10 :  std_logic;
signal bh1112_w39_28_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_copy1361_c9, Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_copy1361_c10 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1364_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w39_29_c10 :  std_logic;
signal bh1112_w40_19_c10 :  std_logic;
signal bh1112_w41_18_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_copy1365_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_copy1365_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1366_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w39_30_c10 :  std_logic;
signal bh1112_w40_20_c10 :  std_logic;
signal bh1112_w41_19_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_copy1367_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_copy1367_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1368_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1368_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w39_31_c9, bh1112_w39_31_c10 :  std_logic;
signal bh1112_w40_21_c9, bh1112_w40_21_c10 :  std_logic;
signal bh1112_w41_20_c9, bh1112_w41_20_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1368_Out0_copy1369_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1370_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1370_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w39_32_c9, bh1112_w39_32_c10 :  std_logic;
signal bh1112_w40_22_c9, bh1112_w40_22_c10 :  std_logic;
signal bh1112_w41_21_c9, bh1112_w41_21_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1370_Out0_copy1371_c9 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1374_In0_c9 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1374_In1_c9 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w39_33_c10 :  std_logic;
signal bh1112_w40_23_c10 :  std_logic;
signal bh1112_w41_22_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_copy1375_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_copy1375_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1376_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1376_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w40_24_c9, bh1112_w40_24_c10 :  std_logic;
signal bh1112_w41_23_c9, bh1112_w41_23_c10 :  std_logic;
signal bh1112_w42_22_c9, bh1112_w42_22_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1376_Out0_copy1377_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1378_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1378_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w40_25_c9, bh1112_w40_25_c10 :  std_logic;
signal bh1112_w41_24_c9, bh1112_w41_24_c10 :  std_logic;
signal bh1112_w42_23_c9, bh1112_w42_23_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1378_Out0_copy1379_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1380_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w40_26_c10 :  std_logic;
signal bh1112_w41_25_c10 :  std_logic;
signal bh1112_w42_24_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_copy1381_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_copy1381_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1382_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1382_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w41_26_c9, bh1112_w41_26_c10 :  std_logic;
signal bh1112_w42_25_c9, bh1112_w42_25_c10 :  std_logic;
signal bh1112_w43_21_c9, bh1112_w43_21_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1382_Out0_copy1383_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1384_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w41_27_c10 :  std_logic;
signal bh1112_w42_26_c10 :  std_logic;
signal bh1112_w43_22_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_copy1385_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_copy1385_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1386_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w41_28_c10 :  std_logic;
signal bh1112_w42_27_c10 :  std_logic;
signal bh1112_w43_23_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_copy1387_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_copy1387_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1388_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w42_28_c10 :  std_logic;
signal bh1112_w43_24_c10 :  std_logic;
signal bh1112_w44_20_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_copy1389_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_copy1389_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1390_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1390_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w42_29_c9, bh1112_w42_29_c10 :  std_logic;
signal bh1112_w43_25_c9, bh1112_w43_25_c10 :  std_logic;
signal bh1112_w44_21_c9, bh1112_w44_21_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1390_Out0_copy1391_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1392_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w42_30_c10 :  std_logic;
signal bh1112_w43_26_c10 :  std_logic;
signal bh1112_w44_22_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_copy1393_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_copy1393_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In0_c9 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c0, Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c1, Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c2, Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c3, Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c4, Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c5, Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c6, Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c7, Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c8, Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c9 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1394_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w42_31_c9, bh1112_w42_31_c10 :  std_logic;
signal bh1112_w43_27_c9, bh1112_w43_27_c10 :  std_logic;
signal bh1112_w44_23_c9 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1394_Out0_copy1395_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1396_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1396_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w43_28_c9, bh1112_w43_28_c10 :  std_logic;
signal bh1112_w44_24_c9, bh1112_w44_24_c10 :  std_logic;
signal bh1112_w45_18_c9, bh1112_w45_18_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1396_Out0_copy1397_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1398_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1398_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w43_29_c9, bh1112_w43_29_c10 :  std_logic;
signal bh1112_w44_25_c9 :  std_logic;
signal bh1112_w45_19_c9, bh1112_w45_19_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1398_Out0_copy1399_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1400_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w43_30_c10 :  std_logic;
signal bh1112_w44_26_c10 :  std_logic;
signal bh1112_w45_20_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_copy1401_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_copy1401_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1402_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1402_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1402_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w43_31_c9, bh1112_w43_31_c10 :  std_logic;
signal bh1112_w44_27_c9 :  std_logic;
signal bh1112_w45_21_c9, bh1112_w45_21_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1402_Out0_copy1403_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1404_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w44_28_c10 :  std_logic;
signal bh1112_w45_22_c10 :  std_logic;
signal bh1112_w46_18_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_copy1405_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_copy1405_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1406_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1406_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w44_29_c9 :  std_logic;
signal bh1112_w45_23_c9, bh1112_w45_23_c10 :  std_logic;
signal bh1112_w46_19_c9, bh1112_w46_19_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1406_Out0_copy1407_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1408_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w44_30_c10 :  std_logic;
signal bh1112_w45_24_c10 :  std_logic;
signal bh1112_w46_20_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_copy1409_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_copy1409_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1410_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1410_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w45_25_c9, bh1112_w45_25_c10 :  std_logic;
signal bh1112_w46_21_c9, bh1112_w46_21_c10 :  std_logic;
signal bh1112_w47_15_c9, bh1112_w47_15_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1410_Out0_copy1411_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1412_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w45_26_c10 :  std_logic;
signal bh1112_w46_22_c10 :  std_logic;
signal bh1112_w47_16_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_copy1413_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_copy1413_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1414_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w45_27_c10 :  std_logic;
signal bh1112_w46_23_c10 :  std_logic;
signal bh1112_w47_17_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_copy1415_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_copy1415_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1416_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w46_24_c10 :  std_logic;
signal bh1112_w47_18_c10 :  std_logic;
signal bh1112_w48_15_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_copy1417_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_copy1417_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1418_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1418_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w46_25_c9, bh1112_w46_25_c10 :  std_logic;
signal bh1112_w47_19_c9, bh1112_w47_19_c10 :  std_logic;
signal bh1112_w48_16_c9, bh1112_w48_16_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1418_Out0_copy1419_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1420_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w46_26_c10 :  std_logic;
signal bh1112_w47_20_c10 :  std_logic;
signal bh1112_w48_17_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_copy1421_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_copy1421_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1422_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1422_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w47_21_c9, bh1112_w47_21_c10 :  std_logic;
signal bh1112_w48_18_c9, bh1112_w48_18_c10 :  std_logic;
signal bh1112_w49_13_c9, bh1112_w49_13_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1422_Out0_copy1423_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1424_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w47_22_c10 :  std_logic;
signal bh1112_w48_19_c10 :  std_logic;
signal bh1112_w49_14_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_copy1425_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_copy1425_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1426_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1426_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w47_23_c10 :  std_logic;
signal bh1112_w48_20_c10 :  std_logic;
signal bh1112_w49_15_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_copy1427_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_copy1427_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1428_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1428_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w48_21_c9, bh1112_w48_21_c10 :  std_logic;
signal bh1112_w49_16_c9, bh1112_w49_16_c10 :  std_logic;
signal bh1112_w50_11_c9, bh1112_w50_11_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1428_Out0_copy1429_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1430_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w48_22_c10 :  std_logic;
signal bh1112_w49_17_c10 :  std_logic;
signal bh1112_w50_12_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_copy1431_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_copy1431_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1432_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w49_18_c10 :  std_logic;
signal bh1112_w50_13_c10 :  std_logic;
signal bh1112_w51_9_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_copy1433_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_copy1433_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1434_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1434_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w49_19_c9, bh1112_w49_19_c10 :  std_logic;
signal bh1112_w50_14_c9, bh1112_w50_14_c10 :  std_logic;
signal bh1112_w51_10_c9, bh1112_w51_10_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1434_Out0_copy1435_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1436_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w50_15_c10 :  std_logic;
signal bh1112_w51_11_c10 :  std_logic;
signal bh1112_w52_9_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_copy1437_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_copy1437_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1438_In0_c9 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1438_In1_c9 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w50_16_c10 :  std_logic;
signal bh1112_w51_12_c10 :  std_logic;
signal bh1112_w52_10_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_copy1439_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_copy1439_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1440_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1440_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w50_17_c10 :  std_logic;
signal bh1112_w51_13_c10 :  std_logic;
signal bh1112_w52_11_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_copy1441_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_copy1441_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1442_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1442_Out0_c9 :  std_logic_vector(2 downto 0);
signal bh1112_w51_14_c9, bh1112_w51_14_c10 :  std_logic;
signal bh1112_w52_12_c9, bh1112_w52_12_c10 :  std_logic;
signal bh1112_w53_7_c9, bh1112_w53_7_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1442_Out0_copy1443_c9 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1444_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w52_13_c10 :  std_logic;
signal bh1112_w53_8_c10 :  std_logic;
signal bh1112_w54_7_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_copy1445_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_copy1445_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1446_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1446_Out0_c9 :  std_logic_vector(1 downto 0);
signal bh1112_w52_14_c9, bh1112_w52_14_c10 :  std_logic;
signal bh1112_w53_9_c9, bh1112_w53_9_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1446_Out0_copy1447_c9 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1448_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w53_10_c10 :  std_logic;
signal bh1112_w54_8_c10 :  std_logic;
signal bh1112_w55_6_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_copy1449_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_copy1449_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1450_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w54_9_c10 :  std_logic;
signal bh1112_w55_7_c10 :  std_logic;
signal bh1112_w56_5_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_copy1451_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_copy1451_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1452_In0_c9 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w55_8_c10 :  std_logic;
signal bh1112_w56_6_c10 :  std_logic;
signal bh1112_w57_4_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_copy1453_c9, Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_copy1453_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1454_In0_c9 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1454_In1_c9 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w56_7_c10 :  std_logic;
signal bh1112_w57_5_c10 :  std_logic;
signal bh1112_w58_4_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_copy1455_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_copy1455_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1456_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w57_6_c10 :  std_logic;
signal bh1112_w58_5_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_copy1457_c9, Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_copy1457_c10 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In0_c9 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c0, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c1, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c2, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c3, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c4, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c5, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c6, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c7, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c8, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c9 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w58_6_c10 :  std_logic;
signal bh1112_w59_3_c10 :  std_logic;
signal bh1112_w60_3_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_copy1459_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_copy1459_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1460_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w59_4_c10 :  std_logic;
signal bh1112_w60_4_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_copy1461_c9, Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_copy1461_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1462_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1462_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w60_5_c10 :  std_logic;
signal bh1112_w61_3_c10 :  std_logic;
signal bh1112_w62_3_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_copy1463_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_copy1463_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1464_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1464_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w62_4_c10 :  std_logic;
signal bh1112_w63_3_c10 :  std_logic;
signal bh1112_w64_3_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_copy1465_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_copy1465_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1466_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1466_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w64_4_c10 :  std_logic;
signal bh1112_w65_3_c10 :  std_logic;
signal bh1112_w66_3_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_copy1467_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_copy1467_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1468_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1468_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w66_4_c10 :  std_logic;
signal bh1112_w67_3_c10 :  std_logic;
signal bh1112_w68_3_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_copy1469_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_copy1469_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1470_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1470_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w68_4_c10 :  std_logic;
signal bh1112_w69_3_c10 :  std_logic;
signal bh1112_w70_2_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_copy1471_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_copy1471_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1472_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1472_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w70_3_c10 :  std_logic;
signal bh1112_w71_2_c10 :  std_logic;
signal bh1112_w72_2_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_copy1473_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_copy1473_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1474_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1474_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w72_3_c10 :  std_logic;
signal bh1112_w73_2_c10 :  std_logic;
signal bh1112_w74_2_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_copy1475_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_copy1475_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1476_In0_c9 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1476_In1_c9 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w74_3_c10 :  std_logic;
signal bh1112_w75_2_c10 :  std_logic;
signal bh1112_w76_1_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_copy1477_c9, Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_copy1477_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1478_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1478_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1478_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w37_3_c10 :  std_logic;
signal bh1112_w38_4_c10 :  std_logic;
signal bh1112_w39_34_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1478_Out0_copy1479_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1480_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1480_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w39_35_c10 :  std_logic;
signal bh1112_w40_27_c10 :  std_logic;
signal bh1112_w41_29_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1480_Out0_copy1481_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1482_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1482_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w40_28_c10 :  std_logic;
signal bh1112_w41_30_c10 :  std_logic;
signal bh1112_w42_32_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1482_Out0_copy1483_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1484_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1484_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1484_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w40_29_c10 :  std_logic;
signal bh1112_w41_31_c10 :  std_logic;
signal bh1112_w42_33_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1484_Out0_copy1485_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1486_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1486_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w41_32_c10 :  std_logic;
signal bh1112_w42_34_c10 :  std_logic;
signal bh1112_w43_32_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1486_Out0_copy1487_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1488_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1488_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1488_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w41_33_c10 :  std_logic;
signal bh1112_w42_35_c10 :  std_logic;
signal bh1112_w43_33_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1488_Out0_copy1489_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1490_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1490_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w42_36_c10 :  std_logic;
signal bh1112_w43_34_c10 :  std_logic;
signal bh1112_w44_31_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1490_Out0_copy1491_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1492_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1492_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w42_37_c10 :  std_logic;
signal bh1112_w43_35_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1492_Out0_copy1493_c10 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1494_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1494_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w43_36_c10 :  std_logic;
signal bh1112_w44_32_c10 :  std_logic;
signal bh1112_w45_28_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1494_Out0_copy1495_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1496_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1496_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1496_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w43_37_c10 :  std_logic;
signal bh1112_w44_33_c10 :  std_logic;
signal bh1112_w45_29_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1496_Out0_copy1497_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1498_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1498_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w44_34_c10 :  std_logic;
signal bh1112_w45_30_c10 :  std_logic;
signal bh1112_w46_27_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1498_Out0_copy1499_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1500_In0_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1500_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1500_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1500_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w44_35_c10 :  std_logic;
signal bh1112_w45_31_c10 :  std_logic;
signal bh1112_w46_28_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1500_Out0_copy1501_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1502_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1502_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w45_32_c10 :  std_logic;
signal bh1112_w46_29_c10 :  std_logic;
signal bh1112_w47_24_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1502_Out0_copy1503_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1504_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1504_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1504_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w45_33_c10 :  std_logic;
signal bh1112_w46_30_c10 :  std_logic;
signal bh1112_w47_25_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1504_Out0_copy1505_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1506_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1506_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w46_31_c10 :  std_logic;
signal bh1112_w47_26_c10 :  std_logic;
signal bh1112_w48_23_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1506_Out0_copy1507_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1508_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1508_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w47_27_c10 :  std_logic;
signal bh1112_w48_24_c10 :  std_logic;
signal bh1112_w49_20_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1508_Out0_copy1509_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1510_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1510_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1510_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w47_28_c10 :  std_logic;
signal bh1112_w48_25_c10 :  std_logic;
signal bh1112_w49_21_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1510_Out0_copy1511_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1512_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1512_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w48_26_c10 :  std_logic;
signal bh1112_w49_22_c10 :  std_logic;
signal bh1112_w50_18_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1512_Out0_copy1513_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1514_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1514_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w49_23_c10 :  std_logic;
signal bh1112_w50_19_c10 :  std_logic;
signal bh1112_w51_15_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1514_Out0_copy1515_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1516_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1516_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1516_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w49_24_c10 :  std_logic;
signal bh1112_w50_20_c10 :  std_logic;
signal bh1112_w51_16_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1516_Out0_copy1517_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1518_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1518_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w50_21_c10 :  std_logic;
signal bh1112_w51_17_c10 :  std_logic;
signal bh1112_w52_15_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1518_Out0_copy1519_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1520_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1520_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w51_18_c10 :  std_logic;
signal bh1112_w52_16_c10 :  std_logic;
signal bh1112_w53_11_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1520_Out0_copy1521_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1522_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1522_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w52_17_c10 :  std_logic;
signal bh1112_w53_12_c10 :  std_logic;
signal bh1112_w54_10_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1522_Out0_copy1523_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1524_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1524_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1524_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1524_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w53_13_c10 :  std_logic;
signal bh1112_w54_11_c10 :  std_logic;
signal bh1112_w55_9_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1524_Out0_copy1525_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1526_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1526_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1526_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w54_12_c10 :  std_logic;
signal bh1112_w55_10_c10 :  std_logic;
signal bh1112_w56_8_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1526_Out0_copy1527_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c0, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c1, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c2, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c3, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c4, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c5, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c6, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c7, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c8, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1528_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w56_9_c10 :  std_logic;
signal bh1112_w57_7_c10 :  std_logic;
signal bh1112_w58_7_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1528_Out0_copy1529_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1530_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1530_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w57_8_c10 :  std_logic;
signal bh1112_w58_8_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1530_Out0_copy1531_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1532_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1532_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1532_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w58_9_c10 :  std_logic;
signal bh1112_w59_5_c10 :  std_logic;
signal bh1112_w60_6_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1532_Out0_copy1533_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1534_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1534_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1534_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w60_7_c10 :  std_logic;
signal bh1112_w61_4_c10 :  std_logic;
signal bh1112_w62_5_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1534_Out0_copy1535_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1536_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1536_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1536_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w62_6_c10 :  std_logic;
signal bh1112_w63_4_c10 :  std_logic;
signal bh1112_w64_5_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1536_Out0_copy1537_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1538_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1538_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1538_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w64_6_c10 :  std_logic;
signal bh1112_w65_4_c10 :  std_logic;
signal bh1112_w66_5_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1538_Out0_copy1539_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1540_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1540_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1540_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w66_6_c10 :  std_logic;
signal bh1112_w67_4_c10 :  std_logic;
signal bh1112_w68_5_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1540_Out0_copy1541_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1542_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1542_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1542_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w68_6_c10 :  std_logic;
signal bh1112_w69_4_c10 :  std_logic;
signal bh1112_w70_4_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1542_Out0_copy1543_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1544_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1544_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1544_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w70_5_c10 :  std_logic;
signal bh1112_w71_3_c10 :  std_logic;
signal bh1112_w72_4_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1544_Out0_copy1545_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1546_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1546_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1546_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w72_5_c10 :  std_logic;
signal bh1112_w73_3_c10 :  std_logic;
signal bh1112_w74_4_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1546_Out0_copy1547_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1548_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1548_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1548_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w74_5_c10 :  std_logic;
signal bh1112_w75_3_c10 :  std_logic;
signal bh1112_w76_2_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1548_Out0_copy1549_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1550_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1550_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1550_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1550_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w76_3_c10 :  std_logic;
signal bh1112_w77_1_c10 :  std_logic;
signal bh1112_w78_1_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1550_Out0_copy1551_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1552_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1552_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1552_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w38_5_c10 :  std_logic;
signal bh1112_w39_36_c10 :  std_logic;
signal bh1112_w40_30_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1552_Out0_copy1553_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1554_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1554_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w40_31_c10 :  std_logic;
signal bh1112_w41_34_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1554_Out0_copy1555_c10 :  std_logic_vector(1 downto 0);
signal Compressor_5_3_Freq300_uid1557_bh1112_uid1558_In0_c10 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid1557_bh1112_uid1558_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w41_35_c10 :  std_logic;
signal bh1112_w42_38_c10 :  std_logic;
signal bh1112_w43_38_c10 :  std_logic;
signal Compressor_5_3_Freq300_uid1557_bh1112_uid1558_Out0_copy1559_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1560_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1560_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w42_39_c10 :  std_logic;
signal bh1112_w43_39_c10 :  std_logic;
signal bh1112_w44_36_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1560_Out0_copy1561_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1562_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1562_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w43_40_c10 :  std_logic;
signal bh1112_w44_37_c10 :  std_logic;
signal bh1112_w45_34_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1562_Out0_copy1563_c10 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid1557_bh1112_uid1564_In0_c10 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid1557_bh1112_uid1564_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w44_38_c10 :  std_logic;
signal bh1112_w45_35_c10 :  std_logic;
signal bh1112_w46_32_c10 :  std_logic;
signal Compressor_5_3_Freq300_uid1557_bh1112_uid1564_Out0_copy1565_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1566_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1566_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w45_36_c10 :  std_logic;
signal bh1112_w46_33_c10 :  std_logic;
signal bh1112_w47_29_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1566_Out0_copy1567_c10 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1568_In0_c10 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1568_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w46_34_c10 :  std_logic;
signal bh1112_w47_30_c10 :  std_logic;
signal bh1112_w48_27_c10 :  std_logic;
signal Compressor_6_3_Freq300_uid1363_bh1112_uid1568_Out0_copy1569_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1570_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1570_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1570_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w47_31_c10 :  std_logic;
signal bh1112_w48_28_c10 :  std_logic;
signal bh1112_w49_25_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1570_Out0_copy1571_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1572_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1572_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1572_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w48_29_c10 :  std_logic;
signal bh1112_w49_26_c10 :  std_logic;
signal bh1112_w50_22_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1572_Out0_copy1573_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1574_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1574_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1574_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w49_27_c10 :  std_logic;
signal bh1112_w50_23_c10 :  std_logic;
signal bh1112_w51_19_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1574_Out0_copy1575_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1576_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1576_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w50_24_c10 :  std_logic;
signal bh1112_w51_20_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1576_Out0_copy1577_c10 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c0, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c1, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c2, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c3, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c4, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c5, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c6, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c7, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c8, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1578_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w51_21_c10 :  std_logic;
signal bh1112_w52_18_c10 :  std_logic;
signal bh1112_w53_14_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1578_Out0_copy1579_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1580_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1580_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w52_19_c10 :  std_logic;
signal bh1112_w53_15_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1580_Out0_copy1581_c10 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c0, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c1, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c2, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c3, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c4, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c5, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c6, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c7, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c8, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1582_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w53_16_c10 :  std_logic;
signal bh1112_w54_13_c10 :  std_logic;
signal bh1112_w55_11_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1582_Out0_copy1583_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1584_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1584_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w54_14_c10 :  std_logic;
signal bh1112_w55_12_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1584_Out0_copy1585_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1586_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1586_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1586_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w55_13_c10 :  std_logic;
signal bh1112_w56_10_c10 :  std_logic;
signal bh1112_w57_9_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1586_Out0_copy1587_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1588_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1588_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w57_10_c10 :  std_logic;
signal bh1112_w58_10_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1588_Out0_copy1589_c10 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1590_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1590_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w58_11_c10 :  std_logic;
signal bh1112_w59_6_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1590_Out0_copy1591_c10 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1592_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1592_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1592_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w60_8_c10 :  std_logic;
signal bh1112_w61_5_c10 :  std_logic;
signal bh1112_w62_7_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1592_Out0_copy1593_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1594_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1594_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1594_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w62_8_c10 :  std_logic;
signal bh1112_w63_5_c10 :  std_logic;
signal bh1112_w64_7_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1594_Out0_copy1595_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1596_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1596_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1596_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w64_8_c10 :  std_logic;
signal bh1112_w65_5_c10 :  std_logic;
signal bh1112_w66_7_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1596_Out0_copy1597_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1598_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1598_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1598_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w66_8_c10 :  std_logic;
signal bh1112_w67_5_c10 :  std_logic;
signal bh1112_w68_7_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1598_Out0_copy1599_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1600_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1600_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1600_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w68_8_c10 :  std_logic;
signal bh1112_w69_5_c10 :  std_logic;
signal bh1112_w70_6_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1600_Out0_copy1601_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1602_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1602_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1602_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w70_7_c10 :  std_logic;
signal bh1112_w71_4_c10 :  std_logic;
signal bh1112_w72_6_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1602_Out0_copy1603_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1604_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1604_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1604_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w72_7_c10 :  std_logic;
signal bh1112_w73_4_c10 :  std_logic;
signal bh1112_w74_6_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1604_Out0_copy1605_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1606_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1606_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1606_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w74_7_c10 :  std_logic;
signal bh1112_w75_4_c10 :  std_logic;
signal bh1112_w76_4_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1606_Out0_copy1607_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1608_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1608_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1608_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w76_5_c10 :  std_logic;
signal bh1112_w77_2_c10 :  std_logic;
signal bh1112_w78_2_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1608_Out0_copy1609_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1610_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1610_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1610_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1610_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w78_3_c10 :  std_logic;
signal bh1112_w79_1_c10 :  std_logic;
signal bh1112_w80_1_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1610_Out0_copy1611_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1612_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1612_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1612_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w40_32_c10 :  std_logic;
signal bh1112_w41_36_c10 :  std_logic;
signal bh1112_w42_40_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1612_Out0_copy1613_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1614_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1614_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w42_41_c10 :  std_logic;
signal bh1112_w43_41_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1614_Out0_copy1615_c10 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c0, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c1, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c2, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c3, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c4, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c5, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c6, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c7, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c8, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1616_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w43_42_c10 :  std_logic;
signal bh1112_w44_39_c10 :  std_logic;
signal bh1112_w45_37_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1616_Out0_copy1617_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1618_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1618_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w44_40_c10 :  std_logic;
signal bh1112_w45_38_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1618_Out0_copy1619_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1620_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1620_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1620_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w45_39_c10 :  std_logic;
signal bh1112_w46_35_c10 :  std_logic;
signal bh1112_w47_32_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1620_Out0_copy1621_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c0, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c1, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c2, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c3, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c4, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c5, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c6, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c7, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c8, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1622_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w47_33_c10 :  std_logic;
signal bh1112_w48_30_c10 :  std_logic;
signal bh1112_w49_28_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1622_Out0_copy1623_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1624_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1624_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w48_31_c10 :  std_logic;
signal bh1112_w49_29_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1624_Out0_copy1625_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1626_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1626_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1626_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w49_30_c10 :  std_logic;
signal bh1112_w50_25_c10 :  std_logic;
signal bh1112_w51_22_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1626_Out0_copy1627_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1628_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1628_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1628_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w51_23_c10 :  std_logic;
signal bh1112_w52_20_c10 :  std_logic;
signal bh1112_w53_17_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1628_Out0_copy1629_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1630_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1630_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1630_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w53_18_c10 :  std_logic;
signal bh1112_w54_15_c10 :  std_logic;
signal bh1112_w55_14_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1630_Out0_copy1631_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1632_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1632_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w55_15_c10 :  std_logic;
signal bh1112_w56_11_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1632_Out0_copy1633_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1634_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1634_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1634_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w57_11_c10 :  std_logic;
signal bh1112_w58_12_c10 :  std_logic;
signal bh1112_w59_7_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1634_Out0_copy1635_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1636_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1636_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1636_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w59_8_c10 :  std_logic;
signal bh1112_w60_9_c10 :  std_logic;
signal bh1112_w61_6_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1636_Out0_copy1637_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1638_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1638_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1638_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w62_9_c10 :  std_logic;
signal bh1112_w63_6_c10 :  std_logic;
signal bh1112_w64_9_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1638_Out0_copy1639_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1640_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1640_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1640_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w64_10_c10 :  std_logic;
signal bh1112_w65_6_c10 :  std_logic;
signal bh1112_w66_9_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1640_Out0_copy1641_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1642_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1642_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1642_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w66_10_c10 :  std_logic;
signal bh1112_w67_6_c10 :  std_logic;
signal bh1112_w68_9_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1642_Out0_copy1643_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1644_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1644_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1644_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w68_10_c10 :  std_logic;
signal bh1112_w69_6_c10 :  std_logic;
signal bh1112_w70_8_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1644_Out0_copy1645_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1646_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1646_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1646_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w70_9_c10 :  std_logic;
signal bh1112_w71_5_c10 :  std_logic;
signal bh1112_w72_8_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1646_Out0_copy1647_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1648_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1648_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1648_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w72_9_c10 :  std_logic;
signal bh1112_w73_5_c10 :  std_logic;
signal bh1112_w74_8_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1648_Out0_copy1649_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1650_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1650_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1650_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w74_9_c10 :  std_logic;
signal bh1112_w75_5_c10 :  std_logic;
signal bh1112_w76_6_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1650_Out0_copy1651_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1652_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1652_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1652_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w76_7_c10 :  std_logic;
signal bh1112_w77_3_c10 :  std_logic;
signal bh1112_w78_4_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1652_Out0_copy1653_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1654_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1654_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1654_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w78_5_c10 :  std_logic;
signal bh1112_w79_2_c10 :  std_logic;
signal bh1112_w80_2_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1654_Out0_copy1655_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1656_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1656_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1656_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1656_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w80_3_c10 :  std_logic;
signal bh1112_w81_1_c10 :  std_logic;
signal bh1112_w82_1_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1656_Out0_copy1657_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1658_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1658_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1658_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w42_42_c10 :  std_logic;
signal bh1112_w43_43_c10 :  std_logic;
signal bh1112_w44_41_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1658_Out0_copy1659_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1660_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1660_Out0_c10 :  std_logic_vector(1 downto 0);
signal bh1112_w44_42_c10 :  std_logic;
signal bh1112_w45_40_c10 :  std_logic;
signal Compressor_3_2_Freq300_uid1359_bh1112_uid1660_Out0_copy1661_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1662_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1662_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1662_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w45_41_c10 :  std_logic;
signal bh1112_w46_36_c10 :  std_logic;
signal bh1112_w47_34_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1662_Out0_copy1663_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1664_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1664_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1664_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w47_35_c10 :  std_logic;
signal bh1112_w48_32_c10 :  std_logic;
signal bh1112_w49_31_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1664_Out0_copy1665_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1666_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1666_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1666_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w49_32_c10 :  std_logic;
signal bh1112_w50_26_c10 :  std_logic;
signal bh1112_w51_24_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1666_Out0_copy1667_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1668_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1668_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1668_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w51_25_c10 :  std_logic;
signal bh1112_w52_21_c10 :  std_logic;
signal bh1112_w53_19_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1668_Out0_copy1669_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1670_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1670_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1670_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w53_20_c10 :  std_logic;
signal bh1112_w54_16_c10 :  std_logic;
signal bh1112_w55_16_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1670_Out0_copy1671_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1672_In0_c10 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1672_In1_c10 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1672_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w55_17_c10 :  std_logic;
signal bh1112_w56_12_c10 :  std_logic;
signal bh1112_w57_12_c10 :  std_logic;
signal Compressor_23_3_Freq300_uid1355_bh1112_uid1672_Out0_copy1673_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1674_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1674_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1674_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w59_9_c10 :  std_logic;
signal bh1112_w60_10_c10 :  std_logic;
signal bh1112_w61_7_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1674_Out0_copy1675_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1676_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1676_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1676_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w61_8_c10 :  std_logic;
signal bh1112_w62_10_c10 :  std_logic;
signal bh1112_w63_7_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1676_Out0_copy1677_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1678_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1678_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1678_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w64_11_c10 :  std_logic;
signal bh1112_w65_7_c10 :  std_logic;
signal bh1112_w66_11_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1678_Out0_copy1679_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1680_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1680_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1680_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w66_12_c10 :  std_logic;
signal bh1112_w67_7_c10 :  std_logic;
signal bh1112_w68_11_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1680_Out0_copy1681_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1682_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1682_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1682_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w68_12_c10 :  std_logic;
signal bh1112_w69_7_c10 :  std_logic;
signal bh1112_w70_10_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1682_Out0_copy1683_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1684_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1684_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1684_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w70_11_c10 :  std_logic;
signal bh1112_w71_6_c10 :  std_logic;
signal bh1112_w72_10_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1684_Out0_copy1685_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1686_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1686_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1686_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w72_11_c10 :  std_logic;
signal bh1112_w73_6_c10 :  std_logic;
signal bh1112_w74_10_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1686_Out0_copy1687_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1688_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1688_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1688_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w74_11_c10 :  std_logic;
signal bh1112_w75_6_c10 :  std_logic;
signal bh1112_w76_8_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1688_Out0_copy1689_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1690_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1690_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1690_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w76_9_c10 :  std_logic;
signal bh1112_w77_4_c10 :  std_logic;
signal bh1112_w78_6_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1690_Out0_copy1691_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1692_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1692_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1692_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w78_7_c10 :  std_logic;
signal bh1112_w79_3_c10 :  std_logic;
signal bh1112_w80_4_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1692_Out0_copy1693_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1694_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1694_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1694_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w80_5_c10 :  std_logic;
signal bh1112_w81_2_c10 :  std_logic;
signal bh1112_w82_2_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1694_Out0_copy1695_c10 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1696_In0_c10 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1696_In1_c9, Compressor_14_3_Freq300_uid1373_bh1112_uid1696_In1_c10 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1696_Out0_c10 :  std_logic_vector(2 downto 0);
signal bh1112_w82_3_c10 :  std_logic;
signal bh1112_w83_1_c10 :  std_logic;
signal bh1112_w84_1_c10 :  std_logic;
signal Compressor_14_3_Freq300_uid1373_bh1112_uid1696_Out0_copy1697_c10 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh1112_43_c10, tmp_bitheapResult_bh1112_43_c11 :  std_logic_vector(43 downto 0);
signal bitheapFinalAdd_bh1112_In0_c10 :  std_logic_vector(49 downto 0);
signal bitheapFinalAdd_bh1112_In1_c10 :  std_logic_vector(49 downto 0);
signal bitheapFinalAdd_bh1112_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh1112_Out_c11 :  std_logic_vector(49 downto 0);
signal bitheapResult_bh1112_c11 :  std_logic_vector(92 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               bh1112_w39_27_c6 <= bh1112_w39_27_c5;
               bh1112_w40_18_c6 <= bh1112_w40_18_c5;
               bh1112_w41_17_c6 <= bh1112_w41_17_c5;
               bh1112_w42_21_c6 <= bh1112_w42_21_c5;
               bh1112_w43_20_c6 <= bh1112_w43_20_c5;
               bh1112_w44_19_c6 <= bh1112_w44_19_c5;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c6 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c5;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c6 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c5;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c6 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c5;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c6 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c5;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c6 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c5;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c6 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c5;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c6 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c5;
            end if;
            if ce_7 = '1' then
               bh1112_w39_27_c7 <= bh1112_w39_27_c6;
               bh1112_w40_18_c7 <= bh1112_w40_18_c6;
               bh1112_w41_17_c7 <= bh1112_w41_17_c6;
               bh1112_w42_21_c7 <= bh1112_w42_21_c6;
               bh1112_w43_20_c7 <= bh1112_w43_20_c6;
               bh1112_w44_19_c7 <= bh1112_w44_19_c6;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c7 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c6;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c7 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c6;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c7 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c6;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c7 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c6;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c7 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c6;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c7 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c6;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c7 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c6;
            end if;
            if ce_8 = '1' then
               bh1112_w39_27_c8 <= bh1112_w39_27_c7;
               bh1112_w40_18_c8 <= bh1112_w40_18_c7;
               bh1112_w41_17_c8 <= bh1112_w41_17_c7;
               bh1112_w42_21_c8 <= bh1112_w42_21_c7;
               bh1112_w43_20_c8 <= bh1112_w43_20_c7;
               bh1112_w44_19_c8 <= bh1112_w44_19_c7;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c8 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c7;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c8 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c7;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c8 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c7;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c8 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c7;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c8 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c7;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c8 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c7;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c8 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c7;
            end if;
            if ce_9 = '1' then
               bh1112_w39_27_c9 <= bh1112_w39_27_c8;
               bh1112_w40_18_c9 <= bh1112_w40_18_c8;
               bh1112_w41_17_c9 <= bh1112_w41_17_c8;
               bh1112_w42_21_c9 <= bh1112_w42_21_c8;
               bh1112_w43_20_c9 <= bh1112_w43_20_c8;
               bh1112_w44_19_c9 <= bh1112_w44_19_c8;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c8;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c8;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c8;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c8;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c8;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c8;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c8;
            end if;
            if ce_10 = '1' then
               bh1112_w29_0_c10 <= bh1112_w29_0_c9;
               bh1112_w30_0_c10 <= bh1112_w30_0_c9;
               bh1112_w31_0_c10 <= bh1112_w31_0_c9;
               bh1112_w32_0_c10 <= bh1112_w32_0_c9;
               bh1112_w33_0_c10 <= bh1112_w33_0_c9;
               bh1112_w34_0_c10 <= bh1112_w34_0_c9;
               bh1112_w35_0_c10 <= bh1112_w35_0_c9;
               bh1112_w76_0_c10 <= bh1112_w76_0_c9;
               bh1112_w78_0_c10 <= bh1112_w78_0_c9;
               bh1112_w80_0_c10 <= bh1112_w80_0_c9;
               bh1112_w82_0_c10 <= bh1112_w82_0_c9;
               bh1112_w84_0_c10 <= bh1112_w84_0_c9;
               bh1112_w85_0_c10 <= bh1112_w85_0_c9;
               bh1112_w86_0_c10 <= bh1112_w86_0_c9;
               bh1112_w87_0_c10 <= bh1112_w87_0_c9;
               bh1112_w88_0_c10 <= bh1112_w88_0_c9;
               bh1112_w89_0_c10 <= bh1112_w89_0_c9;
               bh1112_w90_0_c10 <= bh1112_w90_0_c9;
               bh1112_w91_0_c10 <= bh1112_w91_0_c9;
               bh1112_w92_0_c10 <= bh1112_w92_0_c9;
               bh1112_w61_2_c10 <= bh1112_w61_2_c9;
               bh1112_w63_2_c10 <= bh1112_w63_2_c9;
               bh1112_w65_2_c10 <= bh1112_w65_2_c9;
               bh1112_w67_2_c10 <= bh1112_w67_2_c9;
               bh1112_w69_2_c10 <= bh1112_w69_2_c9;
               bh1112_w49_6_c10 <= bh1112_w49_6_c9;
               bh1112_w48_9_c10 <= bh1112_w48_9_c9;
               bh1112_w53_6_c10 <= bh1112_w53_6_c9;
               bh1112_w56_4_c10 <= bh1112_w56_4_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_copy1357_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_copy1357_c9;
               Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_copy1361_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_copy1361_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_copy1365_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_copy1365_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_copy1367_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_copy1367_c9;
               bh1112_w39_31_c10 <= bh1112_w39_31_c9;
               bh1112_w40_21_c10 <= bh1112_w40_21_c9;
               bh1112_w41_20_c10 <= bh1112_w41_20_c9;
               bh1112_w39_32_c10 <= bh1112_w39_32_c9;
               bh1112_w40_22_c10 <= bh1112_w40_22_c9;
               bh1112_w41_21_c10 <= bh1112_w41_21_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_copy1375_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_copy1375_c9;
               bh1112_w40_24_c10 <= bh1112_w40_24_c9;
               bh1112_w41_23_c10 <= bh1112_w41_23_c9;
               bh1112_w42_22_c10 <= bh1112_w42_22_c9;
               bh1112_w40_25_c10 <= bh1112_w40_25_c9;
               bh1112_w41_24_c10 <= bh1112_w41_24_c9;
               bh1112_w42_23_c10 <= bh1112_w42_23_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_copy1381_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_copy1381_c9;
               bh1112_w41_26_c10 <= bh1112_w41_26_c9;
               bh1112_w42_25_c10 <= bh1112_w42_25_c9;
               bh1112_w43_21_c10 <= bh1112_w43_21_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_copy1385_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_copy1385_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_copy1387_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_copy1387_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_copy1389_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_copy1389_c9;
               bh1112_w42_29_c10 <= bh1112_w42_29_c9;
               bh1112_w43_25_c10 <= bh1112_w43_25_c9;
               bh1112_w44_21_c10 <= bh1112_w44_21_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_copy1393_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_copy1393_c9;
               bh1112_w42_31_c10 <= bh1112_w42_31_c9;
               bh1112_w43_27_c10 <= bh1112_w43_27_c9;
               bh1112_w43_28_c10 <= bh1112_w43_28_c9;
               bh1112_w44_24_c10 <= bh1112_w44_24_c9;
               bh1112_w45_18_c10 <= bh1112_w45_18_c9;
               bh1112_w43_29_c10 <= bh1112_w43_29_c9;
               bh1112_w45_19_c10 <= bh1112_w45_19_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_copy1401_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_copy1401_c9;
               bh1112_w43_31_c10 <= bh1112_w43_31_c9;
               bh1112_w45_21_c10 <= bh1112_w45_21_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_copy1405_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_copy1405_c9;
               bh1112_w45_23_c10 <= bh1112_w45_23_c9;
               bh1112_w46_19_c10 <= bh1112_w46_19_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_copy1409_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_copy1409_c9;
               bh1112_w45_25_c10 <= bh1112_w45_25_c9;
               bh1112_w46_21_c10 <= bh1112_w46_21_c9;
               bh1112_w47_15_c10 <= bh1112_w47_15_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_copy1413_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_copy1413_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_copy1415_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_copy1415_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_copy1417_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_copy1417_c9;
               bh1112_w46_25_c10 <= bh1112_w46_25_c9;
               bh1112_w47_19_c10 <= bh1112_w47_19_c9;
               bh1112_w48_16_c10 <= bh1112_w48_16_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_copy1421_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_copy1421_c9;
               bh1112_w47_21_c10 <= bh1112_w47_21_c9;
               bh1112_w48_18_c10 <= bh1112_w48_18_c9;
               bh1112_w49_13_c10 <= bh1112_w49_13_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_copy1425_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_copy1425_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_copy1427_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_copy1427_c9;
               bh1112_w48_21_c10 <= bh1112_w48_21_c9;
               bh1112_w49_16_c10 <= bh1112_w49_16_c9;
               bh1112_w50_11_c10 <= bh1112_w50_11_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_copy1431_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_copy1431_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_copy1433_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_copy1433_c9;
               bh1112_w49_19_c10 <= bh1112_w49_19_c9;
               bh1112_w50_14_c10 <= bh1112_w50_14_c9;
               bh1112_w51_10_c10 <= bh1112_w51_10_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_copy1437_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_copy1437_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_copy1439_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_copy1439_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_copy1441_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_copy1441_c9;
               bh1112_w51_14_c10 <= bh1112_w51_14_c9;
               bh1112_w52_12_c10 <= bh1112_w52_12_c9;
               bh1112_w53_7_c10 <= bh1112_w53_7_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_copy1445_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_copy1445_c9;
               bh1112_w52_14_c10 <= bh1112_w52_14_c9;
               bh1112_w53_9_c10 <= bh1112_w53_9_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_copy1449_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_copy1449_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_copy1451_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_copy1451_c9;
               Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_copy1453_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_copy1453_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_copy1455_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_copy1455_c9;
               Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_copy1457_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_copy1457_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_copy1459_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_copy1459_c9;
               Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_copy1461_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_copy1461_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_copy1463_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_copy1463_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_copy1465_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_copy1465_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_copy1467_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_copy1467_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_copy1469_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_copy1469_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_copy1471_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_copy1471_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_copy1473_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_copy1473_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_copy1475_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_copy1475_c9;
               Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_copy1477_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_copy1477_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1500_In0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1500_In0_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1524_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1524_In1_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1550_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1550_In1_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1610_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1610_In1_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1656_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1656_In1_c9;
               Compressor_14_3_Freq300_uid1373_bh1112_uid1696_In1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1696_In1_c9;
            end if;
            if ce_11 = '1' then
               tmp_bitheapResult_bh1112_43_c11 <= tmp_bitheapResult_bh1112_43_c10;
            end if;
         end if;
      end process;
   XX_m1111_c5 <= X ;
   YY_m1111_c9 <= Y ;
   tile_0_X_c5 <= X(45 downto 29);
   tile_0_Y_c9 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid1114
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_0_X_c5,
                 Y => tile_0_Y_c9,
                 R => tile_0_output_c9);

   tile_0_filtered_output_c9 <= unsigned(tile_0_output_c9(40 downto 0));
   bh1112_w29_0_c9 <= tile_0_filtered_output_c9(0);
   bh1112_w30_0_c9 <= tile_0_filtered_output_c9(1);
   bh1112_w31_0_c9 <= tile_0_filtered_output_c9(2);
   bh1112_w32_0_c9 <= tile_0_filtered_output_c9(3);
   bh1112_w33_0_c9 <= tile_0_filtered_output_c9(4);
   bh1112_w34_0_c9 <= tile_0_filtered_output_c9(5);
   bh1112_w35_0_c9 <= tile_0_filtered_output_c9(6);
   bh1112_w36_0_c9 <= tile_0_filtered_output_c9(7);
   bh1112_w37_0_c9 <= tile_0_filtered_output_c9(8);
   bh1112_w38_0_c9 <= tile_0_filtered_output_c9(9);
   bh1112_w39_0_c9 <= tile_0_filtered_output_c9(10);
   bh1112_w40_0_c9 <= tile_0_filtered_output_c9(11);
   bh1112_w41_0_c9 <= tile_0_filtered_output_c9(12);
   bh1112_w42_0_c9 <= tile_0_filtered_output_c9(13);
   bh1112_w43_0_c9 <= tile_0_filtered_output_c9(14);
   bh1112_w44_0_c9 <= tile_0_filtered_output_c9(15);
   bh1112_w45_0_c9 <= tile_0_filtered_output_c9(16);
   bh1112_w46_0_c9 <= tile_0_filtered_output_c9(17);
   bh1112_w47_0_c9 <= tile_0_filtered_output_c9(18);
   bh1112_w48_0_c9 <= tile_0_filtered_output_c9(19);
   bh1112_w49_0_c9 <= tile_0_filtered_output_c9(20);
   bh1112_w50_0_c9 <= tile_0_filtered_output_c9(21);
   bh1112_w51_0_c9 <= tile_0_filtered_output_c9(22);
   bh1112_w52_0_c9 <= tile_0_filtered_output_c9(23);
   bh1112_w53_0_c9 <= tile_0_filtered_output_c9(24);
   bh1112_w54_0_c9 <= tile_0_filtered_output_c9(25);
   bh1112_w55_0_c9 <= tile_0_filtered_output_c9(26);
   bh1112_w56_0_c9 <= tile_0_filtered_output_c9(27);
   bh1112_w57_0_c9 <= tile_0_filtered_output_c9(28);
   bh1112_w58_0_c9 <= tile_0_filtered_output_c9(29);
   bh1112_w59_0_c9 <= tile_0_filtered_output_c9(30);
   bh1112_w60_0_c9 <= tile_0_filtered_output_c9(31);
   bh1112_w61_0_c9 <= tile_0_filtered_output_c9(32);
   bh1112_w62_0_c9 <= tile_0_filtered_output_c9(33);
   bh1112_w63_0_c9 <= tile_0_filtered_output_c9(34);
   bh1112_w64_0_c9 <= tile_0_filtered_output_c9(35);
   bh1112_w65_0_c9 <= tile_0_filtered_output_c9(36);
   bh1112_w66_0_c9 <= tile_0_filtered_output_c9(37);
   bh1112_w67_0_c9 <= tile_0_filtered_output_c9(38);
   bh1112_w68_0_c9 <= tile_0_filtered_output_c9(39);
   bh1112_w69_0_c9 <= tile_0_filtered_output_c9(40);
   tile_1_X_c5 <= X(28 downto 28);
   tile_1_Y_c9 <= Y(11 downto 11);
   tile_1_mult: IntMultiplierLUT_1x1_Freq300_uid1116
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_1_X_c5,
                 Y => tile_1_Y_c9,
                 R => tile_1_output_c9);

   tile_1_filtered_output_c9 <= unsigned(tile_1_output_c9(0 downto 0));
   bh1112_w39_1_c9 <= tile_1_filtered_output_c9(0);
   tile_2_X_c5 <= X(26 downto 26);
   tile_2_Y_c9 <= Y(13 downto 13);
   tile_2_mult: IntMultiplierLUT_1x1_Freq300_uid1118
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_2_X_c5,
                 Y => tile_2_Y_c9,
                 R => tile_2_output_c9);

   tile_2_filtered_output_c9 <= unsigned(tile_2_output_c9(0 downto 0));
   bh1112_w39_2_c9 <= tile_2_filtered_output_c9(0);
   tile_3_X_c5 <= X(28 downto 27);
   tile_3_Y_c9 <= Y(13 downto 12);
   tile_3_mult: IntMultiplierLUT_2x2_Freq300_uid1120
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_3_X_c5,
                 Y => tile_3_Y_c9,
                 R => tile_3_output_c9);

   tile_3_filtered_output_c9 <= unsigned(tile_3_output_c9(3 downto 0));
   bh1112_w39_3_c9 <= tile_3_filtered_output_c9(0);
   bh1112_w40_1_c9 <= tile_3_filtered_output_c9(1);
   bh1112_w41_1_c9 <= tile_3_filtered_output_c9(2);
   bh1112_w42_1_c9 <= tile_3_filtered_output_c9(3);
   tile_4_X_c5 <= X(25 downto 25);
   tile_4_Y_c9 <= Y(14 downto 14);
   tile_4_mult: IntMultiplierLUT_1x1_Freq300_uid1125
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_4_X_c5,
                 Y => tile_4_Y_c9,
                 R => tile_4_output_c9);

   tile_4_filtered_output_c9 <= unsigned(tile_4_output_c9(0 downto 0));
   bh1112_w39_4_c9 <= tile_4_filtered_output_c9(0);
   tile_5_X_c5 <= X(25 downto 24);
   tile_5_Y_c9 <= Y(15 downto 15);
   tile_5_mult: IntMultiplierLUT_2x1_Freq300_uid1127
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_5_X_c5,
                 Y => tile_5_Y_c9,
                 R => tile_5_output_c9);

   tile_5_filtered_output_c9 <= unsigned(tile_5_output_c9(1 downto 0));
   bh1112_w39_5_c9 <= tile_5_filtered_output_c9(0);
   bh1112_w40_2_c9 <= tile_5_filtered_output_c9(1);
   tile_6_X_c5 <= X(28 downto 26);
   tile_6_Y_c9 <= Y(15 downto 14);
   tile_6_mult: IntMultiplierLUT_3x2_Freq300_uid1129
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_6_X_c5,
                 Y => tile_6_Y_c9,
                 R => tile_6_output_c9);

   tile_6_filtered_output_c9 <= unsigned(tile_6_output_c9(4 downto 0));
   bh1112_w40_3_c9 <= tile_6_filtered_output_c9(0);
   bh1112_w41_2_c9 <= tile_6_filtered_output_c9(1);
   bh1112_w42_2_c9 <= tile_6_filtered_output_c9(2);
   bh1112_w43_1_c9 <= tile_6_filtered_output_c9(3);
   bh1112_w44_1_c9 <= tile_6_filtered_output_c9(4);
   tile_7_X_c5 <= X(22 downto 22);
   tile_7_Y_c9 <= Y(17 downto 17);
   tile_7_mult: IntMultiplierLUT_1x1_Freq300_uid1134
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_7_X_c5,
                 Y => tile_7_Y_c9,
                 R => tile_7_output_c9);

   tile_7_filtered_output_c9 <= unsigned(tile_7_output_c9(0 downto 0));
   bh1112_w39_6_c9 <= tile_7_filtered_output_c9(0);
   tile_8_X_c5 <= X(25 downto 23);
   tile_8_Y_c9 <= Y(17 downto 16);
   tile_8_mult: IntMultiplierLUT_3x2_Freq300_uid1136
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_8_X_c5,
                 Y => tile_8_Y_c9,
                 R => tile_8_output_c9);

   tile_8_filtered_output_c9 <= unsigned(tile_8_output_c9(4 downto 0));
   bh1112_w39_7_c9 <= tile_8_filtered_output_c9(0);
   bh1112_w40_4_c9 <= tile_8_filtered_output_c9(1);
   bh1112_w41_3_c9 <= tile_8_filtered_output_c9(2);
   bh1112_w42_3_c9 <= tile_8_filtered_output_c9(3);
   bh1112_w43_2_c9 <= tile_8_filtered_output_c9(4);
   tile_9_X_c5 <= X(28 downto 26);
   tile_9_Y_c9 <= Y(17 downto 16);
   tile_9_mult: IntMultiplierLUT_3x2_Freq300_uid1141
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_9_X_c5,
                 Y => tile_9_Y_c9,
                 R => tile_9_output_c9);

   tile_9_filtered_output_c9 <= unsigned(tile_9_output_c9(4 downto 0));
   bh1112_w42_4_c9 <= tile_9_filtered_output_c9(0);
   bh1112_w43_3_c9 <= tile_9_filtered_output_c9(1);
   bh1112_w44_2_c9 <= tile_9_filtered_output_c9(2);
   bh1112_w45_1_c9 <= tile_9_filtered_output_c9(3);
   bh1112_w46_1_c9 <= tile_9_filtered_output_c9(4);
   tile_10_X_c5 <= X(20 downto 20);
   tile_10_Y_c9 <= Y(19 downto 19);
   tile_10_mult: IntMultiplierLUT_1x1_Freq300_uid1146
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_10_X_c5,
                 Y => tile_10_Y_c9,
                 R => tile_10_output_c9);

   tile_10_filtered_output_c9 <= unsigned(tile_10_output_c9(0 downto 0));
   bh1112_w39_8_c9 <= tile_10_filtered_output_c9(0);
   tile_11_X_c5 <= X(22 downto 21);
   tile_11_Y_c9 <= Y(19 downto 18);
   tile_11_mult: IntMultiplierLUT_2x2_Freq300_uid1148
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_11_X_c5,
                 Y => tile_11_Y_c9,
                 R => tile_11_output_c9);

   tile_11_filtered_output_c9 <= unsigned(tile_11_output_c9(3 downto 0));
   bh1112_w39_9_c9 <= tile_11_filtered_output_c9(0);
   bh1112_w40_5_c9 <= tile_11_filtered_output_c9(1);
   bh1112_w41_4_c9 <= tile_11_filtered_output_c9(2);
   bh1112_w42_5_c9 <= tile_11_filtered_output_c9(3);
   tile_12_X_c5 <= X(25 downto 23);
   tile_12_Y_c9 <= Y(19 downto 18);
   tile_12_mult: IntMultiplierLUT_3x2_Freq300_uid1153
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_12_X_c5,
                 Y => tile_12_Y_c9,
                 R => tile_12_output_c9);

   tile_12_filtered_output_c9 <= unsigned(tile_12_output_c9(4 downto 0));
   bh1112_w41_5_c9 <= tile_12_filtered_output_c9(0);
   bh1112_w42_6_c9 <= tile_12_filtered_output_c9(1);
   bh1112_w43_4_c9 <= tile_12_filtered_output_c9(2);
   bh1112_w44_3_c9 <= tile_12_filtered_output_c9(3);
   bh1112_w45_2_c9 <= tile_12_filtered_output_c9(4);
   tile_13_X_c5 <= X(28 downto 26);
   tile_13_Y_c9 <= Y(19 downto 18);
   tile_13_mult: IntMultiplierLUT_3x2_Freq300_uid1158
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_13_X_c5,
                 Y => tile_13_Y_c9,
                 R => tile_13_output_c9);

   tile_13_filtered_output_c9 <= unsigned(tile_13_output_c9(4 downto 0));
   bh1112_w44_4_c9 <= tile_13_filtered_output_c9(0);
   bh1112_w45_3_c9 <= tile_13_filtered_output_c9(1);
   bh1112_w46_2_c9 <= tile_13_filtered_output_c9(2);
   bh1112_w47_1_c9 <= tile_13_filtered_output_c9(3);
   bh1112_w48_1_c9 <= tile_13_filtered_output_c9(4);
   tile_14_X_c5 <= X(19 downto 19);
   tile_14_Y_c9 <= Y(20 downto 20);
   tile_14_mult: IntMultiplierLUT_1x1_Freq300_uid1163
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_14_X_c5,
                 Y => tile_14_Y_c9,
                 R => tile_14_output_c9);

   tile_14_filtered_output_c9 <= unsigned(tile_14_output_c9(0 downto 0));
   bh1112_w39_10_c9 <= tile_14_filtered_output_c9(0);
   tile_15_X_c5 <= X(19 downto 18);
   tile_15_Y_c9 <= Y(21 downto 21);
   tile_15_mult: IntMultiplierLUT_2x1_Freq300_uid1165
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_15_X_c5,
                 Y => tile_15_Y_c9,
                 R => tile_15_output_c9);

   tile_15_filtered_output_c9 <= unsigned(tile_15_output_c9(1 downto 0));
   bh1112_w39_11_c9 <= tile_15_filtered_output_c9(0);
   bh1112_w40_6_c9 <= tile_15_filtered_output_c9(1);
   tile_16_X_c5 <= X(22 downto 20);
   tile_16_Y_c9 <= Y(21 downto 20);
   tile_16_mult: IntMultiplierLUT_3x2_Freq300_uid1167
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_16_X_c5,
                 Y => tile_16_Y_c9,
                 R => tile_16_output_c9);

   tile_16_filtered_output_c9 <= unsigned(tile_16_output_c9(4 downto 0));
   bh1112_w40_7_c9 <= tile_16_filtered_output_c9(0);
   bh1112_w41_6_c9 <= tile_16_filtered_output_c9(1);
   bh1112_w42_7_c9 <= tile_16_filtered_output_c9(2);
   bh1112_w43_5_c9 <= tile_16_filtered_output_c9(3);
   bh1112_w44_5_c9 <= tile_16_filtered_output_c9(4);
   tile_17_X_c5 <= X(25 downto 23);
   tile_17_Y_c9 <= Y(21 downto 20);
   tile_17_mult: IntMultiplierLUT_3x2_Freq300_uid1172
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_17_X_c5,
                 Y => tile_17_Y_c9,
                 R => tile_17_output_c9);

   tile_17_filtered_output_c9 <= unsigned(tile_17_output_c9(4 downto 0));
   bh1112_w43_6_c9 <= tile_17_filtered_output_c9(0);
   bh1112_w44_6_c9 <= tile_17_filtered_output_c9(1);
   bh1112_w45_4_c9 <= tile_17_filtered_output_c9(2);
   bh1112_w46_3_c9 <= tile_17_filtered_output_c9(3);
   bh1112_w47_2_c9 <= tile_17_filtered_output_c9(4);
   tile_18_X_c5 <= X(28 downto 26);
   tile_18_Y_c9 <= Y(21 downto 20);
   tile_18_mult: IntMultiplierLUT_3x2_Freq300_uid1177
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_18_X_c5,
                 Y => tile_18_Y_c9,
                 R => tile_18_output_c9);

   tile_18_filtered_output_c9 <= unsigned(tile_18_output_c9(4 downto 0));
   bh1112_w46_4_c9 <= tile_18_filtered_output_c9(0);
   bh1112_w47_3_c9 <= tile_18_filtered_output_c9(1);
   bh1112_w48_2_c9 <= tile_18_filtered_output_c9(2);
   bh1112_w49_1_c9 <= tile_18_filtered_output_c9(3);
   bh1112_w50_1_c9 <= tile_18_filtered_output_c9(4);
   tile_19_X_c5 <= X(16 downto 16);
   tile_19_Y_c9 <= Y(23 downto 23);
   tile_19_mult: IntMultiplierLUT_1x1_Freq300_uid1182
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_19_X_c5,
                 Y => tile_19_Y_c9,
                 R => tile_19_output_c9);

   tile_19_filtered_output_c9 <= unsigned(tile_19_output_c9(0 downto 0));
   bh1112_w39_12_c9 <= tile_19_filtered_output_c9(0);
   tile_20_X_c5 <= X(19 downto 17);
   tile_20_Y_c9 <= Y(23 downto 22);
   tile_20_mult: IntMultiplierLUT_3x2_Freq300_uid1184
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_20_X_c5,
                 Y => tile_20_Y_c9,
                 R => tile_20_output_c9);

   tile_20_filtered_output_c9 <= unsigned(tile_20_output_c9(4 downto 0));
   bh1112_w39_13_c9 <= tile_20_filtered_output_c9(0);
   bh1112_w40_8_c9 <= tile_20_filtered_output_c9(1);
   bh1112_w41_7_c9 <= tile_20_filtered_output_c9(2);
   bh1112_w42_8_c9 <= tile_20_filtered_output_c9(3);
   bh1112_w43_7_c9 <= tile_20_filtered_output_c9(4);
   tile_21_X_c5 <= X(22 downto 20);
   tile_21_Y_c9 <= Y(23 downto 22);
   tile_21_mult: IntMultiplierLUT_3x2_Freq300_uid1189
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_21_X_c5,
                 Y => tile_21_Y_c9,
                 R => tile_21_output_c9);

   tile_21_filtered_output_c9 <= unsigned(tile_21_output_c9(4 downto 0));
   bh1112_w42_9_c9 <= tile_21_filtered_output_c9(0);
   bh1112_w43_8_c9 <= tile_21_filtered_output_c9(1);
   bh1112_w44_7_c9 <= tile_21_filtered_output_c9(2);
   bh1112_w45_5_c9 <= tile_21_filtered_output_c9(3);
   bh1112_w46_5_c9 <= tile_21_filtered_output_c9(4);
   tile_22_X_c5 <= X(25 downto 23);
   tile_22_Y_c9 <= Y(23 downto 22);
   tile_22_mult: IntMultiplierLUT_3x2_Freq300_uid1194
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_22_X_c5,
                 Y => tile_22_Y_c9,
                 R => tile_22_output_c9);

   tile_22_filtered_output_c9 <= unsigned(tile_22_output_c9(4 downto 0));
   bh1112_w45_6_c9 <= tile_22_filtered_output_c9(0);
   bh1112_w46_6_c9 <= tile_22_filtered_output_c9(1);
   bh1112_w47_4_c9 <= tile_22_filtered_output_c9(2);
   bh1112_w48_3_c9 <= tile_22_filtered_output_c9(3);
   bh1112_w49_2_c9 <= tile_22_filtered_output_c9(4);
   tile_23_X_c5 <= X(28 downto 26);
   tile_23_Y_c9 <= Y(23 downto 22);
   tile_23_mult: IntMultiplierLUT_3x2_Freq300_uid1199
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_23_X_c5,
                 Y => tile_23_Y_c9,
                 R => tile_23_output_c9);

   tile_23_filtered_output_c9 <= unsigned(tile_23_output_c9(4 downto 0));
   bh1112_w48_4_c9 <= tile_23_filtered_output_c9(0);
   bh1112_w49_3_c9 <= tile_23_filtered_output_c9(1);
   bh1112_w50_2_c9 <= tile_23_filtered_output_c9(2);
   bh1112_w51_1_c9 <= tile_23_filtered_output_c9(3);
   bh1112_w52_1_c9 <= tile_23_filtered_output_c9(4);
   tile_24_X_c5 <= X(45 downto 29);
   tile_24_Y_c9 <= Y(46 downto 24);
   tile_24_mult: DSPBlock_17x23_Freq300_uid1204
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_24_X_c5,
                 Y => tile_24_Y_c9,
                 R => tile_24_output_c9);

   tile_24_filtered_output_c9 <= unsigned(tile_24_output_c9(39 downto 0));
   bh1112_w53_1_c9 <= tile_24_filtered_output_c9(0);
   bh1112_w54_1_c9 <= tile_24_filtered_output_c9(1);
   bh1112_w55_1_c9 <= tile_24_filtered_output_c9(2);
   bh1112_w56_1_c9 <= tile_24_filtered_output_c9(3);
   bh1112_w57_1_c9 <= tile_24_filtered_output_c9(4);
   bh1112_w58_1_c9 <= tile_24_filtered_output_c9(5);
   bh1112_w59_1_c9 <= tile_24_filtered_output_c9(6);
   bh1112_w60_1_c9 <= tile_24_filtered_output_c9(7);
   bh1112_w61_1_c9 <= tile_24_filtered_output_c9(8);
   bh1112_w62_1_c9 <= tile_24_filtered_output_c9(9);
   bh1112_w63_1_c9 <= tile_24_filtered_output_c9(10);
   bh1112_w64_1_c9 <= tile_24_filtered_output_c9(11);
   bh1112_w65_1_c9 <= tile_24_filtered_output_c9(12);
   bh1112_w66_1_c9 <= tile_24_filtered_output_c9(13);
   bh1112_w67_1_c9 <= tile_24_filtered_output_c9(14);
   bh1112_w68_1_c9 <= tile_24_filtered_output_c9(15);
   bh1112_w69_1_c9 <= tile_24_filtered_output_c9(16);
   bh1112_w70_0_c9 <= tile_24_filtered_output_c9(17);
   bh1112_w71_0_c9 <= tile_24_filtered_output_c9(18);
   bh1112_w72_0_c9 <= tile_24_filtered_output_c9(19);
   bh1112_w73_0_c9 <= tile_24_filtered_output_c9(20);
   bh1112_w74_0_c9 <= tile_24_filtered_output_c9(21);
   bh1112_w75_0_c9 <= tile_24_filtered_output_c9(22);
   bh1112_w76_0_c9 <= tile_24_filtered_output_c9(23);
   bh1112_w77_0_c9 <= tile_24_filtered_output_c9(24);
   bh1112_w78_0_c9 <= tile_24_filtered_output_c9(25);
   bh1112_w79_0_c9 <= tile_24_filtered_output_c9(26);
   bh1112_w80_0_c9 <= tile_24_filtered_output_c9(27);
   bh1112_w81_0_c9 <= tile_24_filtered_output_c9(28);
   bh1112_w82_0_c9 <= tile_24_filtered_output_c9(29);
   bh1112_w83_0_c9 <= tile_24_filtered_output_c9(30);
   bh1112_w84_0_c9 <= tile_24_filtered_output_c9(31);
   bh1112_w85_0_c9 <= tile_24_filtered_output_c9(32);
   bh1112_w86_0_c9 <= tile_24_filtered_output_c9(33);
   bh1112_w87_0_c9 <= tile_24_filtered_output_c9(34);
   bh1112_w88_0_c9 <= tile_24_filtered_output_c9(35);
   bh1112_w89_0_c9 <= tile_24_filtered_output_c9(36);
   bh1112_w90_0_c9 <= tile_24_filtered_output_c9(37);
   bh1112_w91_0_c9 <= tile_24_filtered_output_c9(38);
   bh1112_w92_0_c9 <= tile_24_filtered_output_c9(39);
   tile_25_X_c5 <= X(28 downto 12);
   tile_25_Y_c9 <= Y(46 downto 24);
   tile_25_mult: DSPBlock_17x23_Freq300_uid1206
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_25_X_c5,
                 Y => tile_25_Y_c9,
                 R => tile_25_output_c9);

   tile_25_filtered_output_c9 <= unsigned(tile_25_output_c9(39 downto 0));
   bh1112_w36_1_c9 <= tile_25_filtered_output_c9(0);
   bh1112_w37_1_c9 <= tile_25_filtered_output_c9(1);
   bh1112_w38_1_c9 <= tile_25_filtered_output_c9(2);
   bh1112_w39_14_c9 <= tile_25_filtered_output_c9(3);
   bh1112_w40_9_c9 <= tile_25_filtered_output_c9(4);
   bh1112_w41_8_c9 <= tile_25_filtered_output_c9(5);
   bh1112_w42_10_c9 <= tile_25_filtered_output_c9(6);
   bh1112_w43_9_c9 <= tile_25_filtered_output_c9(7);
   bh1112_w44_8_c9 <= tile_25_filtered_output_c9(8);
   bh1112_w45_7_c9 <= tile_25_filtered_output_c9(9);
   bh1112_w46_7_c9 <= tile_25_filtered_output_c9(10);
   bh1112_w47_5_c9 <= tile_25_filtered_output_c9(11);
   bh1112_w48_5_c9 <= tile_25_filtered_output_c9(12);
   bh1112_w49_4_c9 <= tile_25_filtered_output_c9(13);
   bh1112_w50_3_c9 <= tile_25_filtered_output_c9(14);
   bh1112_w51_2_c9 <= tile_25_filtered_output_c9(15);
   bh1112_w52_2_c9 <= tile_25_filtered_output_c9(16);
   bh1112_w53_2_c9 <= tile_25_filtered_output_c9(17);
   bh1112_w54_2_c9 <= tile_25_filtered_output_c9(18);
   bh1112_w55_2_c9 <= tile_25_filtered_output_c9(19);
   bh1112_w56_2_c9 <= tile_25_filtered_output_c9(20);
   bh1112_w57_2_c9 <= tile_25_filtered_output_c9(21);
   bh1112_w58_2_c9 <= tile_25_filtered_output_c9(22);
   bh1112_w59_2_c9 <= tile_25_filtered_output_c9(23);
   bh1112_w60_2_c9 <= tile_25_filtered_output_c9(24);
   bh1112_w61_2_c9 <= tile_25_filtered_output_c9(25);
   bh1112_w62_2_c9 <= tile_25_filtered_output_c9(26);
   bh1112_w63_2_c9 <= tile_25_filtered_output_c9(27);
   bh1112_w64_2_c9 <= tile_25_filtered_output_c9(28);
   bh1112_w65_2_c9 <= tile_25_filtered_output_c9(29);
   bh1112_w66_2_c9 <= tile_25_filtered_output_c9(30);
   bh1112_w67_2_c9 <= tile_25_filtered_output_c9(31);
   bh1112_w68_2_c9 <= tile_25_filtered_output_c9(32);
   bh1112_w69_2_c9 <= tile_25_filtered_output_c9(33);
   bh1112_w70_1_c9 <= tile_25_filtered_output_c9(34);
   bh1112_w71_1_c9 <= tile_25_filtered_output_c9(35);
   bh1112_w72_1_c9 <= tile_25_filtered_output_c9(36);
   bh1112_w73_1_c9 <= tile_25_filtered_output_c9(37);
   bh1112_w74_1_c9 <= tile_25_filtered_output_c9(38);
   bh1112_w75_1_c9 <= tile_25_filtered_output_c9(39);
   tile_26_X_c5 <= X(11 downto 11);
   tile_26_Y_c9 <= Y(28 downto 28);
   tile_26_mult: IntMultiplierLUT_1x1_Freq300_uid1208
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_26_X_c5,
                 Y => tile_26_Y_c9,
                 R => tile_26_output_c9);

   tile_26_filtered_output_c9 <= unsigned(tile_26_output_c9(0 downto 0));
   bh1112_w39_15_c9 <= tile_26_filtered_output_c9(0);
   tile_27_X_c5 <= X(9 downto 9);
   tile_27_Y_c9 <= Y(30 downto 30);
   tile_27_mult: IntMultiplierLUT_1x1_Freq300_uid1210
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_27_X_c5,
                 Y => tile_27_Y_c9,
                 R => tile_27_output_c9);

   tile_27_filtered_output_c9 <= unsigned(tile_27_output_c9(0 downto 0));
   bh1112_w39_16_c9 <= tile_27_filtered_output_c9(0);
   tile_28_X_c5 <= X(11 downto 10);
   tile_28_Y_c9 <= Y(30 downto 29);
   tile_28_mult: IntMultiplierLUT_2x2_Freq300_uid1212
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_28_X_c5,
                 Y => tile_28_Y_c9,
                 R => tile_28_output_c9);

   tile_28_filtered_output_c9 <= unsigned(tile_28_output_c9(3 downto 0));
   bh1112_w39_17_c9 <= tile_28_filtered_output_c9(0);
   bh1112_w40_10_c9 <= tile_28_filtered_output_c9(1);
   bh1112_w41_9_c9 <= tile_28_filtered_output_c9(2);
   bh1112_w42_11_c9 <= tile_28_filtered_output_c9(3);
   tile_29_X_c5 <= X(8 downto 8);
   tile_29_Y_c9 <= Y(31 downto 31);
   tile_29_mult: IntMultiplierLUT_1x1_Freq300_uid1217
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_29_X_c5,
                 Y => tile_29_Y_c9,
                 R => tile_29_output_c9);

   tile_29_filtered_output_c9 <= unsigned(tile_29_output_c9(0 downto 0));
   bh1112_w39_18_c9 <= tile_29_filtered_output_c9(0);
   tile_30_X_c5 <= X(8 downto 7);
   tile_30_Y_c9 <= Y(32 downto 32);
   tile_30_mult: IntMultiplierLUT_2x1_Freq300_uid1219
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_30_X_c5,
                 Y => tile_30_Y_c9,
                 R => tile_30_output_c9);

   tile_30_filtered_output_c9 <= unsigned(tile_30_output_c9(1 downto 0));
   bh1112_w39_19_c9 <= tile_30_filtered_output_c9(0);
   bh1112_w40_11_c9 <= tile_30_filtered_output_c9(1);
   tile_31_X_c5 <= X(11 downto 9);
   tile_31_Y_c9 <= Y(32 downto 31);
   tile_31_mult: IntMultiplierLUT_3x2_Freq300_uid1221
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_31_X_c5,
                 Y => tile_31_Y_c9,
                 R => tile_31_output_c9);

   tile_31_filtered_output_c9 <= unsigned(tile_31_output_c9(4 downto 0));
   bh1112_w40_12_c9 <= tile_31_filtered_output_c9(0);
   bh1112_w41_10_c9 <= tile_31_filtered_output_c9(1);
   bh1112_w42_12_c9 <= tile_31_filtered_output_c9(2);
   bh1112_w43_10_c9 <= tile_31_filtered_output_c9(3);
   bh1112_w44_9_c9 <= tile_31_filtered_output_c9(4);
   tile_32_X_c5 <= X(5 downto 5);
   tile_32_Y_c9 <= Y(34 downto 34);
   tile_32_mult: IntMultiplierLUT_1x1_Freq300_uid1226
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_32_X_c5,
                 Y => tile_32_Y_c9,
                 R => tile_32_output_c9);

   tile_32_filtered_output_c9 <= unsigned(tile_32_output_c9(0 downto 0));
   bh1112_w39_20_c9 <= tile_32_filtered_output_c9(0);
   tile_33_X_c5 <= X(8 downto 6);
   tile_33_Y_c9 <= Y(34 downto 33);
   tile_33_mult: IntMultiplierLUT_3x2_Freq300_uid1228
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_33_X_c5,
                 Y => tile_33_Y_c9,
                 R => tile_33_output_c9);

   tile_33_filtered_output_c9 <= unsigned(tile_33_output_c9(4 downto 0));
   bh1112_w39_21_c9 <= tile_33_filtered_output_c9(0);
   bh1112_w40_13_c9 <= tile_33_filtered_output_c9(1);
   bh1112_w41_11_c9 <= tile_33_filtered_output_c9(2);
   bh1112_w42_13_c9 <= tile_33_filtered_output_c9(3);
   bh1112_w43_11_c9 <= tile_33_filtered_output_c9(4);
   tile_34_X_c5 <= X(11 downto 9);
   tile_34_Y_c9 <= Y(34 downto 33);
   tile_34_mult: IntMultiplierLUT_3x2_Freq300_uid1233
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_34_X_c5,
                 Y => tile_34_Y_c9,
                 R => tile_34_output_c9);

   tile_34_filtered_output_c9 <= unsigned(tile_34_output_c9(4 downto 0));
   bh1112_w42_14_c9 <= tile_34_filtered_output_c9(0);
   bh1112_w43_12_c9 <= tile_34_filtered_output_c9(1);
   bh1112_w44_10_c9 <= tile_34_filtered_output_c9(2);
   bh1112_w45_8_c9 <= tile_34_filtered_output_c9(3);
   bh1112_w46_8_c9 <= tile_34_filtered_output_c9(4);
   tile_35_X_c5 <= X(3 downto 3);
   tile_35_Y_c9 <= Y(36 downto 36);
   tile_35_mult: IntMultiplierLUT_1x1_Freq300_uid1238
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_35_X_c5,
                 Y => tile_35_Y_c9,
                 R => tile_35_output_c9);

   tile_35_filtered_output_c9 <= unsigned(tile_35_output_c9(0 downto 0));
   bh1112_w39_22_c9 <= tile_35_filtered_output_c9(0);
   tile_36_X_c5 <= X(5 downto 4);
   tile_36_Y_c9 <= Y(36 downto 35);
   tile_36_mult: IntMultiplierLUT_2x2_Freq300_uid1240
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_36_X_c5,
                 Y => tile_36_Y_c9,
                 R => tile_36_output_c9);

   tile_36_filtered_output_c9 <= unsigned(tile_36_output_c9(3 downto 0));
   bh1112_w39_23_c9 <= tile_36_filtered_output_c9(0);
   bh1112_w40_14_c9 <= tile_36_filtered_output_c9(1);
   bh1112_w41_12_c9 <= tile_36_filtered_output_c9(2);
   bh1112_w42_15_c9 <= tile_36_filtered_output_c9(3);
   tile_37_X_c5 <= X(8 downto 6);
   tile_37_Y_c9 <= Y(36 downto 35);
   tile_37_mult: IntMultiplierLUT_3x2_Freq300_uid1245
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_37_X_c5,
                 Y => tile_37_Y_c9,
                 R => tile_37_output_c9);

   tile_37_filtered_output_c9 <= unsigned(tile_37_output_c9(4 downto 0));
   bh1112_w41_13_c9 <= tile_37_filtered_output_c9(0);
   bh1112_w42_16_c9 <= tile_37_filtered_output_c9(1);
   bh1112_w43_13_c9 <= tile_37_filtered_output_c9(2);
   bh1112_w44_11_c9 <= tile_37_filtered_output_c9(3);
   bh1112_w45_9_c9 <= tile_37_filtered_output_c9(4);
   tile_38_X_c5 <= X(11 downto 9);
   tile_38_Y_c9 <= Y(36 downto 35);
   tile_38_mult: IntMultiplierLUT_3x2_Freq300_uid1250
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_38_X_c5,
                 Y => tile_38_Y_c9,
                 R => tile_38_output_c9);

   tile_38_filtered_output_c9 <= unsigned(tile_38_output_c9(4 downto 0));
   bh1112_w44_12_c9 <= tile_38_filtered_output_c9(0);
   bh1112_w45_10_c9 <= tile_38_filtered_output_c9(1);
   bh1112_w46_9_c9 <= tile_38_filtered_output_c9(2);
   bh1112_w47_6_c9 <= tile_38_filtered_output_c9(3);
   bh1112_w48_6_c9 <= tile_38_filtered_output_c9(4);
   tile_39_X_c5 <= X(2 downto 2);
   tile_39_Y_c9 <= Y(37 downto 37);
   tile_39_mult: IntMultiplierLUT_1x1_Freq300_uid1255
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_39_X_c5,
                 Y => tile_39_Y_c9,
                 R => tile_39_output_c9);

   tile_39_filtered_output_c9 <= unsigned(tile_39_output_c9(0 downto 0));
   bh1112_w39_24_c9 <= tile_39_filtered_output_c9(0);
   tile_40_X_c5 <= X(2 downto 1);
   tile_40_Y_c9 <= Y(38 downto 38);
   tile_40_mult: IntMultiplierLUT_2x1_Freq300_uid1257
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_40_X_c5,
                 Y => tile_40_Y_c9,
                 R => tile_40_output_c9);

   tile_40_filtered_output_c9 <= unsigned(tile_40_output_c9(1 downto 0));
   bh1112_w39_25_c9 <= tile_40_filtered_output_c9(0);
   bh1112_w40_15_c9 <= tile_40_filtered_output_c9(1);
   tile_41_X_c5 <= X(5 downto 3);
   tile_41_Y_c9 <= Y(38 downto 37);
   tile_41_mult: IntMultiplierLUT_3x2_Freq300_uid1259
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_41_X_c5,
                 Y => tile_41_Y_c9,
                 R => tile_41_output_c9);

   tile_41_filtered_output_c9 <= unsigned(tile_41_output_c9(4 downto 0));
   bh1112_w40_16_c9 <= tile_41_filtered_output_c9(0);
   bh1112_w41_14_c9 <= tile_41_filtered_output_c9(1);
   bh1112_w42_17_c9 <= tile_41_filtered_output_c9(2);
   bh1112_w43_14_c9 <= tile_41_filtered_output_c9(3);
   bh1112_w44_13_c9 <= tile_41_filtered_output_c9(4);
   tile_42_X_c5 <= X(8 downto 6);
   tile_42_Y_c9 <= Y(38 downto 37);
   tile_42_mult: IntMultiplierLUT_3x2_Freq300_uid1264
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_42_X_c5,
                 Y => tile_42_Y_c9,
                 R => tile_42_output_c9);

   tile_42_filtered_output_c9 <= unsigned(tile_42_output_c9(4 downto 0));
   bh1112_w43_15_c9 <= tile_42_filtered_output_c9(0);
   bh1112_w44_14_c9 <= tile_42_filtered_output_c9(1);
   bh1112_w45_11_c9 <= tile_42_filtered_output_c9(2);
   bh1112_w46_10_c9 <= tile_42_filtered_output_c9(3);
   bh1112_w47_7_c9 <= tile_42_filtered_output_c9(4);
   tile_43_X_c5 <= X(11 downto 9);
   tile_43_Y_c9 <= Y(38 downto 37);
   tile_43_mult: IntMultiplierLUT_3x2_Freq300_uid1269
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_43_X_c5,
                 Y => tile_43_Y_c9,
                 R => tile_43_output_c9);

   tile_43_filtered_output_c9 <= unsigned(tile_43_output_c9(4 downto 0));
   bh1112_w46_11_c9 <= tile_43_filtered_output_c9(0);
   bh1112_w47_8_c9 <= tile_43_filtered_output_c9(1);
   bh1112_w48_7_c9 <= tile_43_filtered_output_c9(2);
   bh1112_w49_5_c9 <= tile_43_filtered_output_c9(3);
   bh1112_w50_4_c9 <= tile_43_filtered_output_c9(4);
   tile_44_X_c5 <= X(2 downto 0);
   tile_44_Y_c9 <= Y(40 downto 39);
   tile_44_mult: IntMultiplierLUT_3x2_Freq300_uid1274
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_44_X_c5,
                 Y => tile_44_Y_c9,
                 R => tile_44_output_c9);

   tile_44_filtered_output_c9 <= unsigned(tile_44_output_c9(4 downto 0));
   bh1112_w39_26_c9 <= tile_44_filtered_output_c9(0);
   bh1112_w40_17_c9 <= tile_44_filtered_output_c9(1);
   bh1112_w41_15_c9 <= tile_44_filtered_output_c9(2);
   bh1112_w42_18_c9 <= tile_44_filtered_output_c9(3);
   bh1112_w43_16_c9 <= tile_44_filtered_output_c9(4);
   tile_45_X_c5 <= X(5 downto 3);
   tile_45_Y_c9 <= Y(40 downto 39);
   tile_45_mult: IntMultiplierLUT_3x2_Freq300_uid1279
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_45_X_c5,
                 Y => tile_45_Y_c9,
                 R => tile_45_output_c9);

   tile_45_filtered_output_c9 <= unsigned(tile_45_output_c9(4 downto 0));
   bh1112_w42_19_c9 <= tile_45_filtered_output_c9(0);
   bh1112_w43_17_c9 <= tile_45_filtered_output_c9(1);
   bh1112_w44_15_c9 <= tile_45_filtered_output_c9(2);
   bh1112_w45_12_c9 <= tile_45_filtered_output_c9(3);
   bh1112_w46_12_c9 <= tile_45_filtered_output_c9(4);
   tile_46_X_c5 <= X(8 downto 6);
   tile_46_Y_c9 <= Y(40 downto 39);
   tile_46_mult: IntMultiplierLUT_3x2_Freq300_uid1284
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_46_X_c5,
                 Y => tile_46_Y_c9,
                 R => tile_46_output_c9);

   tile_46_filtered_output_c9 <= unsigned(tile_46_output_c9(4 downto 0));
   bh1112_w45_13_c9 <= tile_46_filtered_output_c9(0);
   bh1112_w46_13_c9 <= tile_46_filtered_output_c9(1);
   bh1112_w47_9_c9 <= tile_46_filtered_output_c9(2);
   bh1112_w48_8_c9 <= tile_46_filtered_output_c9(3);
   bh1112_w49_6_c9 <= tile_46_filtered_output_c9(4);
   tile_47_X_c5 <= X(11 downto 9);
   tile_47_Y_c9 <= Y(40 downto 39);
   tile_47_mult: IntMultiplierLUT_3x2_Freq300_uid1289
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_47_X_c5,
                 Y => tile_47_Y_c9,
                 R => tile_47_output_c9);

   tile_47_filtered_output_c9 <= unsigned(tile_47_output_c9(4 downto 0));
   bh1112_w48_9_c9 <= tile_47_filtered_output_c9(0);
   bh1112_w49_7_c9 <= tile_47_filtered_output_c9(1);
   bh1112_w50_5_c9 <= tile_47_filtered_output_c9(2);
   bh1112_w51_3_c9 <= tile_47_filtered_output_c9(3);
   bh1112_w52_3_c9 <= tile_47_filtered_output_c9(4);
   tile_48_X_c5 <= X(2 downto 0);
   tile_48_Y_c9 <= Y(42 downto 41);
   tile_48_mult: IntMultiplierLUT_3x2_Freq300_uid1294
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_48_X_c5,
                 Y => tile_48_Y_c9,
                 R => tile_48_output_c9);

   tile_48_filtered_output_c9 <= unsigned(tile_48_output_c9(4 downto 0));
   bh1112_w41_16_c9 <= tile_48_filtered_output_c9(0);
   bh1112_w42_20_c9 <= tile_48_filtered_output_c9(1);
   bh1112_w43_18_c9 <= tile_48_filtered_output_c9(2);
   bh1112_w44_16_c9 <= tile_48_filtered_output_c9(3);
   bh1112_w45_14_c9 <= tile_48_filtered_output_c9(4);
   tile_49_X_c5 <= X(5 downto 3);
   tile_49_Y_c9 <= Y(42 downto 41);
   tile_49_mult: IntMultiplierLUT_3x2_Freq300_uid1299
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_49_X_c5,
                 Y => tile_49_Y_c9,
                 R => tile_49_output_c9);

   tile_49_filtered_output_c9 <= unsigned(tile_49_output_c9(4 downto 0));
   bh1112_w44_17_c9 <= tile_49_filtered_output_c9(0);
   bh1112_w45_15_c9 <= tile_49_filtered_output_c9(1);
   bh1112_w46_14_c9 <= tile_49_filtered_output_c9(2);
   bh1112_w47_10_c9 <= tile_49_filtered_output_c9(3);
   bh1112_w48_10_c9 <= tile_49_filtered_output_c9(4);
   tile_50_X_c5 <= X(8 downto 6);
   tile_50_Y_c9 <= Y(42 downto 41);
   tile_50_mult: IntMultiplierLUT_3x2_Freq300_uid1304
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_50_X_c5,
                 Y => tile_50_Y_c9,
                 R => tile_50_output_c9);

   tile_50_filtered_output_c9 <= unsigned(tile_50_output_c9(4 downto 0));
   bh1112_w47_11_c9 <= tile_50_filtered_output_c9(0);
   bh1112_w48_11_c9 <= tile_50_filtered_output_c9(1);
   bh1112_w49_8_c9 <= tile_50_filtered_output_c9(2);
   bh1112_w50_6_c9 <= tile_50_filtered_output_c9(3);
   bh1112_w51_4_c9 <= tile_50_filtered_output_c9(4);
   tile_51_X_c5 <= X(11 downto 9);
   tile_51_Y_c9 <= Y(42 downto 41);
   tile_51_mult: IntMultiplierLUT_3x2_Freq300_uid1309
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_51_X_c5,
                 Y => tile_51_Y_c9,
                 R => tile_51_output_c9);

   tile_51_filtered_output_c9 <= unsigned(tile_51_output_c9(4 downto 0));
   bh1112_w50_7_c9 <= tile_51_filtered_output_c9(0);
   bh1112_w51_5_c9 <= tile_51_filtered_output_c9(1);
   bh1112_w52_4_c9 <= tile_51_filtered_output_c9(2);
   bh1112_w53_3_c9 <= tile_51_filtered_output_c9(3);
   bh1112_w54_3_c9 <= tile_51_filtered_output_c9(4);
   tile_52_X_c5 <= X(2 downto 0);
   tile_52_Y_c9 <= Y(44 downto 43);
   tile_52_mult: IntMultiplierLUT_3x2_Freq300_uid1314
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_52_X_c5,
                 Y => tile_52_Y_c9,
                 R => tile_52_output_c9);

   tile_52_filtered_output_c9 <= unsigned(tile_52_output_c9(4 downto 0));
   bh1112_w43_19_c9 <= tile_52_filtered_output_c9(0);
   bh1112_w44_18_c9 <= tile_52_filtered_output_c9(1);
   bh1112_w45_16_c9 <= tile_52_filtered_output_c9(2);
   bh1112_w46_15_c9 <= tile_52_filtered_output_c9(3);
   bh1112_w47_12_c9 <= tile_52_filtered_output_c9(4);
   tile_53_X_c5 <= X(5 downto 3);
   tile_53_Y_c9 <= Y(44 downto 43);
   tile_53_mult: IntMultiplierLUT_3x2_Freq300_uid1319
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_53_X_c5,
                 Y => tile_53_Y_c9,
                 R => tile_53_output_c9);

   tile_53_filtered_output_c9 <= unsigned(tile_53_output_c9(4 downto 0));
   bh1112_w46_16_c9 <= tile_53_filtered_output_c9(0);
   bh1112_w47_13_c9 <= tile_53_filtered_output_c9(1);
   bh1112_w48_12_c9 <= tile_53_filtered_output_c9(2);
   bh1112_w49_9_c9 <= tile_53_filtered_output_c9(3);
   bh1112_w50_8_c9 <= tile_53_filtered_output_c9(4);
   tile_54_X_c5 <= X(8 downto 6);
   tile_54_Y_c9 <= Y(44 downto 43);
   tile_54_mult: IntMultiplierLUT_3x2_Freq300_uid1324
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_54_X_c5,
                 Y => tile_54_Y_c9,
                 R => tile_54_output_c9);

   tile_54_filtered_output_c9 <= unsigned(tile_54_output_c9(4 downto 0));
   bh1112_w49_10_c9 <= tile_54_filtered_output_c9(0);
   bh1112_w50_9_c9 <= tile_54_filtered_output_c9(1);
   bh1112_w51_6_c9 <= tile_54_filtered_output_c9(2);
   bh1112_w52_5_c9 <= tile_54_filtered_output_c9(3);
   bh1112_w53_4_c9 <= tile_54_filtered_output_c9(4);
   tile_55_X_c5 <= X(11 downto 9);
   tile_55_Y_c9 <= Y(44 downto 43);
   tile_55_mult: IntMultiplierLUT_3x2_Freq300_uid1329
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_55_X_c5,
                 Y => tile_55_Y_c9,
                 R => tile_55_output_c9);

   tile_55_filtered_output_c9 <= unsigned(tile_55_output_c9(4 downto 0));
   bh1112_w52_6_c9 <= tile_55_filtered_output_c9(0);
   bh1112_w53_5_c9 <= tile_55_filtered_output_c9(1);
   bh1112_w54_4_c9 <= tile_55_filtered_output_c9(2);
   bh1112_w55_3_c9 <= tile_55_filtered_output_c9(3);
   bh1112_w56_3_c9 <= tile_55_filtered_output_c9(4);
   tile_56_X_c5 <= X(2 downto 0);
   tile_56_Y_c9 <= Y(46 downto 45);
   tile_56_mult: IntMultiplierLUT_3x2_Freq300_uid1334
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_56_X_c5,
                 Y => tile_56_Y_c9,
                 R => tile_56_output_c9);

   tile_56_filtered_output_c9 <= unsigned(tile_56_output_c9(4 downto 0));
   bh1112_w45_17_c9 <= tile_56_filtered_output_c9(0);
   bh1112_w46_17_c9 <= tile_56_filtered_output_c9(1);
   bh1112_w47_14_c9 <= tile_56_filtered_output_c9(2);
   bh1112_w48_13_c9 <= tile_56_filtered_output_c9(3);
   bh1112_w49_11_c9 <= tile_56_filtered_output_c9(4);
   tile_57_X_c5 <= X(5 downto 3);
   tile_57_Y_c9 <= Y(46 downto 45);
   tile_57_mult: IntMultiplierLUT_3x2_Freq300_uid1339
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_57_X_c5,
                 Y => tile_57_Y_c9,
                 R => tile_57_output_c9);

   tile_57_filtered_output_c9 <= unsigned(tile_57_output_c9(4 downto 0));
   bh1112_w48_14_c9 <= tile_57_filtered_output_c9(0);
   bh1112_w49_12_c9 <= tile_57_filtered_output_c9(1);
   bh1112_w50_10_c9 <= tile_57_filtered_output_c9(2);
   bh1112_w51_7_c9 <= tile_57_filtered_output_c9(3);
   bh1112_w52_7_c9 <= tile_57_filtered_output_c9(4);
   tile_58_X_c5 <= X(8 downto 6);
   tile_58_Y_c9 <= Y(46 downto 45);
   tile_58_mult: IntMultiplierLUT_3x2_Freq300_uid1344
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_58_X_c5,
                 Y => tile_58_Y_c9,
                 R => tile_58_output_c9);

   tile_58_filtered_output_c9 <= unsigned(tile_58_output_c9(4 downto 0));
   bh1112_w51_8_c9 <= tile_58_filtered_output_c9(0);
   bh1112_w52_8_c9 <= tile_58_filtered_output_c9(1);
   bh1112_w53_6_c9 <= tile_58_filtered_output_c9(2);
   bh1112_w54_5_c9 <= tile_58_filtered_output_c9(3);
   bh1112_w55_4_c9 <= tile_58_filtered_output_c9(4);
   tile_59_X_c5 <= X(11 downto 9);
   tile_59_Y_c9 <= Y(46 downto 45);
   tile_59_mult: IntMultiplierLUT_3x2_Freq300_uid1349
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 X => tile_59_X_c5,
                 Y => tile_59_Y_c9,
                 R => tile_59_output_c9);

   tile_59_filtered_output_c9 <= unsigned(tile_59_output_c9(4 downto 0));
   bh1112_w54_6_c9 <= tile_59_filtered_output_c9(0);
   bh1112_w55_5_c9 <= tile_59_filtered_output_c9(1);
   bh1112_w56_4_c9 <= tile_59_filtered_output_c9(2);
   bh1112_w57_3_c9 <= tile_59_filtered_output_c9(3);
   bh1112_w58_3_c9 <= tile_59_filtered_output_c9(4);

   -- Adding the constant bits 
   bh1112_w39_27_c0 <= '1';
   bh1112_w40_18_c0 <= '1';
   bh1112_w41_17_c0 <= '1';
   bh1112_w42_21_c0 <= '1';
   bh1112_w43_20_c0 <= '1';
   bh1112_w44_19_c0 <= '1';


   Compressor_23_3_Freq300_uid1355_bh1112_uid1356_In0_c9 <= "" & bh1112_w36_0_c9 & bh1112_w36_1_c9 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1356_In1_c9 <= "" & bh1112_w37_0_c9 & bh1112_w37_1_c9;
   bh1112_w36_2_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_c10(0);
   bh1112_w37_2_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_c10(1);
   bh1112_w38_2_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1356: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1356_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1356_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_copy1357_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1356_Out0_copy1357_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1360_In0_c9 <= "" & bh1112_w38_0_c9 & bh1112_w38_1_c9 & "0";
   bh1112_w38_3_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_c10(0);
   bh1112_w39_28_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1360: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1360_In0_c9,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_copy1361_c9);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1360_Out0_copy1361_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1364_In0_c9 <= "" & bh1112_w39_14_c9 & bh1112_w39_27_c9 & bh1112_w39_26_c9 & bh1112_w39_25_c9 & bh1112_w39_24_c9 & bh1112_w39_23_c9;
   bh1112_w39_29_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_c10(0);
   bh1112_w40_19_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_c10(1);
   bh1112_w41_18_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1364: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1364_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_copy1365_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1364_Out0_copy1365_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1366_In0_c9 <= "" & bh1112_w39_0_c9 & bh1112_w39_1_c9 & bh1112_w39_2_c9 & bh1112_w39_3_c9 & bh1112_w39_4_c9 & bh1112_w39_5_c9;
   bh1112_w39_30_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_c10(0);
   bh1112_w40_20_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_c10(1);
   bh1112_w41_19_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1366: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1366_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_copy1367_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1366_Out0_copy1367_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1368_In0_c9 <= "" & bh1112_w39_22_c9 & bh1112_w39_21_c9 & bh1112_w39_20_c9 & bh1112_w39_19_c9 & bh1112_w39_18_c9 & bh1112_w39_17_c9;
   bh1112_w39_31_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1368_Out0_c9(0);
   bh1112_w40_21_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1368_Out0_c9(1);
   bh1112_w41_20_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1368_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1368: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1368_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1368_Out0_copy1369_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1368_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1368_Out0_copy1369_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1370_In0_c9 <= "" & bh1112_w39_6_c9 & bh1112_w39_7_c9 & bh1112_w39_8_c9 & bh1112_w39_9_c9 & bh1112_w39_10_c9 & bh1112_w39_11_c9;
   bh1112_w39_32_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1370_Out0_c9(0);
   bh1112_w40_22_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1370_Out0_c9(1);
   bh1112_w41_21_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1370_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1370: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1370_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1370_Out0_copy1371_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1370_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1370_Out0_copy1371_c9; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1374_In0_c9 <= "" & bh1112_w39_15_c9 & bh1112_w39_16_c9 & bh1112_w39_13_c9 & bh1112_w39_12_c9;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1374_In1_c9 <= "" & bh1112_w40_0_c9;
   bh1112_w39_33_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_c10(0);
   bh1112_w40_23_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_c10(1);
   bh1112_w41_22_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1374: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1374_In0_c9,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1374_In1_c9,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_copy1375_c9);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1374_Out0_copy1375_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1376_In0_c9 <= "" & bh1112_w40_10_c9 & bh1112_w40_1_c9 & bh1112_w40_2_c9 & bh1112_w40_3_c9 & bh1112_w40_4_c9 & bh1112_w40_5_c9;
   bh1112_w40_24_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1376_Out0_c9(0);
   bh1112_w41_23_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1376_Out0_c9(1);
   bh1112_w42_22_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1376_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1376: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1376_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1376_Out0_copy1377_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1376_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1376_Out0_copy1377_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1378_In0_c9 <= "" & bh1112_w40_18_c9 & bh1112_w40_17_c9 & bh1112_w40_16_c9 & bh1112_w40_15_c9 & bh1112_w40_14_c9 & bh1112_w40_13_c9;
   bh1112_w40_25_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1378_Out0_c9(0);
   bh1112_w41_24_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1378_Out0_c9(1);
   bh1112_w42_23_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1378_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1378: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1378_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1378_Out0_copy1379_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1378_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1378_Out0_copy1379_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1380_In0_c9 <= "" & bh1112_w40_6_c9 & bh1112_w40_7_c9 & bh1112_w40_8_c9 & bh1112_w40_9_c9 & bh1112_w40_11_c9 & bh1112_w40_12_c9;
   bh1112_w40_26_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_c10(0);
   bh1112_w41_25_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_c10(1);
   bh1112_w42_24_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1380: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1380_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_copy1381_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1380_Out0_copy1381_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1382_In0_c9 <= "" & bh1112_w41_9_c9 & bh1112_w41_17_c9 & bh1112_w41_16_c9 & bh1112_w41_15_c9 & bh1112_w41_14_c9 & bh1112_w41_13_c9;
   bh1112_w41_26_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1382_Out0_c9(0);
   bh1112_w42_25_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1382_Out0_c9(1);
   bh1112_w43_21_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1382_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1382: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1382_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1382_Out0_copy1383_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1382_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1382_Out0_copy1383_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1384_In0_c9 <= "" & bh1112_w41_0_c9 & bh1112_w41_1_c9 & bh1112_w41_2_c9 & bh1112_w41_3_c9 & bh1112_w41_4_c9 & bh1112_w41_5_c9;
   bh1112_w41_27_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_c10(0);
   bh1112_w42_26_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_c10(1);
   bh1112_w43_22_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1384: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1384_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_copy1385_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1384_Out0_copy1385_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1386_In0_c9 <= "" & bh1112_w41_12_c9 & bh1112_w41_11_c9 & bh1112_w41_10_c9 & bh1112_w41_8_c9 & bh1112_w41_7_c9 & bh1112_w41_6_c9;
   bh1112_w41_28_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_c10(0);
   bh1112_w42_27_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_c10(1);
   bh1112_w43_23_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1386: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1386_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_copy1387_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1386_Out0_copy1387_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1388_In0_c9 <= "" & bh1112_w42_0_c9 & bh1112_w42_1_c9 & bh1112_w42_2_c9 & bh1112_w42_3_c9 & bh1112_w42_4_c9 & bh1112_w42_5_c9;
   bh1112_w42_28_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_c10(0);
   bh1112_w43_24_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_c10(1);
   bh1112_w44_20_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1388: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1388_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_copy1389_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1388_Out0_copy1389_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1390_In0_c9 <= "" & bh1112_w42_11_c9 & bh1112_w42_21_c9 & bh1112_w42_20_c9 & bh1112_w42_19_c9 & bh1112_w42_18_c9 & bh1112_w42_17_c9;
   bh1112_w42_29_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1390_Out0_c9(0);
   bh1112_w43_25_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1390_Out0_c9(1);
   bh1112_w44_21_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1390_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1390: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1390_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1390_Out0_copy1391_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1390_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1390_Out0_copy1391_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1392_In0_c9 <= "" & bh1112_w42_6_c9 & bh1112_w42_7_c9 & bh1112_w42_8_c9 & bh1112_w42_9_c9 & bh1112_w42_10_c9 & bh1112_w42_12_c9;
   bh1112_w42_30_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_c10(0);
   bh1112_w43_26_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_c10(1);
   bh1112_w44_22_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1392: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1392_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_copy1393_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1392_Out0_copy1393_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In0_c9 <= "" & bh1112_w42_16_c9 & bh1112_w42_15_c9 & bh1112_w42_14_c9 & bh1112_w42_13_c9;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c0 <= "" & "0";
   bh1112_w42_31_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1394_Out0_c9(0);
   bh1112_w43_27_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1394_Out0_c9(1);
   bh1112_w44_23_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1394_Out0_c9(2);
   Compressor_14_3_Freq300_uid1373_uid1394: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In0_c9,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1394_In1_c9,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1394_Out0_copy1395_c9);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1394_Out0_c9 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1394_Out0_copy1395_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1396_In0_c9 <= "" & bh1112_w43_10_c9 & bh1112_w43_1_c9 & bh1112_w43_2_c9 & bh1112_w43_3_c9 & bh1112_w43_4_c9 & bh1112_w43_5_c9;
   bh1112_w43_28_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1396_Out0_c9(0);
   bh1112_w44_24_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1396_Out0_c9(1);
   bh1112_w45_18_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1396_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1396: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1396_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1396_Out0_copy1397_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1396_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1396_Out0_copy1397_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1398_In0_c9 <= "" & bh1112_w43_11_c9 & bh1112_w43_20_c9 & bh1112_w43_19_c9 & bh1112_w43_18_c9 & bh1112_w43_17_c9 & bh1112_w43_16_c9;
   bh1112_w43_29_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1398_Out0_c9(0);
   bh1112_w44_25_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1398_Out0_c9(1);
   bh1112_w45_19_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1398_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1398: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1398_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1398_Out0_copy1399_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1398_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1398_Out0_copy1399_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1400_In0_c9 <= "" & bh1112_w43_6_c9 & bh1112_w43_7_c9 & bh1112_w43_8_c9 & bh1112_w43_9_c9 & bh1112_w43_0_c9 & bh1112_w43_12_c9;
   bh1112_w43_30_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_c10(0);
   bh1112_w44_26_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_c10(1);
   bh1112_w45_20_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1400: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1400_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_copy1401_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1400_Out0_copy1401_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1402_In0_c9 <= "" & bh1112_w43_15_c9 & bh1112_w43_14_c9 & bh1112_w43_13_c9;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1402_In1_c9 <= "" & bh1112_w44_10_c9 & bh1112_w44_19_c9;
   bh1112_w43_31_c9 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1402_Out0_c9(0);
   bh1112_w44_27_c9 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1402_Out0_c9(1);
   bh1112_w45_21_c9 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1402_Out0_c9(2);
   Compressor_23_3_Freq300_uid1355_uid1402: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1402_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1402_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1402_Out0_copy1403_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1402_Out0_c9 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1402_Out0_copy1403_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1404_In0_c9 <= "" & bh1112_w44_0_c9 & bh1112_w44_1_c9 & bh1112_w44_2_c9 & bh1112_w44_3_c9 & bh1112_w44_4_c9 & bh1112_w44_5_c9;
   bh1112_w44_28_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_c10(0);
   bh1112_w45_22_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_c10(1);
   bh1112_w46_18_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1404: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1404_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_copy1405_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1404_Out0_copy1405_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1406_In0_c9 <= "" & bh1112_w44_18_c9 & bh1112_w44_17_c9 & bh1112_w44_16_c9 & bh1112_w44_15_c9 & bh1112_w44_14_c9 & bh1112_w44_13_c9;
   bh1112_w44_29_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1406_Out0_c9(0);
   bh1112_w45_23_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1406_Out0_c9(1);
   bh1112_w46_19_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1406_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1406: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1406_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1406_Out0_copy1407_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1406_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1406_Out0_copy1407_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1408_In0_c9 <= "" & bh1112_w44_6_c9 & bh1112_w44_7_c9 & bh1112_w44_8_c9 & bh1112_w44_9_c9 & bh1112_w44_11_c9 & bh1112_w44_12_c9;
   bh1112_w44_30_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_c10(0);
   bh1112_w45_24_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_c10(1);
   bh1112_w46_20_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1408: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1408_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_copy1409_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1408_Out0_copy1409_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1410_In0_c9 <= "" & bh1112_w45_9_c9 & bh1112_w45_17_c9 & bh1112_w45_16_c9 & bh1112_w45_15_c9 & bh1112_w45_14_c9 & bh1112_w45_13_c9;
   bh1112_w45_25_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1410_Out0_c9(0);
   bh1112_w46_21_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1410_Out0_c9(1);
   bh1112_w47_15_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1410_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1410: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1410_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1410_Out0_copy1411_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1410_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1410_Out0_copy1411_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1412_In0_c9 <= "" & bh1112_w45_0_c9 & bh1112_w45_1_c9 & bh1112_w45_2_c9 & bh1112_w45_3_c9 & bh1112_w45_4_c9 & bh1112_w45_5_c9;
   bh1112_w45_26_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_c10(0);
   bh1112_w46_22_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_c10(1);
   bh1112_w47_16_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1412: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1412_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_copy1413_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1412_Out0_copy1413_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1414_In0_c9 <= "" & bh1112_w45_12_c9 & bh1112_w45_11_c9 & bh1112_w45_10_c9 & bh1112_w45_8_c9 & bh1112_w45_7_c9 & bh1112_w45_6_c9;
   bh1112_w45_27_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_c10(0);
   bh1112_w46_23_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_c10(1);
   bh1112_w47_17_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1414: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1414_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_copy1415_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1414_Out0_copy1415_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1416_In0_c9 <= "" & bh1112_w46_0_c9 & bh1112_w46_1_c9 & bh1112_w46_2_c9 & bh1112_w46_3_c9 & bh1112_w46_4_c9 & bh1112_w46_5_c9;
   bh1112_w46_24_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_c10(0);
   bh1112_w47_18_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_c10(1);
   bh1112_w48_15_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1416: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1416_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_copy1417_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1416_Out0_copy1417_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1418_In0_c9 <= "" & bh1112_w46_9_c9 & bh1112_w46_17_c9 & bh1112_w46_16_c9 & bh1112_w46_15_c9 & bh1112_w46_14_c9 & bh1112_w46_13_c9;
   bh1112_w46_25_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1418_Out0_c9(0);
   bh1112_w47_19_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1418_Out0_c9(1);
   bh1112_w48_16_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1418_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1418: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1418_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1418_Out0_copy1419_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1418_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1418_Out0_copy1419_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1420_In0_c9 <= "" & bh1112_w46_6_c9 & bh1112_w46_7_c9 & bh1112_w46_8_c9 & bh1112_w46_10_c9 & bh1112_w46_11_c9 & bh1112_w46_12_c9;
   bh1112_w46_26_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_c10(0);
   bh1112_w47_20_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_c10(1);
   bh1112_w48_17_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1420: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1420_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_copy1421_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1420_Out0_copy1421_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1422_In0_c9 <= "" & bh1112_w47_8_c9 & bh1112_w47_14_c9 & bh1112_w47_13_c9 & bh1112_w47_12_c9 & bh1112_w47_11_c9 & bh1112_w47_10_c9;
   bh1112_w47_21_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1422_Out0_c9(0);
   bh1112_w48_18_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1422_Out0_c9(1);
   bh1112_w49_13_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1422_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1422: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1422_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1422_Out0_copy1423_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1422_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1422_Out0_copy1423_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1424_In0_c9 <= "" & bh1112_w47_0_c9 & bh1112_w47_1_c9 & bh1112_w47_2_c9 & bh1112_w47_3_c9 & bh1112_w47_4_c9 & bh1112_w47_5_c9;
   bh1112_w47_22_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_c10(0);
   bh1112_w48_19_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_c10(1);
   bh1112_w49_14_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1424: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1424_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_copy1425_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1424_Out0_copy1425_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1426_In0_c9 <= "" & bh1112_w47_9_c9 & bh1112_w47_7_c9 & bh1112_w47_6_c9;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1426_In1_c9 <= "" & bh1112_w48_0_c9 & bh1112_w48_1_c9;
   bh1112_w47_23_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_c10(0);
   bh1112_w48_20_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_c10(1);
   bh1112_w49_15_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1426: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1426_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1426_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_copy1427_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1426_Out0_copy1427_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1428_In0_c9 <= "" & bh1112_w48_8_c9 & bh1112_w48_14_c9 & bh1112_w48_13_c9 & bh1112_w48_12_c9 & bh1112_w48_11_c9 & bh1112_w48_10_c9;
   bh1112_w48_21_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1428_Out0_c9(0);
   bh1112_w49_16_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1428_Out0_c9(1);
   bh1112_w50_11_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1428_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1428: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1428_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1428_Out0_copy1429_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1428_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1428_Out0_copy1429_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1430_In0_c9 <= "" & bh1112_w48_2_c9 & bh1112_w48_3_c9 & bh1112_w48_4_c9 & bh1112_w48_5_c9 & bh1112_w48_6_c9 & bh1112_w48_7_c9;
   bh1112_w48_22_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_c10(0);
   bh1112_w49_17_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_c10(1);
   bh1112_w50_12_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1430: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1430_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_copy1431_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1430_Out0_copy1431_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1432_In0_c9 <= "" & bh1112_w49_0_c9 & bh1112_w49_1_c9 & bh1112_w49_2_c9 & bh1112_w49_3_c9 & bh1112_w49_4_c9 & bh1112_w49_5_c9;
   bh1112_w49_18_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_c10(0);
   bh1112_w50_13_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_c10(1);
   bh1112_w51_9_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1432: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1432_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_copy1433_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1432_Out0_copy1433_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1434_In0_c9 <= "" & bh1112_w49_8_c9 & bh1112_w49_12_c9 & bh1112_w49_11_c9 & bh1112_w49_10_c9 & bh1112_w49_9_c9 & bh1112_w49_7_c9;
   bh1112_w49_19_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1434_Out0_c9(0);
   bh1112_w50_14_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1434_Out0_c9(1);
   bh1112_w51_10_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1434_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1434: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1434_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1434_Out0_copy1435_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1434_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1434_Out0_copy1435_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1436_In0_c9 <= "" & bh1112_w50_0_c9 & bh1112_w50_1_c9 & bh1112_w50_2_c9 & bh1112_w50_3_c9 & "0" & "0";
   bh1112_w50_15_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_c10(0);
   bh1112_w51_11_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_c10(1);
   bh1112_w52_9_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1436: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1436_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_copy1437_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1436_Out0_copy1437_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1438_In0_c9 <= "" & bh1112_w50_4_c9 & bh1112_w50_5_c9 & bh1112_w50_6_c9 & bh1112_w50_7_c9;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1438_In1_c9 <= "" & bh1112_w51_0_c9;
   bh1112_w50_16_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_c10(0);
   bh1112_w51_12_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_c10(1);
   bh1112_w52_10_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1438: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1438_In0_c9,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1438_In1_c9,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_copy1439_c9);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1438_Out0_copy1439_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1440_In0_c9 <= "" & bh1112_w50_8_c9 & bh1112_w50_10_c9 & bh1112_w50_9_c9;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1440_In1_c9 <= "" & bh1112_w51_1_c9 & bh1112_w51_2_c9;
   bh1112_w50_17_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_c10(0);
   bh1112_w51_13_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_c10(1);
   bh1112_w52_11_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1440: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1440_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1440_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_copy1441_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1440_Out0_copy1441_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1442_In0_c9 <= "" & bh1112_w51_3_c9 & bh1112_w51_4_c9 & bh1112_w51_5_c9 & bh1112_w51_6_c9 & bh1112_w51_7_c9 & bh1112_w51_8_c9;
   bh1112_w51_14_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1442_Out0_c9(0);
   bh1112_w52_12_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1442_Out0_c9(1);
   bh1112_w53_7_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1442_Out0_c9(2);
   Compressor_6_3_Freq300_uid1363_uid1442: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1442_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1442_Out0_copy1443_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1442_Out0_c9 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1442_Out0_copy1443_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1444_In0_c9 <= "" & bh1112_w52_0_c9 & bh1112_w52_1_c9 & bh1112_w52_2_c9 & bh1112_w52_3_c9 & bh1112_w52_4_c9 & bh1112_w52_5_c9;
   bh1112_w52_13_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_c10(0);
   bh1112_w53_8_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_c10(1);
   bh1112_w54_7_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1444: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1444_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_copy1445_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1444_Out0_copy1445_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1446_In0_c9 <= "" & bh1112_w52_6_c9 & bh1112_w52_7_c9 & bh1112_w52_8_c9;
   bh1112_w52_14_c9 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1446_Out0_c9(0);
   bh1112_w53_9_c9 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1446_Out0_c9(1);
   Compressor_3_2_Freq300_uid1359_uid1446: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1446_In0_c9,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1446_Out0_copy1447_c9);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1446_Out0_c9 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1446_Out0_copy1447_c9; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1448_In0_c9 <= "" & bh1112_w53_0_c9 & bh1112_w53_1_c9 & bh1112_w53_2_c9 & bh1112_w53_3_c9 & bh1112_w53_4_c9 & bh1112_w53_5_c9;
   bh1112_w53_10_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_c10(0);
   bh1112_w54_8_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_c10(1);
   bh1112_w55_6_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1448: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1448_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_copy1449_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1448_Out0_copy1449_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1450_In0_c9 <= "" & bh1112_w54_0_c9 & bh1112_w54_1_c9 & bh1112_w54_2_c9 & bh1112_w54_3_c9 & bh1112_w54_4_c9 & bh1112_w54_5_c9;
   bh1112_w54_9_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_c10(0);
   bh1112_w55_7_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_c10(1);
   bh1112_w56_5_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1450: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1450_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_copy1451_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1450_Out0_copy1451_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1452_In0_c9 <= "" & bh1112_w55_0_c9 & bh1112_w55_1_c9 & bh1112_w55_2_c9 & bh1112_w55_3_c9 & bh1112_w55_4_c9 & bh1112_w55_5_c9;
   bh1112_w55_8_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_c10(0);
   bh1112_w56_6_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_c10(1);
   bh1112_w57_4_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1452: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1452_In0_c9,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_copy1453_c9);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1452_Out0_copy1453_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1454_In0_c9 <= "" & bh1112_w56_0_c9 & bh1112_w56_1_c9 & bh1112_w56_2_c9 & bh1112_w56_3_c9;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1454_In1_c9 <= "" & bh1112_w57_0_c9;
   bh1112_w56_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_c10(0);
   bh1112_w57_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_c10(1);
   bh1112_w58_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1454: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1454_In0_c9,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1454_In1_c9,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_copy1455_c9);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1454_Out0_copy1455_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1456_In0_c9 <= "" & bh1112_w57_1_c9 & bh1112_w57_2_c9 & bh1112_w57_3_c9;
   bh1112_w57_6_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_c10(0);
   bh1112_w58_5_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1456: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1456_In0_c9,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_copy1457_c9);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1456_Out0_copy1457_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In0_c9 <= "" & bh1112_w58_0_c9 & bh1112_w58_1_c9 & bh1112_w58_2_c9 & bh1112_w58_3_c9;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c0 <= "" & "0";
   bh1112_w58_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_c10(0);
   bh1112_w59_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_c10(1);
   bh1112_w60_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1458: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In0_c9,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1458_In1_c9,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_copy1459_c9);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1458_Out0_copy1459_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1460_In0_c9 <= "" & bh1112_w59_0_c9 & bh1112_w59_1_c9 & bh1112_w59_2_c9;
   bh1112_w59_4_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_c10(0);
   bh1112_w60_4_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1460: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1460_In0_c9,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_copy1461_c9);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1460_Out0_copy1461_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1462_In0_c9 <= "" & bh1112_w60_0_c9 & bh1112_w60_1_c9 & bh1112_w60_2_c9;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1462_In1_c9 <= "" & bh1112_w61_0_c9 & bh1112_w61_1_c9;
   bh1112_w60_5_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_c10(0);
   bh1112_w61_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_c10(1);
   bh1112_w62_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1462: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1462_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1462_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_copy1463_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1462_Out0_copy1463_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1464_In0_c9 <= "" & bh1112_w62_0_c9 & bh1112_w62_1_c9 & bh1112_w62_2_c9;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1464_In1_c9 <= "" & bh1112_w63_0_c9 & bh1112_w63_1_c9;
   bh1112_w62_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_c10(0);
   bh1112_w63_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_c10(1);
   bh1112_w64_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1464: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1464_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1464_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_copy1465_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1464_Out0_copy1465_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1466_In0_c9 <= "" & bh1112_w64_0_c9 & bh1112_w64_1_c9 & bh1112_w64_2_c9;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1466_In1_c9 <= "" & bh1112_w65_0_c9 & bh1112_w65_1_c9;
   bh1112_w64_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_c10(0);
   bh1112_w65_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_c10(1);
   bh1112_w66_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1466: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1466_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1466_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_copy1467_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1466_Out0_copy1467_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1468_In0_c9 <= "" & bh1112_w66_0_c9 & bh1112_w66_1_c9 & bh1112_w66_2_c9;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1468_In1_c9 <= "" & bh1112_w67_0_c9 & bh1112_w67_1_c9;
   bh1112_w66_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_c10(0);
   bh1112_w67_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_c10(1);
   bh1112_w68_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1468: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1468_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1468_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_copy1469_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1468_Out0_copy1469_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1470_In0_c9 <= "" & bh1112_w68_0_c9 & bh1112_w68_1_c9 & bh1112_w68_2_c9;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1470_In1_c9 <= "" & bh1112_w69_0_c9 & bh1112_w69_1_c9;
   bh1112_w68_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_c10(0);
   bh1112_w69_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_c10(1);
   bh1112_w70_2_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1470: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1470_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1470_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_copy1471_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1470_Out0_copy1471_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1472_In0_c9 <= "" & bh1112_w70_0_c9 & bh1112_w70_1_c9 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1472_In1_c9 <= "" & bh1112_w71_0_c9 & bh1112_w71_1_c9;
   bh1112_w70_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_c10(0);
   bh1112_w71_2_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_c10(1);
   bh1112_w72_2_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1472: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1472_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1472_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_copy1473_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1472_Out0_copy1473_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1474_In0_c9 <= "" & bh1112_w72_0_c9 & bh1112_w72_1_c9 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1474_In1_c9 <= "" & bh1112_w73_0_c9 & bh1112_w73_1_c9;
   bh1112_w72_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_c10(0);
   bh1112_w73_2_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_c10(1);
   bh1112_w74_2_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1474: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1474_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1474_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_copy1475_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1474_Out0_copy1475_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1476_In0_c9 <= "" & bh1112_w74_0_c9 & bh1112_w74_1_c9 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1476_In1_c9 <= "" & bh1112_w75_0_c9 & bh1112_w75_1_c9;
   bh1112_w74_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_c10(0);
   bh1112_w75_2_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_c10(1);
   bh1112_w76_1_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1476: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1476_In0_c9,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1476_In1_c9,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_copy1477_c9);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1476_Out0_copy1477_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1478_In0_c10 <= "" & bh1112_w37_2_c10 & "0" & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1478_In1_c10 <= "" & bh1112_w38_2_c10 & bh1112_w38_3_c10;
   bh1112_w37_3_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1478_Out0_c10(0);
   bh1112_w38_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1478_Out0_c10(1);
   bh1112_w39_34_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1478_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1478: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1478_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1478_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1478_Out0_copy1479_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1478_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1478_Out0_copy1479_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1480_In0_c10 <= "" & bh1112_w39_28_c10 & bh1112_w39_30_c10 & bh1112_w39_32_c10 & bh1112_w39_29_c10 & bh1112_w39_31_c10 & bh1112_w39_33_c10;
   bh1112_w39_35_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1480_Out0_c10(0);
   bh1112_w40_27_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1480_Out0_c10(1);
   bh1112_w41_29_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1480_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1480: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1480_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1480_Out0_copy1481_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1480_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1480_Out0_copy1481_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1482_In0_c10 <= "" & bh1112_w40_26_c10 & bh1112_w40_24_c10 & bh1112_w40_22_c10 & bh1112_w40_20_c10 & "0" & "0";
   bh1112_w40_28_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1482_Out0_c10(0);
   bh1112_w41_30_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1482_Out0_c10(1);
   bh1112_w42_32_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1482_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1482: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1482_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1482_Out0_copy1483_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1482_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1482_Out0_copy1483_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1484_In0_c10 <= "" & bh1112_w40_19_c10 & bh1112_w40_21_c10 & bh1112_w40_23_c10 & bh1112_w40_25_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1484_In1_c10 <= "" & bh1112_w41_27_c10;
   bh1112_w40_29_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1484_Out0_c10(0);
   bh1112_w41_31_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1484_Out0_c10(1);
   bh1112_w42_33_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1484_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1484: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1484_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1484_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1484_Out0_copy1485_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1484_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1484_Out0_copy1485_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1486_In0_c10 <= "" & bh1112_w41_25_c10 & bh1112_w41_23_c10 & bh1112_w41_21_c10 & bh1112_w41_19_c10 & bh1112_w41_18_c10 & bh1112_w41_20_c10;
   bh1112_w41_32_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1486_Out0_c10(0);
   bh1112_w42_34_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1486_Out0_c10(1);
   bh1112_w43_32_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1486_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1486: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1486_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1486_Out0_copy1487_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1486_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1486_Out0_copy1487_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1488_In0_c10 <= "" & bh1112_w41_22_c10 & bh1112_w41_24_c10 & bh1112_w41_26_c10 & bh1112_w41_28_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1488_In1_c10 <= "" & bh1112_w42_30_c10;
   bh1112_w41_33_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1488_Out0_c10(0);
   bh1112_w42_35_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1488_Out0_c10(1);
   bh1112_w43_33_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1488_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1488: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1488_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1488_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1488_Out0_copy1489_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1488_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1488_Out0_copy1489_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1490_In0_c10 <= "" & bh1112_w42_28_c10 & bh1112_w42_26_c10 & bh1112_w42_24_c10 & bh1112_w42_22_c10 & bh1112_w42_23_c10 & bh1112_w42_25_c10;
   bh1112_w42_36_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1490_Out0_c10(0);
   bh1112_w43_34_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1490_Out0_c10(1);
   bh1112_w44_31_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1490_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1490: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1490_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1490_Out0_copy1491_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1490_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1490_Out0_copy1491_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1492_In0_c10 <= "" & bh1112_w42_27_c10 & bh1112_w42_29_c10 & bh1112_w42_31_c10;
   bh1112_w42_37_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1492_Out0_c10(0);
   bh1112_w43_35_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1492_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1492: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1492_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1492_Out0_copy1493_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1492_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1492_Out0_copy1493_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1494_In0_c10 <= "" & bh1112_w43_30_c10 & bh1112_w43_28_c10 & bh1112_w43_26_c10 & bh1112_w43_24_c10 & bh1112_w43_22_c10 & bh1112_w43_21_c10;
   bh1112_w43_36_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1494_Out0_c10(0);
   bh1112_w44_32_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1494_Out0_c10(1);
   bh1112_w45_28_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1494_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1494: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1494_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1494_Out0_copy1495_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1494_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1494_Out0_copy1495_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1496_In0_c10 <= "" & bh1112_w43_23_c10 & bh1112_w43_25_c10 & bh1112_w43_27_c10 & bh1112_w43_29_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1496_In1_c10 <= "" & bh1112_w44_30_c10;
   bh1112_w43_37_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1496_Out0_c10(0);
   bh1112_w44_33_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1496_Out0_c10(1);
   bh1112_w45_29_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1496_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1496: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1496_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1496_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1496_Out0_copy1497_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1496_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1496_Out0_copy1497_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1498_In0_c10 <= "" & bh1112_w44_28_c10 & bh1112_w44_26_c10 & bh1112_w44_24_c10 & bh1112_w44_22_c10 & bh1112_w44_20_c10 & bh1112_w44_21_c10;
   bh1112_w44_34_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1498_Out0_c10(0);
   bh1112_w45_30_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1498_Out0_c10(1);
   bh1112_w46_27_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1498_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1498: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1498_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1498_Out0_copy1499_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1498_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1498_Out0_copy1499_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1500_In0_c9 <= "" & bh1112_w44_23_c9 & bh1112_w44_25_c9 & bh1112_w44_27_c9 & bh1112_w44_29_c9;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1500_In1_c10 <= "" & bh1112_w45_26_c10;
   bh1112_w44_35_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1500_Out0_c10(0);
   bh1112_w45_31_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1500_Out0_c10(1);
   bh1112_w46_28_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1500_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1500: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1500_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1500_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1500_Out0_copy1501_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1500_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1500_Out0_copy1501_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1502_In0_c10 <= "" & bh1112_w45_24_c10 & bh1112_w45_22_c10 & bh1112_w45_20_c10 & bh1112_w45_18_c10 & bh1112_w45_19_c10 & bh1112_w45_21_c10;
   bh1112_w45_32_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1502_Out0_c10(0);
   bh1112_w46_29_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1502_Out0_c10(1);
   bh1112_w47_24_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1502_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1502: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1502_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1502_Out0_copy1503_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1502_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1502_Out0_copy1503_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1504_In0_c10 <= "" & bh1112_w45_23_c10 & bh1112_w45_25_c10 & bh1112_w45_27_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1504_In1_c10 <= "" & bh1112_w46_26_c10 & bh1112_w46_24_c10;
   bh1112_w45_33_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1504_Out0_c10(0);
   bh1112_w46_30_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1504_Out0_c10(1);
   bh1112_w47_25_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1504_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1504: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1504_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1504_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1504_Out0_copy1505_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1504_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1504_Out0_copy1505_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1506_In0_c10 <= "" & bh1112_w46_22_c10 & bh1112_w46_20_c10 & bh1112_w46_18_c10 & bh1112_w46_19_c10 & bh1112_w46_21_c10 & bh1112_w46_23_c10;
   bh1112_w46_31_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1506_Out0_c10(0);
   bh1112_w47_26_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1506_Out0_c10(1);
   bh1112_w48_23_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1506_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1506: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1506_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1506_Out0_copy1507_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1506_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1506_Out0_copy1507_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1508_In0_c10 <= "" & bh1112_w47_22_c10 & bh1112_w47_20_c10 & bh1112_w47_18_c10 & bh1112_w47_16_c10 & bh1112_w47_15_c10 & bh1112_w47_17_c10;
   bh1112_w47_27_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1508_Out0_c10(0);
   bh1112_w48_24_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1508_Out0_c10(1);
   bh1112_w49_20_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1508_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1508: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1508_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1508_Out0_copy1509_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1508_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1508_Out0_copy1509_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1510_In0_c10 <= "" & bh1112_w47_19_c10 & bh1112_w47_21_c10 & bh1112_w47_23_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1510_In1_c10 <= "" & bh1112_w48_21_c10 & bh1112_w48_19_c10;
   bh1112_w47_28_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1510_Out0_c10(0);
   bh1112_w48_25_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1510_Out0_c10(1);
   bh1112_w49_21_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1510_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1510: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1510_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1510_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1510_Out0_copy1511_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1510_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1510_Out0_copy1511_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1512_In0_c10 <= "" & bh1112_w48_17_c10 & bh1112_w48_9_c10 & bh1112_w48_15_c10 & bh1112_w48_16_c10 & bh1112_w48_18_c10 & bh1112_w48_20_c10;
   bh1112_w48_26_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1512_Out0_c10(0);
   bh1112_w49_22_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1512_Out0_c10(1);
   bh1112_w50_18_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1512_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1512: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1512_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1512_Out0_copy1513_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1512_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1512_Out0_copy1513_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1514_In0_c10 <= "" & bh1112_w49_18_c10 & bh1112_w49_16_c10 & bh1112_w49_15_c10 & bh1112_w49_14_c10 & "0" & "0";
   bh1112_w49_23_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1514_Out0_c10(0);
   bh1112_w50_19_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1514_Out0_c10(1);
   bh1112_w51_15_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1514_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1514: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1514_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1514_Out0_copy1515_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1514_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1514_Out0_copy1515_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1516_In0_c10 <= "" & bh1112_w49_13_c10 & bh1112_w49_6_c10 & bh1112_w49_17_c10 & bh1112_w49_19_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1516_In1_c10 <= "" & bh1112_w50_17_c10;
   bh1112_w49_24_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1516_Out0_c10(0);
   bh1112_w50_20_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1516_Out0_c10(1);
   bh1112_w51_16_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1516_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1516: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1516_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1516_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1516_Out0_copy1517_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1516_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1516_Out0_copy1517_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1518_In0_c10 <= "" & bh1112_w50_11_c10 & bh1112_w50_12_c10 & bh1112_w50_13_c10 & bh1112_w50_14_c10 & bh1112_w50_15_c10 & bh1112_w50_16_c10;
   bh1112_w50_21_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1518_Out0_c10(0);
   bh1112_w51_17_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1518_Out0_c10(1);
   bh1112_w52_15_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1518_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1518: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1518_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1518_Out0_copy1519_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1518_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1518_Out0_copy1519_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1520_In0_c10 <= "" & bh1112_w51_9_c10 & bh1112_w51_10_c10 & bh1112_w51_11_c10 & bh1112_w51_12_c10 & bh1112_w51_13_c10 & bh1112_w51_14_c10;
   bh1112_w51_18_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1520_Out0_c10(0);
   bh1112_w52_16_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1520_Out0_c10(1);
   bh1112_w53_11_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1520_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1520: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1520_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1520_Out0_copy1521_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1520_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1520_Out0_copy1521_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1522_In0_c10 <= "" & bh1112_w52_9_c10 & bh1112_w52_10_c10 & bh1112_w52_11_c10 & bh1112_w52_12_c10 & bh1112_w52_13_c10 & bh1112_w52_14_c10;
   bh1112_w52_17_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1522_Out0_c10(0);
   bh1112_w53_12_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1522_Out0_c10(1);
   bh1112_w54_10_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1522_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1522: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1522_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1522_Out0_copy1523_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1522_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1522_Out0_copy1523_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1524_In0_c10 <= "" & bh1112_w53_6_c10 & bh1112_w53_7_c10 & bh1112_w53_8_c10 & bh1112_w53_9_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1524_In1_c9 <= "" & bh1112_w54_6_c9;
   bh1112_w53_13_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1524_Out0_c10(0);
   bh1112_w54_11_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1524_Out0_c10(1);
   bh1112_w55_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1524_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1524: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1524_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1524_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1524_Out0_copy1525_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1524_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1524_Out0_copy1525_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1526_In0_c10 <= "" & bh1112_w54_7_c10 & bh1112_w54_8_c10 & bh1112_w54_9_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1526_In1_c10 <= "" & bh1112_w55_6_c10 & bh1112_w55_7_c10;
   bh1112_w54_12_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1526_Out0_c10(0);
   bh1112_w55_10_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1526_Out0_c10(1);
   bh1112_w56_8_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1526_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1526: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1526_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1526_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1526_Out0_copy1527_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1526_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1526_Out0_copy1527_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In0_c10 <= "" & bh1112_w56_4_c10 & bh1112_w56_5_c10 & bh1112_w56_6_c10 & bh1112_w56_7_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c0 <= "" & "0";
   bh1112_w56_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1528_Out0_c10(0);
   bh1112_w57_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1528_Out0_c10(1);
   bh1112_w58_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1528_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1528: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1528_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1528_Out0_copy1529_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1528_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1528_Out0_copy1529_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1530_In0_c10 <= "" & bh1112_w57_4_c10 & bh1112_w57_5_c10 & bh1112_w57_6_c10;
   bh1112_w57_8_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1530_Out0_c10(0);
   bh1112_w58_8_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1530_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1530: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1530_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1530_Out0_copy1531_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1530_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1530_Out0_copy1531_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1532_In0_c10 <= "" & bh1112_w58_4_c10 & bh1112_w58_5_c10 & bh1112_w58_6_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1532_In1_c10 <= "" & bh1112_w59_3_c10 & bh1112_w59_4_c10;
   bh1112_w58_9_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1532_Out0_c10(0);
   bh1112_w59_5_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1532_Out0_c10(1);
   bh1112_w60_6_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1532_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1532: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1532_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1532_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1532_Out0_copy1533_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1532_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1532_Out0_copy1533_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1534_In0_c10 <= "" & bh1112_w60_3_c10 & bh1112_w60_4_c10 & bh1112_w60_5_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1534_In1_c10 <= "" & bh1112_w61_2_c10 & bh1112_w61_3_c10;
   bh1112_w60_7_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1534_Out0_c10(0);
   bh1112_w61_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1534_Out0_c10(1);
   bh1112_w62_5_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1534_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1534: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1534_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1534_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1534_Out0_copy1535_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1534_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1534_Out0_copy1535_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1536_In0_c10 <= "" & bh1112_w62_3_c10 & bh1112_w62_4_c10 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1536_In1_c10 <= "" & bh1112_w63_2_c10 & bh1112_w63_3_c10;
   bh1112_w62_6_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1536_Out0_c10(0);
   bh1112_w63_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1536_Out0_c10(1);
   bh1112_w64_5_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1536_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1536: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1536_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1536_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1536_Out0_copy1537_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1536_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1536_Out0_copy1537_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1538_In0_c10 <= "" & bh1112_w64_3_c10 & bh1112_w64_4_c10 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1538_In1_c10 <= "" & bh1112_w65_2_c10 & bh1112_w65_3_c10;
   bh1112_w64_6_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1538_Out0_c10(0);
   bh1112_w65_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1538_Out0_c10(1);
   bh1112_w66_5_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1538_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1538: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1538_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1538_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1538_Out0_copy1539_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1538_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1538_Out0_copy1539_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1540_In0_c10 <= "" & bh1112_w66_3_c10 & bh1112_w66_4_c10 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1540_In1_c10 <= "" & bh1112_w67_2_c10 & bh1112_w67_3_c10;
   bh1112_w66_6_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1540_Out0_c10(0);
   bh1112_w67_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1540_Out0_c10(1);
   bh1112_w68_5_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1540_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1540: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1540_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1540_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1540_Out0_copy1541_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1540_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1540_Out0_copy1541_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1542_In0_c10 <= "" & bh1112_w68_3_c10 & bh1112_w68_4_c10 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1542_In1_c10 <= "" & bh1112_w69_2_c10 & bh1112_w69_3_c10;
   bh1112_w68_6_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1542_Out0_c10(0);
   bh1112_w69_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1542_Out0_c10(1);
   bh1112_w70_4_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1542_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1542: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1542_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1542_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1542_Out0_copy1543_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1542_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1542_Out0_copy1543_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1544_In0_c10 <= "" & bh1112_w70_2_c10 & bh1112_w70_3_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1544_In1_c10 <= "" & bh1112_w71_2_c10;
   bh1112_w70_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1544_Out0_c10(0);
   bh1112_w71_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1544_Out0_c10(1);
   bh1112_w72_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1544_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1544: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1544_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1544_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1544_Out0_copy1545_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1544_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1544_Out0_copy1545_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1546_In0_c10 <= "" & bh1112_w72_2_c10 & bh1112_w72_3_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1546_In1_c10 <= "" & bh1112_w73_2_c10;
   bh1112_w72_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1546_Out0_c10(0);
   bh1112_w73_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1546_Out0_c10(1);
   bh1112_w74_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1546_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1546: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1546_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1546_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1546_Out0_copy1547_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1546_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1546_Out0_copy1547_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1548_In0_c10 <= "" & bh1112_w74_2_c10 & bh1112_w74_3_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1548_In1_c10 <= "" & bh1112_w75_2_c10;
   bh1112_w74_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1548_Out0_c10(0);
   bh1112_w75_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1548_Out0_c10(1);
   bh1112_w76_2_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1548_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1548: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1548_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1548_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1548_Out0_copy1549_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1548_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1548_Out0_copy1549_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1550_In0_c10 <= "" & bh1112_w76_0_c10 & bh1112_w76_1_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1550_In1_c9 <= "" & bh1112_w77_0_c9;
   bh1112_w76_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1550_Out0_c10(0);
   bh1112_w77_1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1550_Out0_c10(1);
   bh1112_w78_1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1550_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1550: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1550_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1550_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1550_Out0_copy1551_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1550_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1550_Out0_copy1551_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1552_In0_c10 <= "" & bh1112_w38_4_c10 & "0" & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1552_In1_c10 <= "" & bh1112_w39_34_c10 & bh1112_w39_35_c10;
   bh1112_w38_5_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1552_Out0_c10(0);
   bh1112_w39_36_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1552_Out0_c10(1);
   bh1112_w40_30_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1552_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1552: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1552_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1552_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1552_Out0_copy1553_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1552_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1552_Out0_copy1553_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1554_In0_c10 <= "" & bh1112_w40_27_c10 & bh1112_w40_28_c10 & bh1112_w40_29_c10;
   bh1112_w40_31_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1554_Out0_c10(0);
   bh1112_w41_34_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1554_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1554: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1554_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1554_Out0_copy1555_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1554_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1554_Out0_copy1555_c10; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid1557_bh1112_uid1558_In0_c10 <= "" & bh1112_w41_29_c10 & bh1112_w41_30_c10 & bh1112_w41_31_c10 & bh1112_w41_32_c10 & bh1112_w41_33_c10;
   bh1112_w41_35_c10 <= Compressor_5_3_Freq300_uid1557_bh1112_uid1558_Out0_c10(0);
   bh1112_w42_38_c10 <= Compressor_5_3_Freq300_uid1557_bh1112_uid1558_Out0_c10(1);
   bh1112_w43_38_c10 <= Compressor_5_3_Freq300_uid1557_bh1112_uid1558_Out0_c10(2);
   Compressor_5_3_Freq300_uid1557_uid1558: Compressor_5_3_Freq300_uid1557
      port map ( X0 => Compressor_5_3_Freq300_uid1557_bh1112_uid1558_In0_c10,
                 R => Compressor_5_3_Freq300_uid1557_bh1112_uid1558_Out0_copy1559_c10);
   Compressor_5_3_Freq300_uid1557_bh1112_uid1558_Out0_c10 <= Compressor_5_3_Freq300_uid1557_bh1112_uid1558_Out0_copy1559_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1560_In0_c10 <= "" & bh1112_w42_32_c10 & bh1112_w42_33_c10 & bh1112_w42_34_c10 & bh1112_w42_35_c10 & bh1112_w42_36_c10 & bh1112_w42_37_c10;
   bh1112_w42_39_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1560_Out0_c10(0);
   bh1112_w43_39_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1560_Out0_c10(1);
   bh1112_w44_36_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1560_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1560: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1560_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1560_Out0_copy1561_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1560_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1560_Out0_copy1561_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1562_In0_c10 <= "" & bh1112_w43_31_c10 & bh1112_w43_32_c10 & bh1112_w43_33_c10 & bh1112_w43_34_c10 & bh1112_w43_35_c10 & bh1112_w43_36_c10;
   bh1112_w43_40_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1562_Out0_c10(0);
   bh1112_w44_37_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1562_Out0_c10(1);
   bh1112_w45_34_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1562_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1562: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1562_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1562_Out0_copy1563_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1562_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1562_Out0_copy1563_c10; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid1557_bh1112_uid1564_In0_c10 <= "" & bh1112_w44_31_c10 & bh1112_w44_32_c10 & bh1112_w44_33_c10 & bh1112_w44_34_c10 & bh1112_w44_35_c10;
   bh1112_w44_38_c10 <= Compressor_5_3_Freq300_uid1557_bh1112_uid1564_Out0_c10(0);
   bh1112_w45_35_c10 <= Compressor_5_3_Freq300_uid1557_bh1112_uid1564_Out0_c10(1);
   bh1112_w46_32_c10 <= Compressor_5_3_Freq300_uid1557_bh1112_uid1564_Out0_c10(2);
   Compressor_5_3_Freq300_uid1557_uid1564: Compressor_5_3_Freq300_uid1557
      port map ( X0 => Compressor_5_3_Freq300_uid1557_bh1112_uid1564_In0_c10,
                 R => Compressor_5_3_Freq300_uid1557_bh1112_uid1564_Out0_copy1565_c10);
   Compressor_5_3_Freq300_uid1557_bh1112_uid1564_Out0_c10 <= Compressor_5_3_Freq300_uid1557_bh1112_uid1564_Out0_copy1565_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1566_In0_c10 <= "" & bh1112_w45_28_c10 & bh1112_w45_29_c10 & bh1112_w45_30_c10 & bh1112_w45_31_c10 & bh1112_w45_32_c10 & bh1112_w45_33_c10;
   bh1112_w45_36_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1566_Out0_c10(0);
   bh1112_w46_33_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1566_Out0_c10(1);
   bh1112_w47_29_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1566_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1566: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1566_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1566_Out0_copy1567_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1566_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1566_Out0_copy1567_c10; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid1363_bh1112_uid1568_In0_c10 <= "" & bh1112_w46_25_c10 & bh1112_w46_27_c10 & bh1112_w46_28_c10 & bh1112_w46_29_c10 & bh1112_w46_30_c10 & bh1112_w46_31_c10;
   bh1112_w46_34_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1568_Out0_c10(0);
   bh1112_w47_30_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1568_Out0_c10(1);
   bh1112_w48_27_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1568_Out0_c10(2);
   Compressor_6_3_Freq300_uid1363_uid1568: Compressor_6_3_Freq300_uid1363
      port map ( X0 => Compressor_6_3_Freq300_uid1363_bh1112_uid1568_In0_c10,
                 R => Compressor_6_3_Freq300_uid1363_bh1112_uid1568_Out0_copy1569_c10);
   Compressor_6_3_Freq300_uid1363_bh1112_uid1568_Out0_c10 <= Compressor_6_3_Freq300_uid1363_bh1112_uid1568_Out0_copy1569_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1570_In0_c10 <= "" & bh1112_w47_24_c10 & bh1112_w47_25_c10 & bh1112_w47_26_c10 & bh1112_w47_27_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1570_In1_c10 <= "" & bh1112_w48_22_c10;
   bh1112_w47_31_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1570_Out0_c10(0);
   bh1112_w48_28_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1570_Out0_c10(1);
   bh1112_w49_25_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1570_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1570: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1570_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1570_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1570_Out0_copy1571_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1570_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1570_Out0_copy1571_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1572_In0_c10 <= "" & bh1112_w48_23_c10 & bh1112_w48_24_c10 & bh1112_w48_25_c10 & bh1112_w48_26_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1572_In1_c10 <= "" & bh1112_w49_20_c10;
   bh1112_w48_29_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1572_Out0_c10(0);
   bh1112_w49_26_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1572_Out0_c10(1);
   bh1112_w50_22_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1572_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1572: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1572_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1572_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1572_Out0_copy1573_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1572_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1572_Out0_copy1573_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1574_In0_c10 <= "" & bh1112_w49_21_c10 & bh1112_w49_22_c10 & bh1112_w49_23_c10 & bh1112_w49_24_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1574_In1_c10 <= "" & bh1112_w50_18_c10;
   bh1112_w49_27_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1574_Out0_c10(0);
   bh1112_w50_23_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1574_Out0_c10(1);
   bh1112_w51_19_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1574_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1574: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1574_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1574_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1574_Out0_copy1575_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1574_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1574_Out0_copy1575_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1576_In0_c10 <= "" & bh1112_w50_19_c10 & bh1112_w50_20_c10 & bh1112_w50_21_c10;
   bh1112_w50_24_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1576_Out0_c10(0);
   bh1112_w51_20_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1576_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1576: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1576_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1576_Out0_copy1577_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1576_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1576_Out0_copy1577_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In0_c10 <= "" & bh1112_w51_15_c10 & bh1112_w51_16_c10 & bh1112_w51_17_c10 & bh1112_w51_18_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c0 <= "" & "0";
   bh1112_w51_21_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1578_Out0_c10(0);
   bh1112_w52_18_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1578_Out0_c10(1);
   bh1112_w53_14_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1578_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1578: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1578_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1578_Out0_copy1579_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1578_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1578_Out0_copy1579_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1580_In0_c10 <= "" & bh1112_w52_15_c10 & bh1112_w52_16_c10 & bh1112_w52_17_c10;
   bh1112_w52_19_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1580_Out0_c10(0);
   bh1112_w53_15_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1580_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1580: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1580_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1580_Out0_copy1581_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1580_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1580_Out0_copy1581_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In0_c10 <= "" & bh1112_w53_10_c10 & bh1112_w53_11_c10 & bh1112_w53_12_c10 & bh1112_w53_13_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c0 <= "" & "0";
   bh1112_w53_16_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1582_Out0_c10(0);
   bh1112_w54_13_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1582_Out0_c10(1);
   bh1112_w55_11_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1582_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1582: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1582_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1582_Out0_copy1583_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1582_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1582_Out0_copy1583_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1584_In0_c10 <= "" & bh1112_w54_10_c10 & bh1112_w54_11_c10 & bh1112_w54_12_c10;
   bh1112_w54_14_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1584_Out0_c10(0);
   bh1112_w55_12_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1584_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1584: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1584_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1584_Out0_copy1585_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1584_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1584_Out0_copy1585_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1586_In0_c10 <= "" & bh1112_w55_8_c10 & bh1112_w55_9_c10 & bh1112_w55_10_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1586_In1_c10 <= "" & bh1112_w56_8_c10 & bh1112_w56_9_c10;
   bh1112_w55_13_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1586_Out0_c10(0);
   bh1112_w56_10_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1586_Out0_c10(1);
   bh1112_w57_9_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1586_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1586: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1586_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1586_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1586_Out0_copy1587_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1586_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1586_Out0_copy1587_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1588_In0_c10 <= "" & bh1112_w57_7_c10 & bh1112_w57_8_c10 & "0";
   bh1112_w57_10_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1588_Out0_c10(0);
   bh1112_w58_10_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1588_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1588: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1588_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1588_Out0_copy1589_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1588_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1588_Out0_copy1589_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1590_In0_c10 <= "" & bh1112_w58_7_c10 & bh1112_w58_8_c10 & bh1112_w58_9_c10;
   bh1112_w58_11_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1590_Out0_c10(0);
   bh1112_w59_6_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1590_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1590: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1590_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1590_Out0_copy1591_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1590_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1590_Out0_copy1591_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1592_In0_c10 <= "" & bh1112_w60_6_c10 & bh1112_w60_7_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1592_In1_c10 <= "" & bh1112_w61_4_c10;
   bh1112_w60_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1592_Out0_c10(0);
   bh1112_w61_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1592_Out0_c10(1);
   bh1112_w62_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1592_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1592: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1592_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1592_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1592_Out0_copy1593_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1592_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1592_Out0_copy1593_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1594_In0_c10 <= "" & bh1112_w62_5_c10 & bh1112_w62_6_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1594_In1_c10 <= "" & bh1112_w63_4_c10;
   bh1112_w62_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1594_Out0_c10(0);
   bh1112_w63_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1594_Out0_c10(1);
   bh1112_w64_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1594_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1594: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1594_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1594_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1594_Out0_copy1595_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1594_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1594_Out0_copy1595_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1596_In0_c10 <= "" & bh1112_w64_5_c10 & bh1112_w64_6_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1596_In1_c10 <= "" & bh1112_w65_4_c10;
   bh1112_w64_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1596_Out0_c10(0);
   bh1112_w65_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1596_Out0_c10(1);
   bh1112_w66_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1596_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1596: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1596_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1596_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1596_Out0_copy1597_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1596_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1596_Out0_copy1597_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1598_In0_c10 <= "" & bh1112_w66_5_c10 & bh1112_w66_6_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1598_In1_c10 <= "" & bh1112_w67_4_c10;
   bh1112_w66_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1598_Out0_c10(0);
   bh1112_w67_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1598_Out0_c10(1);
   bh1112_w68_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1598_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1598: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1598_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1598_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1598_Out0_copy1599_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1598_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1598_Out0_copy1599_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1600_In0_c10 <= "" & bh1112_w68_5_c10 & bh1112_w68_6_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1600_In1_c10 <= "" & bh1112_w69_4_c10;
   bh1112_w68_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1600_Out0_c10(0);
   bh1112_w69_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1600_Out0_c10(1);
   bh1112_w70_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1600_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1600: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1600_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1600_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1600_Out0_copy1601_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1600_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1600_Out0_copy1601_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1602_In0_c10 <= "" & bh1112_w70_4_c10 & bh1112_w70_5_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1602_In1_c10 <= "" & bh1112_w71_3_c10;
   bh1112_w70_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1602_Out0_c10(0);
   bh1112_w71_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1602_Out0_c10(1);
   bh1112_w72_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1602_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1602: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1602_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1602_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1602_Out0_copy1603_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1602_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1602_Out0_copy1603_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1604_In0_c10 <= "" & bh1112_w72_4_c10 & bh1112_w72_5_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1604_In1_c10 <= "" & bh1112_w73_3_c10;
   bh1112_w72_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1604_Out0_c10(0);
   bh1112_w73_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1604_Out0_c10(1);
   bh1112_w74_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1604_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1604: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1604_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1604_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1604_Out0_copy1605_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1604_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1604_Out0_copy1605_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1606_In0_c10 <= "" & bh1112_w74_4_c10 & bh1112_w74_5_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1606_In1_c10 <= "" & bh1112_w75_3_c10;
   bh1112_w74_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1606_Out0_c10(0);
   bh1112_w75_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1606_Out0_c10(1);
   bh1112_w76_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1606_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1606: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1606_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1606_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1606_Out0_copy1607_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1606_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1606_Out0_copy1607_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1608_In0_c10 <= "" & bh1112_w76_2_c10 & bh1112_w76_3_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1608_In1_c10 <= "" & bh1112_w77_1_c10;
   bh1112_w76_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1608_Out0_c10(0);
   bh1112_w77_2_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1608_Out0_c10(1);
   bh1112_w78_2_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1608_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1608: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1608_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1608_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1608_Out0_copy1609_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1608_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1608_Out0_copy1609_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1610_In0_c10 <= "" & bh1112_w78_0_c10 & bh1112_w78_1_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1610_In1_c9 <= "" & bh1112_w79_0_c9;
   bh1112_w78_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1610_Out0_c10(0);
   bh1112_w79_1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1610_Out0_c10(1);
   bh1112_w80_1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1610_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1610: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1610_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1610_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1610_Out0_copy1611_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1610_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1610_Out0_copy1611_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1612_In0_c10 <= "" & bh1112_w40_30_c10 & bh1112_w40_31_c10 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1612_In1_c10 <= "" & bh1112_w41_34_c10 & bh1112_w41_35_c10;
   bh1112_w40_32_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1612_Out0_c10(0);
   bh1112_w41_36_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1612_Out0_c10(1);
   bh1112_w42_40_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1612_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1612: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1612_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1612_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1612_Out0_copy1613_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1612_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1612_Out0_copy1613_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1614_In0_c10 <= "" & bh1112_w42_38_c10 & bh1112_w42_39_c10 & "0";
   bh1112_w42_41_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1614_Out0_c10(0);
   bh1112_w43_41_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1614_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1614: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1614_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1614_Out0_copy1615_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1614_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1614_Out0_copy1615_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In0_c10 <= "" & bh1112_w43_37_c10 & bh1112_w43_38_c10 & bh1112_w43_39_c10 & bh1112_w43_40_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c0 <= "" & "0";
   bh1112_w43_42_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1616_Out0_c10(0);
   bh1112_w44_39_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1616_Out0_c10(1);
   bh1112_w45_37_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1616_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1616: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1616_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1616_Out0_copy1617_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1616_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1616_Out0_copy1617_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1618_In0_c10 <= "" & bh1112_w44_36_c10 & bh1112_w44_37_c10 & bh1112_w44_38_c10;
   bh1112_w44_40_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1618_Out0_c10(0);
   bh1112_w45_38_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1618_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1618: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1618_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1618_Out0_copy1619_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1618_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1618_Out0_copy1619_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1620_In0_c10 <= "" & bh1112_w45_34_c10 & bh1112_w45_35_c10 & bh1112_w45_36_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1620_In1_c10 <= "" & bh1112_w46_32_c10 & bh1112_w46_33_c10;
   bh1112_w45_39_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1620_Out0_c10(0);
   bh1112_w46_35_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1620_Out0_c10(1);
   bh1112_w47_32_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1620_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1620: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1620_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1620_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1620_Out0_copy1621_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1620_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1620_Out0_copy1621_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In0_c10 <= "" & bh1112_w47_28_c10 & bh1112_w47_29_c10 & bh1112_w47_30_c10 & bh1112_w47_31_c10;
   Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c0 <= "" & "0";
   bh1112_w47_33_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1622_Out0_c10(0);
   bh1112_w48_30_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1622_Out0_c10(1);
   bh1112_w49_28_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1622_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1622: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1622_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1622_Out0_copy1623_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1622_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1622_Out0_copy1623_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1624_In0_c10 <= "" & bh1112_w48_27_c10 & bh1112_w48_28_c10 & bh1112_w48_29_c10;
   bh1112_w48_31_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1624_Out0_c10(0);
   bh1112_w49_29_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1624_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1624: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1624_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1624_Out0_copy1625_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1624_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1624_Out0_copy1625_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1626_In0_c10 <= "" & bh1112_w49_25_c10 & bh1112_w49_26_c10 & bh1112_w49_27_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1626_In1_c10 <= "" & bh1112_w50_22_c10 & bh1112_w50_23_c10;
   bh1112_w49_30_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1626_Out0_c10(0);
   bh1112_w50_25_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1626_Out0_c10(1);
   bh1112_w51_22_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1626_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1626: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1626_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1626_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1626_Out0_copy1627_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1626_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1626_Out0_copy1627_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1628_In0_c10 <= "" & bh1112_w51_19_c10 & bh1112_w51_20_c10 & bh1112_w51_21_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1628_In1_c10 <= "" & bh1112_w52_18_c10 & bh1112_w52_19_c10;
   bh1112_w51_23_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1628_Out0_c10(0);
   bh1112_w52_20_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1628_Out0_c10(1);
   bh1112_w53_17_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1628_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1628: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1628_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1628_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1628_Out0_copy1629_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1628_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1628_Out0_copy1629_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1630_In0_c10 <= "" & bh1112_w53_14_c10 & bh1112_w53_15_c10 & bh1112_w53_16_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1630_In1_c10 <= "" & bh1112_w54_13_c10 & bh1112_w54_14_c10;
   bh1112_w53_18_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1630_Out0_c10(0);
   bh1112_w54_15_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1630_Out0_c10(1);
   bh1112_w55_14_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1630_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1630: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1630_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1630_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1630_Out0_copy1631_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1630_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1630_Out0_copy1631_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1632_In0_c10 <= "" & bh1112_w55_11_c10 & bh1112_w55_12_c10 & bh1112_w55_13_c10;
   bh1112_w55_15_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1632_Out0_c10(0);
   bh1112_w56_11_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1632_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1632: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1632_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1632_Out0_copy1633_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1632_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1632_Out0_copy1633_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1634_In0_c10 <= "" & bh1112_w57_9_c10 & bh1112_w57_10_c10 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1634_In1_c10 <= "" & bh1112_w58_10_c10 & bh1112_w58_11_c10;
   bh1112_w57_11_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1634_Out0_c10(0);
   bh1112_w58_12_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1634_Out0_c10(1);
   bh1112_w59_7_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1634_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1634: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1634_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1634_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1634_Out0_copy1635_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1634_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1634_Out0_copy1635_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1636_In0_c10 <= "" & bh1112_w59_5_c10 & bh1112_w59_6_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1636_In1_c10 <= "" & bh1112_w60_8_c10;
   bh1112_w59_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1636_Out0_c10(0);
   bh1112_w60_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1636_Out0_c10(1);
   bh1112_w61_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1636_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1636: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1636_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1636_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1636_Out0_copy1637_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1636_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1636_Out0_copy1637_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1638_In0_c10 <= "" & bh1112_w62_7_c10 & bh1112_w62_8_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1638_In1_c10 <= "" & bh1112_w63_5_c10;
   bh1112_w62_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1638_Out0_c10(0);
   bh1112_w63_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1638_Out0_c10(1);
   bh1112_w64_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1638_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1638: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1638_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1638_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1638_Out0_copy1639_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1638_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1638_Out0_copy1639_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1640_In0_c10 <= "" & bh1112_w64_7_c10 & bh1112_w64_8_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1640_In1_c10 <= "" & bh1112_w65_5_c10;
   bh1112_w64_10_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1640_Out0_c10(0);
   bh1112_w65_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1640_Out0_c10(1);
   bh1112_w66_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1640_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1640: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1640_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1640_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1640_Out0_copy1641_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1640_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1640_Out0_copy1641_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1642_In0_c10 <= "" & bh1112_w66_7_c10 & bh1112_w66_8_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1642_In1_c10 <= "" & bh1112_w67_5_c10;
   bh1112_w66_10_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1642_Out0_c10(0);
   bh1112_w67_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1642_Out0_c10(1);
   bh1112_w68_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1642_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1642: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1642_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1642_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1642_Out0_copy1643_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1642_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1642_Out0_copy1643_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1644_In0_c10 <= "" & bh1112_w68_7_c10 & bh1112_w68_8_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1644_In1_c10 <= "" & bh1112_w69_5_c10;
   bh1112_w68_10_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1644_Out0_c10(0);
   bh1112_w69_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1644_Out0_c10(1);
   bh1112_w70_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1644_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1644: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1644_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1644_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1644_Out0_copy1645_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1644_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1644_Out0_copy1645_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1646_In0_c10 <= "" & bh1112_w70_6_c10 & bh1112_w70_7_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1646_In1_c10 <= "" & bh1112_w71_4_c10;
   bh1112_w70_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1646_Out0_c10(0);
   bh1112_w71_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1646_Out0_c10(1);
   bh1112_w72_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1646_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1646: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1646_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1646_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1646_Out0_copy1647_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1646_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1646_Out0_copy1647_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1648_In0_c10 <= "" & bh1112_w72_6_c10 & bh1112_w72_7_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1648_In1_c10 <= "" & bh1112_w73_4_c10;
   bh1112_w72_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1648_Out0_c10(0);
   bh1112_w73_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1648_Out0_c10(1);
   bh1112_w74_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1648_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1648: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1648_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1648_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1648_Out0_copy1649_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1648_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1648_Out0_copy1649_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1650_In0_c10 <= "" & bh1112_w74_6_c10 & bh1112_w74_7_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1650_In1_c10 <= "" & bh1112_w75_4_c10;
   bh1112_w74_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1650_Out0_c10(0);
   bh1112_w75_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1650_Out0_c10(1);
   bh1112_w76_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1650_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1650: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1650_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1650_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1650_Out0_copy1651_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1650_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1650_Out0_copy1651_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1652_In0_c10 <= "" & bh1112_w76_4_c10 & bh1112_w76_5_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1652_In1_c10 <= "" & bh1112_w77_2_c10;
   bh1112_w76_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1652_Out0_c10(0);
   bh1112_w77_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1652_Out0_c10(1);
   bh1112_w78_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1652_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1652: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1652_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1652_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1652_Out0_copy1653_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1652_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1652_Out0_copy1653_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1654_In0_c10 <= "" & bh1112_w78_2_c10 & bh1112_w78_3_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1654_In1_c10 <= "" & bh1112_w79_1_c10;
   bh1112_w78_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1654_Out0_c10(0);
   bh1112_w79_2_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1654_Out0_c10(1);
   bh1112_w80_2_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1654_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1654: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1654_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1654_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1654_Out0_copy1655_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1654_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1654_Out0_copy1655_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1656_In0_c10 <= "" & bh1112_w80_0_c10 & bh1112_w80_1_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1656_In1_c9 <= "" & bh1112_w81_0_c9;
   bh1112_w80_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1656_Out0_c10(0);
   bh1112_w81_1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1656_Out0_c10(1);
   bh1112_w82_1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1656_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1656: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1656_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1656_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1656_Out0_copy1657_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1656_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1656_Out0_copy1657_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1658_In0_c10 <= "" & bh1112_w42_40_c10 & bh1112_w42_41_c10 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1658_In1_c10 <= "" & bh1112_w43_41_c10 & bh1112_w43_42_c10;
   bh1112_w42_42_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1658_Out0_c10(0);
   bh1112_w43_43_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1658_Out0_c10(1);
   bh1112_w44_41_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1658_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1658: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1658_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1658_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1658_Out0_copy1659_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1658_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1658_Out0_copy1659_c10; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid1359_bh1112_uid1660_In0_c10 <= "" & bh1112_w44_39_c10 & bh1112_w44_40_c10 & "0";
   bh1112_w44_42_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1660_Out0_c10(0);
   bh1112_w45_40_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1660_Out0_c10(1);
   Compressor_3_2_Freq300_uid1359_uid1660: Compressor_3_2_Freq300_uid1359
      port map ( X0 => Compressor_3_2_Freq300_uid1359_bh1112_uid1660_In0_c10,
                 R => Compressor_3_2_Freq300_uid1359_bh1112_uid1660_Out0_copy1661_c10);
   Compressor_3_2_Freq300_uid1359_bh1112_uid1660_Out0_c10 <= Compressor_3_2_Freq300_uid1359_bh1112_uid1660_Out0_copy1661_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1662_In0_c10 <= "" & bh1112_w45_37_c10 & bh1112_w45_38_c10 & bh1112_w45_39_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1662_In1_c10 <= "" & bh1112_w46_34_c10 & bh1112_w46_35_c10;
   bh1112_w45_41_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1662_Out0_c10(0);
   bh1112_w46_36_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1662_Out0_c10(1);
   bh1112_w47_34_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1662_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1662: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1662_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1662_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1662_Out0_copy1663_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1662_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1662_Out0_copy1663_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1664_In0_c10 <= "" & bh1112_w47_32_c10 & bh1112_w47_33_c10 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1664_In1_c10 <= "" & bh1112_w48_30_c10 & bh1112_w48_31_c10;
   bh1112_w47_35_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1664_Out0_c10(0);
   bh1112_w48_32_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1664_Out0_c10(1);
   bh1112_w49_31_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1664_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1664: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1664_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1664_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1664_Out0_copy1665_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1664_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1664_Out0_copy1665_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1666_In0_c10 <= "" & bh1112_w49_28_c10 & bh1112_w49_29_c10 & bh1112_w49_30_c10;
   Compressor_23_3_Freq300_uid1355_bh1112_uid1666_In1_c10 <= "" & bh1112_w50_24_c10 & bh1112_w50_25_c10;
   bh1112_w49_32_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1666_Out0_c10(0);
   bh1112_w50_26_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1666_Out0_c10(1);
   bh1112_w51_24_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1666_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1666: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1666_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1666_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1666_Out0_copy1667_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1666_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1666_Out0_copy1667_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1668_In0_c10 <= "" & bh1112_w51_22_c10 & bh1112_w51_23_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1668_In1_c10 <= "" & bh1112_w52_20_c10;
   bh1112_w51_25_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1668_Out0_c10(0);
   bh1112_w52_21_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1668_Out0_c10(1);
   bh1112_w53_19_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1668_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1668: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1668_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1668_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1668_Out0_copy1669_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1668_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1668_Out0_copy1669_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1670_In0_c10 <= "" & bh1112_w53_17_c10 & bh1112_w53_18_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1670_In1_c10 <= "" & bh1112_w54_15_c10;
   bh1112_w53_20_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1670_Out0_c10(0);
   bh1112_w54_16_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1670_Out0_c10(1);
   bh1112_w55_16_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1670_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1670: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1670_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1670_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1670_Out0_copy1671_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1670_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1670_Out0_copy1671_c10; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid1355_bh1112_uid1672_In0_c10 <= "" & bh1112_w55_14_c10 & bh1112_w55_15_c10 & "0";
   Compressor_23_3_Freq300_uid1355_bh1112_uid1672_In1_c10 <= "" & bh1112_w56_10_c10 & bh1112_w56_11_c10;
   bh1112_w55_17_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1672_Out0_c10(0);
   bh1112_w56_12_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1672_Out0_c10(1);
   bh1112_w57_12_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1672_Out0_c10(2);
   Compressor_23_3_Freq300_uid1355_uid1672: Compressor_23_3_Freq300_uid1355
      port map ( X0 => Compressor_23_3_Freq300_uid1355_bh1112_uid1672_In0_c10,
                 X1 => Compressor_23_3_Freq300_uid1355_bh1112_uid1672_In1_c10,
                 R => Compressor_23_3_Freq300_uid1355_bh1112_uid1672_Out0_copy1673_c10);
   Compressor_23_3_Freq300_uid1355_bh1112_uid1672_Out0_c10 <= Compressor_23_3_Freq300_uid1355_bh1112_uid1672_Out0_copy1673_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1674_In0_c10 <= "" & bh1112_w59_7_c10 & bh1112_w59_8_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1674_In1_c10 <= "" & bh1112_w60_9_c10;
   bh1112_w59_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1674_Out0_c10(0);
   bh1112_w60_10_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1674_Out0_c10(1);
   bh1112_w61_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1674_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1674: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1674_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1674_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1674_Out0_copy1675_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1674_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1674_Out0_copy1675_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1676_In0_c10 <= "" & bh1112_w61_5_c10 & bh1112_w61_6_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1676_In1_c10 <= "" & bh1112_w62_9_c10;
   bh1112_w61_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1676_Out0_c10(0);
   bh1112_w62_10_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1676_Out0_c10(1);
   bh1112_w63_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1676_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1676: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1676_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1676_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1676_Out0_copy1677_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1676_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1676_Out0_copy1677_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1678_In0_c10 <= "" & bh1112_w64_9_c10 & bh1112_w64_10_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1678_In1_c10 <= "" & bh1112_w65_6_c10;
   bh1112_w64_11_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1678_Out0_c10(0);
   bh1112_w65_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1678_Out0_c10(1);
   bh1112_w66_11_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1678_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1678: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1678_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1678_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1678_Out0_copy1679_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1678_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1678_Out0_copy1679_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1680_In0_c10 <= "" & bh1112_w66_9_c10 & bh1112_w66_10_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1680_In1_c10 <= "" & bh1112_w67_6_c10;
   bh1112_w66_12_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1680_Out0_c10(0);
   bh1112_w67_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1680_Out0_c10(1);
   bh1112_w68_11_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1680_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1680: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1680_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1680_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1680_Out0_copy1681_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1680_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1680_Out0_copy1681_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1682_In0_c10 <= "" & bh1112_w68_9_c10 & bh1112_w68_10_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1682_In1_c10 <= "" & bh1112_w69_6_c10;
   bh1112_w68_12_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1682_Out0_c10(0);
   bh1112_w69_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1682_Out0_c10(1);
   bh1112_w70_10_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1682_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1682: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1682_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1682_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1682_Out0_copy1683_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1682_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1682_Out0_copy1683_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1684_In0_c10 <= "" & bh1112_w70_8_c10 & bh1112_w70_9_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1684_In1_c10 <= "" & bh1112_w71_5_c10;
   bh1112_w70_11_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1684_Out0_c10(0);
   bh1112_w71_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1684_Out0_c10(1);
   bh1112_w72_10_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1684_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1684: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1684_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1684_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1684_Out0_copy1685_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1684_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1684_Out0_copy1685_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1686_In0_c10 <= "" & bh1112_w72_8_c10 & bh1112_w72_9_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1686_In1_c10 <= "" & bh1112_w73_5_c10;
   bh1112_w72_11_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1686_Out0_c10(0);
   bh1112_w73_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1686_Out0_c10(1);
   bh1112_w74_10_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1686_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1686: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1686_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1686_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1686_Out0_copy1687_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1686_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1686_Out0_copy1687_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1688_In0_c10 <= "" & bh1112_w74_8_c10 & bh1112_w74_9_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1688_In1_c10 <= "" & bh1112_w75_5_c10;
   bh1112_w74_11_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1688_Out0_c10(0);
   bh1112_w75_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1688_Out0_c10(1);
   bh1112_w76_8_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1688_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1688: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1688_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1688_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1688_Out0_copy1689_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1688_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1688_Out0_copy1689_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1690_In0_c10 <= "" & bh1112_w76_6_c10 & bh1112_w76_7_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1690_In1_c10 <= "" & bh1112_w77_3_c10;
   bh1112_w76_9_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1690_Out0_c10(0);
   bh1112_w77_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1690_Out0_c10(1);
   bh1112_w78_6_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1690_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1690: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1690_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1690_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1690_Out0_copy1691_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1690_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1690_Out0_copy1691_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1692_In0_c10 <= "" & bh1112_w78_4_c10 & bh1112_w78_5_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1692_In1_c10 <= "" & bh1112_w79_2_c10;
   bh1112_w78_7_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1692_Out0_c10(0);
   bh1112_w79_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1692_Out0_c10(1);
   bh1112_w80_4_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1692_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1692: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1692_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1692_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1692_Out0_copy1693_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1692_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1692_Out0_copy1693_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1694_In0_c10 <= "" & bh1112_w80_2_c10 & bh1112_w80_3_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1694_In1_c10 <= "" & bh1112_w81_1_c10;
   bh1112_w80_5_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1694_Out0_c10(0);
   bh1112_w81_2_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1694_Out0_c10(1);
   bh1112_w82_2_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1694_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1694: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1694_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1694_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1694_Out0_copy1695_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1694_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1694_Out0_copy1695_c10; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid1373_bh1112_uid1696_In0_c10 <= "" & bh1112_w82_0_c10 & bh1112_w82_1_c10 & "0" & "0";
   Compressor_14_3_Freq300_uid1373_bh1112_uid1696_In1_c9 <= "" & bh1112_w83_0_c9;
   bh1112_w82_3_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1696_Out0_c10(0);
   bh1112_w83_1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1696_Out0_c10(1);
   bh1112_w84_1_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1696_Out0_c10(2);
   Compressor_14_3_Freq300_uid1373_uid1696: Compressor_14_3_Freq300_uid1373
      port map ( X0 => Compressor_14_3_Freq300_uid1373_bh1112_uid1696_In0_c10,
                 X1 => Compressor_14_3_Freq300_uid1373_bh1112_uid1696_In1_c10,
                 R => Compressor_14_3_Freq300_uid1373_bh1112_uid1696_Out0_copy1697_c10);
   Compressor_14_3_Freq300_uid1373_bh1112_uid1696_Out0_c10 <= Compressor_14_3_Freq300_uid1373_bh1112_uid1696_Out0_copy1697_c10; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh1112_43_c10 <= bh1112_w43_43_c10 & bh1112_w42_42_c10 & bh1112_w41_36_c10 & bh1112_w40_32_c10 & bh1112_w39_36_c10 & bh1112_w38_5_c10 & bh1112_w37_3_c10 & bh1112_w36_2_c10 & bh1112_w35_0_c10 & bh1112_w34_0_c10 & bh1112_w33_0_c10 & bh1112_w32_0_c10 & bh1112_w31_0_c10 & bh1112_w30_0_c10 & bh1112_w29_0_c10 & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0";

   bitheapFinalAdd_bh1112_In0_c10 <= "0" & bh1112_w92_0_c10 & bh1112_w91_0_c10 & bh1112_w90_0_c10 & bh1112_w89_0_c10 & bh1112_w88_0_c10 & bh1112_w87_0_c10 & bh1112_w86_0_c10 & bh1112_w85_0_c10 & bh1112_w84_0_c10 & bh1112_w83_1_c10 & bh1112_w82_2_c10 & bh1112_w81_2_c10 & bh1112_w80_4_c10 & bh1112_w79_3_c10 & bh1112_w78_6_c10 & bh1112_w77_4_c10 & bh1112_w76_8_c10 & bh1112_w75_6_c10 & bh1112_w74_10_c10 & bh1112_w73_6_c10 & bh1112_w72_10_c10 & bh1112_w71_6_c10 & bh1112_w70_10_c10 & bh1112_w69_7_c10 & bh1112_w68_11_c10 & bh1112_w67_7_c10 & bh1112_w66_11_c10 & bh1112_w65_7_c10 & bh1112_w64_11_c10 & bh1112_w63_6_c10 & bh1112_w62_10_c10 & bh1112_w61_7_c10 & bh1112_w60_10_c10 & bh1112_w59_9_c10 & bh1112_w58_12_c10 & bh1112_w57_11_c10 & bh1112_w56_12_c10 & bh1112_w55_16_c10 & bh1112_w54_16_c10 & bh1112_w53_19_c10 & bh1112_w52_21_c10 & bh1112_w51_24_c10 & bh1112_w50_26_c10 & bh1112_w49_31_c10 & bh1112_w48_32_c10 & bh1112_w47_34_c10 & bh1112_w46_36_c10 & bh1112_w45_40_c10 & bh1112_w44_41_c10;
   bitheapFinalAdd_bh1112_In1_c10 <= "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & bh1112_w84_1_c10 & "0" & bh1112_w82_3_c10 & "0" & bh1112_w80_5_c10 & "0" & bh1112_w78_7_c10 & "0" & bh1112_w76_9_c10 & "0" & bh1112_w74_11_c10 & "0" & bh1112_w72_11_c10 & "0" & bh1112_w70_11_c10 & "0" & bh1112_w68_12_c10 & "0" & bh1112_w66_12_c10 & "0" & "0" & bh1112_w63_7_c10 & "0" & bh1112_w61_8_c10 & "0" & "0" & "0" & bh1112_w57_12_c10 & "0" & bh1112_w55_17_c10 & "0" & bh1112_w53_20_c10 & "0" & bh1112_w51_25_c10 & "0" & bh1112_w49_32_c10 & "0" & bh1112_w47_35_c10 & "0" & bh1112_w45_41_c10 & bh1112_w44_42_c10;
   bitheapFinalAdd_bh1112_Cin_c0 <= '0';

   bitheapFinalAdd_bh1112: IntAdder_50_Freq300_uid1699
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 Cin => bitheapFinalAdd_bh1112_Cin_c0,
                 X => bitheapFinalAdd_bh1112_In0_c10,
                 Y => bitheapFinalAdd_bh1112_In1_c10,
                 R => bitheapFinalAdd_bh1112_Out_c11);
   bitheapResult_bh1112_c11 <= bitheapFinalAdd_bh1112_Out_c11(48 downto 0) & tmp_bitheapResult_bh1112_43_c11;
   R <= bitheapResult_bh1112_c11(92 downto 45);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_57_Freq300_uid1702
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_57_Freq300_uid1702 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(56 downto 0);
          Y : in  std_logic_vector(56 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of IntAdder_57_Freq300_uid1702 is
signal Rtmp_c11 :  std_logic_vector(56 downto 0);
signal X_c6, X_c7, X_c8, X_c9, X_c10, X_c11 :  std_logic_vector(56 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               X_c6 <= X;
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               X_c7 <= X_c6;
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               X_c8 <= X_c7;
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               X_c9 <= X_c8;
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               X_c10 <= X_c9;
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               X_c11 <= X_c10;
               Cin_c11 <= Cin_c10;
            end if;
         end if;
      end process;
   Rtmp_c11 <= X_c11 + Y + Cin_c11;
   R <= Rtmp_c11;
end architecture;

--------------------------------------------------------------------------------
--                           Exp_11_52_Freq300_uid6
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca (2008-2021)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: ufixX_i XSign
-- Output signals: expY K

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Exp_11_52_Freq300_uid6 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          ufixX_i : in  std_logic_vector(65 downto 0);
          XSign : in  std_logic;
          expY : out  std_logic_vector(56 downto 0);
          K : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of Exp_11_52_Freq300_uid6 is
   component FixRealKCM_Freq300_uid8 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(12 downto 0);
             R : out  std_logic_vector(10 downto 0)   );
   end component;

   component FixRealKCM_Freq300_uid35 is
      port ( clk, ce_3 : in std_logic;
             X : in  std_logic_vector(10 downto 0);
             R : out  std_logic_vector(66 downto 0)   );
   end component;

   component IntAdder_56_Freq300_uid48 is
      port ( clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
             X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(55 downto 0)   );
   end component;

   component FixFunctionByTable_Freq300_uid50 is
      port ( clk, ce_5 : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(56 downto 0)   );
   end component;

   component FixFunctionByPiecewisePoly_Freq300_uid59 is
      port ( clk, ce_5, ce_6, ce_7, ce_8 : in std_logic;
             X : in  std_logic_vector(35 downto 0);
             Y : out  std_logic_vector(35 downto 0)   );
   end component;

   component IntAdder_47_Freq300_uid1108 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(46 downto 0);
             Y : in  std_logic_vector(46 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(46 downto 0)   );
   end component;

   component IntMultiplier_46x47_48_Freq300_uid1110 is
      port ( clk, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(45 downto 0);
             Y : in  std_logic_vector(46 downto 0);
             R : out  std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_57_Freq300_uid1702 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(56 downto 0);
             Y : in  std_logic_vector(56 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(56 downto 0)   );
   end component;

signal ufixX_c2 :  unsigned(9+56 downto 0);
signal xMulIn_c2 :  unsigned(9+3 downto 0);
signal absK_c2, absK_c3 :  std_logic_vector(10 downto 0);
signal minusAbsK_c3 :  std_logic_vector(11 downto 0);
signal absKLog2_c3 :  std_logic_vector(66 downto 0);
signal subOp1_c2 :  std_logic_vector(55 downto 0);
signal subOp2_c3 :  std_logic_vector(55 downto 0);
signal Y_c4 :  std_logic_vector(55 downto 0);
signal A_c4 :  std_logic_vector(9 downto 0);
signal Z_c4 :  std_logic_vector(45 downto 0);
signal expA_c5 :  std_logic_vector(56 downto 0);
signal Ztrunc_c4 :  std_logic_vector(35 downto 0);
signal expZmZm1_c8 :  std_logic_vector(35 downto 0);
signal expZm1adderX_c4 :  std_logic_vector(46 downto 0);
signal expZm1adderY_c8 :  std_logic_vector(46 downto 0);
signal expZm1_c9 :  std_logic_vector(46 downto 0);
signal expArounded_c5 :  std_logic_vector(45 downto 0);
signal lowerProduct_c11 :  std_logic_vector(47 downto 0);
signal extendedLowerProduct_c11 :  std_logic_vector(56 downto 0);
signal XSign_c1, XSign_c2, XSign_c3 :  std_logic;
constant g: positive := 4;
constant wE: positive := 11;
constant wF: positive := 52;
constant wFIn: positive := 52;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               XSign_c1 <= XSign;
            end if;
            if ce_2 = '1' then
               XSign_c2 <= XSign_c1;
            end if;
            if ce_3 = '1' then
               absK_c3 <= absK_c2;
               XSign_c3 <= XSign_c2;
            end if;
            if ce_4 = '1' then
            end if;
            if ce_5 = '1' then
            end if;
            if ce_6 = '1' then
            end if;
            if ce_7 = '1' then
            end if;
            if ce_8 = '1' then
            end if;
            if ce_9 = '1' then
            end if;
            if ce_10 = '1' then
            end if;
            if ce_11 = '1' then
            end if;
         end if;
      end process;
ufixX_c2 <= unsigned(ufixX_i);
   xMulIn_c2 <= ufixX_c2(65 downto 53); -- fix resize from (9, -56) to (9, -3)
   MulInvLog2: FixRealKCM_Freq300_uid8
      port map ( clk  => clk,
                 X => std_logic_vector(xMulIn_c2),
                 R => absK_c2);
   minusAbsK_c3 <= (11 downto 0 => '0') - ('0' & absK_c3);
   K <= minusAbsK_c3 when  XSign_c3='1'   else ('0' & absK_c3);
   MulLog2: FixRealKCM_Freq300_uid35
      port map ( clk  => clk,
                 ce_3 => ce_3,
                 X => absK_c2,
                 R => absKLog2_c3);
   subOp1_c2 <= std_logic_vector(ufixX_c2(55 downto 0)) when XSign_c2='0' else not (std_logic_vector(ufixX_c2(55 downto 0)));
   subOp2_c3 <= absKLog2_c3(55 downto 0) when XSign_c3='1' else not (absKLog2_c3(55 downto 0));
   theYAdder: IntAdder_56_Freq300_uid48
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 Cin => '1',
                 X => subOp1_c2,
                 Y => subOp2_c3,
                 R => Y_c4);
   -- Now compute the exp of this fixed-point value
   A_c4 <= Y_c4(55 downto 46);
   Z_c4 <= Y_c4(45 downto 0);
   ExpATable: FixFunctionByTable_Freq300_uid50
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 X => A_c4,
                 Y => expA_c5);
   Ztrunc_c4 <= Z_c4(45 downto 10);
   poly: FixFunctionByPiecewisePoly_Freq300_uid59
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 X => Ztrunc_c4,
                 Y => expZmZm1_c8);
   -- Computing Z + (exp(Z)-1-Z)
   expZm1adderX_c4 <= '0' & Z_c4;
   expZm1adderY_c8 <= (10 downto 0 => '0') & expZmZm1_c8 ;
   Adder_expZm1: IntAdder_47_Freq300_uid1108
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 Cin => '0',
                 X => expZm1adderX_c4,
                 Y => expZm1adderY_c8,
                 R => expZm1_c9);
   -- Truncating expA to the same accuracy as expZm1
   expArounded_c5 <= expA_c5(56 downto 11);
   TheLowerProduct: IntMultiplier_46x47_48_Freq300_uid1110
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 X => expArounded_c5,
                 Y => expZm1_c9,
                 R => lowerProduct_c11);
   extendedLowerProduct_c11 <= ((56 downto 48 => '0') & lowerProduct_c11(47 downto 0));
   -- Final addition -- the product MSB bit weight is -k+2 = -8
   TheFinalAdder: IntAdder_57_Freq300_uid1702
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 Cin => '0',
                 X => expA_c5,
                 Y => extendedLowerProduct_c11,
                 R => expY);
end architecture;

--------------------------------------------------------------------------------
--                        IntAdder_65_Freq300_uid1705
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_65_Freq300_uid1705 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
          X : in  std_logic_vector(64 downto 0);
          Y : in  std_logic_vector(64 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(64 downto 0)   );
end entity;

architecture arch of IntAdder_65_Freq300_uid1705 is
signal Rtmp_c12 :  std_logic_vector(64 downto 0);
signal Y_c12 :  std_logic_vector(64 downto 0);
signal Cin_c1, Cin_c2, Cin_c3, Cin_c4, Cin_c5, Cin_c6, Cin_c7, Cin_c8, Cin_c9, Cin_c10, Cin_c11, Cin_c12 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               Cin_c2 <= Cin_c1;
            end if;
            if ce_3 = '1' then
               Cin_c3 <= Cin_c2;
            end if;
            if ce_4 = '1' then
               Cin_c4 <= Cin_c3;
            end if;
            if ce_5 = '1' then
               Cin_c5 <= Cin_c4;
            end if;
            if ce_6 = '1' then
               Cin_c6 <= Cin_c5;
            end if;
            if ce_7 = '1' then
               Cin_c7 <= Cin_c6;
            end if;
            if ce_8 = '1' then
               Cin_c8 <= Cin_c7;
            end if;
            if ce_9 = '1' then
               Cin_c9 <= Cin_c8;
            end if;
            if ce_10 = '1' then
               Cin_c10 <= Cin_c9;
            end if;
            if ce_11 = '1' then
               Cin_c11 <= Cin_c10;
            end if;
            if ce_12 = '1' then
               Y_c12 <= Y;
               Cin_c12 <= Cin_c11;
            end if;
         end if;
      end process;
   Rtmp_c12 <= X + Y_c12 + Cin_c12;
   R <= Rtmp_c12;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointExponential
--                         (FPExp_11_52_Freq300_uid2)
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca (2008-2021)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointExponential is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointExponential is
   component LeftShifter53_by_max_65_Freq300_uid4 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             S : in  std_logic_vector(6 downto 0);
             R : out  std_logic_vector(117 downto 0)   );
   end component;

   component Exp_11_52_Freq300_uid6 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             ufixX_i : in  std_logic_vector(65 downto 0);
             XSign : in  std_logic;
             expY : out  std_logic_vector(56 downto 0);
             K : out  std_logic_vector(11 downto 0)   );
   end component;

   component IntAdder_65_Freq300_uid1705 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
             X : in  std_logic_vector(64 downto 0);
             Y : in  std_logic_vector(64 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(64 downto 0)   );
   end component;

signal Xexn_c0, Xexn_c1, Xexn_c2, Xexn_c3, Xexn_c4, Xexn_c5, Xexn_c6, Xexn_c7, Xexn_c8, Xexn_c9, Xexn_c10, Xexn_c11, Xexn_c12 :  std_logic_vector(1 downto 0);
signal XSign_c0, XSign_c1, XSign_c2, XSign_c3, XSign_c4, XSign_c5, XSign_c6, XSign_c7, XSign_c8, XSign_c9, XSign_c10, XSign_c11, XSign_c12 :  std_logic;
signal XexpField_c0 :  std_logic_vector(10 downto 0);
signal Xfrac_c0 :  unsigned(-1+52 downto 0);
signal e0_c0 :  std_logic_vector(12 downto 0);
signal shiftVal_c0 :  std_logic_vector(12 downto 0);
signal resultWillBeOne_c0, resultWillBeOne_c1, resultWillBeOne_c2 :  std_logic;
signal mXu_c0 :  unsigned(0+52 downto 0);
signal maxShift_c0 :  std_logic_vector(11 downto 0);
signal overflow0_c0 :  std_logic;
signal shiftValIn_c0 :  std_logic_vector(6 downto 0);
signal fixX0_c2 :  std_logic_vector(117 downto 0);
signal ufixX_c2 :  unsigned(9+56 downto 0);
signal expY_c11, expY_c12 :  std_logic_vector(56 downto 0);
signal K_c3, K_c4, K_c5, K_c6, K_c7, K_c8, K_c9, K_c10, K_c11 :  std_logic_vector(11 downto 0);
signal needNoNorm_c11, needNoNorm_c12 :  std_logic;
signal preRoundBiasSig_c12 :  std_logic_vector(64 downto 0);
signal roundBit_c11 :  std_logic;
signal roundNormAddend_c11 :  std_logic_vector(64 downto 0);
signal roundedExpSigRes_c12 :  std_logic_vector(64 downto 0);
signal roundedExpSig_c12 :  std_logic_vector(64 downto 0);
signal ofl1_c0, ofl1_c1, ofl1_c2, ofl1_c3, ofl1_c4, ofl1_c5, ofl1_c6, ofl1_c7, ofl1_c8, ofl1_c9, ofl1_c10, ofl1_c11, ofl1_c12 :  std_logic;
signal ofl2_c12 :  std_logic;
signal ofl3_c0, ofl3_c1, ofl3_c2, ofl3_c3, ofl3_c4, ofl3_c5, ofl3_c6, ofl3_c7, ofl3_c8, ofl3_c9, ofl3_c10, ofl3_c11, ofl3_c12 :  std_logic;
signal ofl_c12 :  std_logic;
signal ufl1_c12 :  std_logic;
signal ufl2_c0, ufl2_c1, ufl2_c2, ufl2_c3, ufl2_c4, ufl2_c5, ufl2_c6, ufl2_c7, ufl2_c8, ufl2_c9, ufl2_c10, ufl2_c11, ufl2_c12 :  std_logic;
signal ufl3_c0, ufl3_c1, ufl3_c2, ufl3_c3, ufl3_c4, ufl3_c5, ufl3_c6, ufl3_c7, ufl3_c8, ufl3_c9, ufl3_c10, ufl3_c11, ufl3_c12 :  std_logic;
signal ufl_c12 :  std_logic;
signal Rexn_c12 :  std_logic_vector(1 downto 0);
constant g: positive := 4;
constant wE: positive := 11;
constant wF: positive := 52;
constant wFIn: positive := 52;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Xexn_c1 <= Xexn_c0;
               XSign_c1 <= XSign_c0;
               resultWillBeOne_c1 <= resultWillBeOne_c0;
               ofl1_c1 <= ofl1_c0;
               ofl3_c1 <= ofl3_c0;
               ufl2_c1 <= ufl2_c0;
               ufl3_c1 <= ufl3_c0;
            end if;
            if ce_2 = '1' then
               Xexn_c2 <= Xexn_c1;
               XSign_c2 <= XSign_c1;
               resultWillBeOne_c2 <= resultWillBeOne_c1;
               ofl1_c2 <= ofl1_c1;
               ofl3_c2 <= ofl3_c1;
               ufl2_c2 <= ufl2_c1;
               ufl3_c2 <= ufl3_c1;
            end if;
            if ce_3 = '1' then
               Xexn_c3 <= Xexn_c2;
               XSign_c3 <= XSign_c2;
               ofl1_c3 <= ofl1_c2;
               ofl3_c3 <= ofl3_c2;
               ufl2_c3 <= ufl2_c2;
               ufl3_c3 <= ufl3_c2;
            end if;
            if ce_4 = '1' then
               Xexn_c4 <= Xexn_c3;
               XSign_c4 <= XSign_c3;
               K_c4 <= K_c3;
               ofl1_c4 <= ofl1_c3;
               ofl3_c4 <= ofl3_c3;
               ufl2_c4 <= ufl2_c3;
               ufl3_c4 <= ufl3_c3;
            end if;
            if ce_5 = '1' then
               Xexn_c5 <= Xexn_c4;
               XSign_c5 <= XSign_c4;
               K_c5 <= K_c4;
               ofl1_c5 <= ofl1_c4;
               ofl3_c5 <= ofl3_c4;
               ufl2_c5 <= ufl2_c4;
               ufl3_c5 <= ufl3_c4;
            end if;
            if ce_6 = '1' then
               Xexn_c6 <= Xexn_c5;
               XSign_c6 <= XSign_c5;
               K_c6 <= K_c5;
               ofl1_c6 <= ofl1_c5;
               ofl3_c6 <= ofl3_c5;
               ufl2_c6 <= ufl2_c5;
               ufl3_c6 <= ufl3_c5;
            end if;
            if ce_7 = '1' then
               Xexn_c7 <= Xexn_c6;
               XSign_c7 <= XSign_c6;
               K_c7 <= K_c6;
               ofl1_c7 <= ofl1_c6;
               ofl3_c7 <= ofl3_c6;
               ufl2_c7 <= ufl2_c6;
               ufl3_c7 <= ufl3_c6;
            end if;
            if ce_8 = '1' then
               Xexn_c8 <= Xexn_c7;
               XSign_c8 <= XSign_c7;
               K_c8 <= K_c7;
               ofl1_c8 <= ofl1_c7;
               ofl3_c8 <= ofl3_c7;
               ufl2_c8 <= ufl2_c7;
               ufl3_c8 <= ufl3_c7;
            end if;
            if ce_9 = '1' then
               Xexn_c9 <= Xexn_c8;
               XSign_c9 <= XSign_c8;
               K_c9 <= K_c8;
               ofl1_c9 <= ofl1_c8;
               ofl3_c9 <= ofl3_c8;
               ufl2_c9 <= ufl2_c8;
               ufl3_c9 <= ufl3_c8;
            end if;
            if ce_10 = '1' then
               Xexn_c10 <= Xexn_c9;
               XSign_c10 <= XSign_c9;
               K_c10 <= K_c9;
               ofl1_c10 <= ofl1_c9;
               ofl3_c10 <= ofl3_c9;
               ufl2_c10 <= ufl2_c9;
               ufl3_c10 <= ufl3_c9;
            end if;
            if ce_11 = '1' then
               Xexn_c11 <= Xexn_c10;
               XSign_c11 <= XSign_c10;
               K_c11 <= K_c10;
               ofl1_c11 <= ofl1_c10;
               ofl3_c11 <= ofl3_c10;
               ufl2_c11 <= ufl2_c10;
               ufl3_c11 <= ufl3_c10;
            end if;
            if ce_12 = '1' then
               Xexn_c12 <= Xexn_c11;
               XSign_c12 <= XSign_c11;
               expY_c12 <= expY_c11;
               needNoNorm_c12 <= needNoNorm_c11;
               ofl1_c12 <= ofl1_c11;
               ofl3_c12 <= ofl3_c11;
               ufl2_c12 <= ufl2_c11;
               ufl3_c12 <= ufl3_c11;
            end if;
         end if;
      end process;
   Xexn_c0 <= X(wE+wFIn+2 downto wE+wFIn+1);
   XSign_c0 <= X(wE+wFIn);
   XexpField_c0 <= X(wE+wFIn-1 downto wFIn);
   Xfrac_c0 <= unsigned(X(wFIn-1 downto 0));
   e0_c0 <= conv_std_logic_vector(967, wE+2);  -- bias - (wF+g)
   shiftVal_c0 <= ("00" & XexpField_c0) - e0_c0; -- for a left shift
   -- underflow when input is shifted to zero (shiftval<0), in which case exp = 1
   resultWillBeOne_c0 <= shiftVal_c0(wE+1);
   --  mantissa with implicit bit
   mXu_c0 <= "1" & Xfrac_c0;
   -- Partial overflow detection
   maxShift_c0 <= conv_std_logic_vector(65, wE+1);  -- wE-2 + wF+g
   overflow0_c0 <= not shiftVal_c0(wE+1) when shiftVal_c0(wE downto 0) > maxShift_c0 else '0';
   shiftValIn_c0 <= shiftVal_c0(6 downto 0);
   mantissa_shift: LeftShifter53_by_max_65_Freq300_uid4
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 S => shiftValIn_c0,
                 X => std_logic_vector(mXu_c0),
                 R => fixX0_c2);
   ufixX_c2 <=  unsigned(fixX0_c2(117 downto 52)) when resultWillBeOne_c2='0' else "000000000000000000000000000000000000000000000000000000000000000000";
   exp_helper: Exp_11_52_Freq300_uid6
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 XSign => XSign_c0,
                 ufixX_i => std_logic_vector(ufixX_c2),
                 K => K_c3,
                 expY => expY_c11);
   needNoNorm_c11 <= expY_c11(56);
   -- Rounding: all this should consume one row of LUTs
   preRoundBiasSig_c12 <= conv_std_logic_vector(1023, wE+2)  & expY_c12(55 downto 4) when needNoNorm_c12 = '1'
      else conv_std_logic_vector(1022, wE+2)  & expY_c12(54 downto 3) ;
   roundBit_c11 <= expY_c11(3)  when needNoNorm_c11 = '1'    else expY_c11(2) ;
   roundNormAddend_c11 <= K_c11(11) & K_c11 & (51 downto 1 => '0') & roundBit_c11;
   roundedExpSigOperandAdder: IntAdder_65_Freq300_uid1705
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 Cin => '0',
                 X => preRoundBiasSig_c12,
                 Y => roundNormAddend_c11,
                 R => roundedExpSigRes_c12);
   roundedExpSig_c12 <= roundedExpSigRes_c12 when Xexn_c12="01" else  "000" & (wE-2 downto 0 => '1') & (wF-1 downto 0 => '0');
   ofl1_c0 <= not XSign_c0 and overflow0_c0 and (not Xexn_c0(1) and Xexn_c0(0)); -- input positive, normal,  very large
   ofl2_c12 <= not XSign_c12 and (roundedExpSig_c12(wE+wF) and not roundedExpSig_c12(wE+wF+1)) and (not Xexn_c12(1) and Xexn_c12(0)); -- input positive, normal, overflowed
   ofl3_c0 <= not XSign_c0 and Xexn_c0(1) and not Xexn_c0(0);  -- input was -infty
   ofl_c12 <= ofl1_c12 or ofl2_c12 or ofl3_c12;
   ufl1_c12 <= (roundedExpSig_c12(wE+wF) and roundedExpSig_c12(wE+wF+1))  and (not Xexn_c12(1) and Xexn_c12(0)); -- input normal
   ufl2_c0 <= XSign_c0 and Xexn_c0(1) and not Xexn_c0(0);  -- input was -infty
   ufl3_c0 <= XSign_c0 and overflow0_c0  and (not Xexn_c0(1) and Xexn_c0(0)); -- input negative, normal,  very large
   ufl_c12 <= ufl1_c12 or ufl2_c12 or ufl3_c12;
   Rexn_c12 <= "11" when Xexn_c12 = "11"
      else "10" when ofl_c12='1'
      else "00" when ufl_c12='1'
      else "01";
   R <= Rexn_c12 & '0' & roundedExpSig_c12(62 downto 0);
end architecture;



