--------------------------------------------------------------------------------
--                  FixRealKCM_Freq800_uid8_T0_Freq800_uid11
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq800_uid8_T0_Freq800_uid11 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq800_uid8_T0_Freq800_uid11 is
signal Y0 :  std_logic_vector(11 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(11 downto 0);
begin
   with X  select  Y0 <= 
      "000000001000" when "00000",
      "000001100100" when "00001",
      "000011000001" when "00010",
      "000100011101" when "00011",
      "000101111001" when "00100",
      "000111010110" when "00101",
      "001000110010" when "00110",
      "001010001110" when "00111",
      "001011101011" when "01000",
      "001101000111" when "01001",
      "001110100011" when "01010",
      "010000000000" when "01011",
      "010001011100" when "01100",
      "010010111000" when "01101",
      "010100010101" when "01110",
      "010101110001" when "01111",
      "010111001101" when "10000",
      "011000101010" when "10001",
      "011010000110" when "10010",
      "011011100010" when "10011",
      "011100111111" when "10100",
      "011110011011" when "10101",
      "011111110111" when "10110",
      "100001010100" when "10111",
      "100010110000" when "11000",
      "100100001100" when "11001",
      "100101101001" when "11010",
      "100111000101" when "11011",
      "101000100001" when "11100",
      "101001111110" when "11101",
      "101011011010" when "11110",
      "101100110110" when "11111",
      "------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                  FixRealKCM_Freq800_uid8_T1_Freq800_uid14
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq800_uid8_T1_Freq800_uid14 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq800_uid8_T1_Freq800_uid14 is
signal Y0 :  std_logic_vector(6 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(6 downto 0);
begin
   with X  select  Y0 <= 
      "0000000" when "00000",
      "0000011" when "00001",
      "0000110" when "00010",
      "0001001" when "00011",
      "0001100" when "00100",
      "0001110" when "00101",
      "0010001" when "00110",
      "0010100" when "00111",
      "0010111" when "01000",
      "0011010" when "01001",
      "0011101" when "01010",
      "0100000" when "01011",
      "0100011" when "01100",
      "0100110" when "01101",
      "0101000" when "01110",
      "0101011" when "01111",
      "0101110" when "10000",
      "0110001" when "10001",
      "0110100" when "10010",
      "0110111" when "10011",
      "0111010" when "10100",
      "0111101" when "10101",
      "0111111" when "10110",
      "1000010" when "10111",
      "1000101" when "11000",
      "1001000" when "11001",
      "1001011" when "11010",
      "1001110" when "11011",
      "1010001" when "11100",
      "1010100" when "11101",
      "1010111" when "11110",
      "1011001" when "11111",
      "-------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq800_uid20_T0_Freq800_uid23
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq800_uid20_T0_Freq800_uid23 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq800_uid20_T0_Freq800_uid23 is
signal Y0 :  std_logic_vector(34 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(34 downto 0);
begin
   with X  select  Y0 <= 
      "00000000000000000000000000000000000" when "00000",
      "00000101100010111001000010111111110" when "00001",
      "00001011000101110010000101111111100" when "00010",
      "00010000101000101011001000111111010" when "00011",
      "00010110001011100100001011111111000" when "00100",
      "00011011101110011101001110111110110" when "00101",
      "00100001010001010110010001111110100" when "00110",
      "00100110110100001111010100111110010" when "00111",
      "00101100010111001000010111111110000" when "01000",
      "00110001111010000001011010111101110" when "01001",
      "00110111011100111010011101111101100" when "01010",
      "00111100111111110011100000111101010" when "01011",
      "01000010100010101100100011111100111" when "01100",
      "01001000000101100101100110111100101" when "01101",
      "01001101101000011110101001111100011" when "01110",
      "01010011001011010111101100111100001" when "01111",
      "01011000101110010000101111111011111" when "10000",
      "01011110010001001001110010111011101" when "10001",
      "01100011110100000010110101111011011" when "10010",
      "01101001010110111011111000111011001" when "10011",
      "01101110111001110100111011111010111" when "10100",
      "01110100011100101101111110111010101" when "10101",
      "01111001111111100111000001111010011" when "10110",
      "01111111100010100000000100111010001" when "10111",
      "10000101000101011001000111111001111" when "11000",
      "10001010101000010010001010111001101" when "11001",
      "10010000001011001011001101111001011" when "11010",
      "10010101101110000100010000111001001" when "11011",
      "10011011010000111101010011111000111" when "11100",
      "10100000110011110110010110111000101" when "11101",
      "10100110010110101111011001111000011" when "11110",
      "10101011111001101000011100111000001" when "11111",
      "-----------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                 FixRealKCM_Freq800_uid20_T1_Freq800_uid26
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq800_uid20_T1_Freq800_uid26 is
    port (X : in  std_logic_vector(2 downto 0);
          Y : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq800_uid20_T1_Freq800_uid26 is
signal Y0 :  std_logic_vector(29 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(29 downto 0);
begin
   with X  select  Y0 <= 
      "000000000000000000000000000000" when "000",
      "000101100010111001000011000000" when "001",
      "001011000101110010000101111111" when "010",
      "010000101000101011001000111111" when "011",
      "010110001011100100001011111111" when "100",
      "011011101110011101001110111111" when "101",
      "100001010001010110010001111110" when "110",
      "100110110100001111010100111110" when "111",
      "------------------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--          compressedTable_Freq800_uid37_subsampling_Freq800_uid39
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity compressedTable_Freq800_uid37_subsampling_Freq800_uid39 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of compressedTable_Freq800_uid37_subsampling_Freq800_uid39 is
signal Y0 :  std_logic_vector(8 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(8 downto 0);
begin
   with X  select  Y0 <= 
      "100000000" when "0000000",
      "100000010" when "0000001",
      "100000100" when "0000010",
      "100000110" when "0000011",
      "100001000" when "0000100",
      "100001010" when "0000101",
      "100001100" when "0000110",
      "100001110" when "0000111",
      "100010000" when "0001000",
      "100010010" when "0001001",
      "100010100" when "0001010",
      "100010110" when "0001011",
      "100011001" when "0001100",
      "100011011" when "0001101",
      "100011101" when "0001110",
      "100011111" when "0001111",
      "100100010" when "0010000",
      "100100100" when "0010001",
      "100100110" when "0010010",
      "100101000" when "0010011",
      "100101011" when "0010100",
      "100101101" when "0010101",
      "100110000" when "0010110",
      "100110010" when "0010111",
      "100110100" when "0011000",
      "100110111" when "0011001",
      "100111001" when "0011010",
      "100111100" when "0011011",
      "100111110" when "0011100",
      "101000001" when "0011101",
      "101000011" when "0011110",
      "101000110" when "0011111",
      "101001000" when "0100000",
      "101001011" when "0100001",
      "101001101" when "0100010",
      "101010000" when "0100011",
      "101010011" when "0100100",
      "101010101" when "0100101",
      "101011000" when "0100110",
      "101011011" when "0100111",
      "101011101" when "0101000",
      "101100000" when "0101001",
      "101100011" when "0101010",
      "101100110" when "0101011",
      "101101001" when "0101100",
      "101101011" when "0101101",
      "101101110" when "0101110",
      "101110001" when "0101111",
      "101110100" when "0110000",
      "101110111" when "0110001",
      "101111010" when "0110010",
      "101111101" when "0110011",
      "110000000" when "0110100",
      "110000011" when "0110101",
      "110000110" when "0110110",
      "110001001" when "0110111",
      "110001100" when "0111000",
      "110001111" when "0111001",
      "110010010" when "0111010",
      "110010101" when "0111011",
      "110011001" when "0111100",
      "110011100" when "0111101",
      "110011111" when "0111110",
      "110100010" when "0111111",
      "010011011" when "1000000",
      "010011100" when "1000001",
      "010011101" when "1000010",
      "010011110" when "1000011",
      "010100000" when "1000100",
      "010100001" when "1000101",
      "010100010" when "1000110",
      "010100011" when "1000111",
      "010100101" when "1001000",
      "010100110" when "1001001",
      "010100111" when "1001010",
      "010101001" when "1001011",
      "010101010" when "1001100",
      "010101011" when "1001101",
      "010101101" when "1001110",
      "010101110" when "1001111",
      "010101111" when "1010000",
      "010110001" when "1010001",
      "010110010" when "1010010",
      "010110100" when "1010011",
      "010110101" when "1010100",
      "010110110" when "1010101",
      "010111000" when "1010110",
      "010111001" when "1010111",
      "010111011" when "1011000",
      "010111100" when "1011001",
      "010111110" when "1011010",
      "010111111" when "1011011",
      "011000001" when "1011100",
      "011000010" when "1011101",
      "011000100" when "1011110",
      "011000101" when "1011111",
      "011000111" when "1100000",
      "011001000" when "1100001",
      "011001010" when "1100010",
      "011001100" when "1100011",
      "011001101" when "1100100",
      "011001111" when "1100101",
      "011010000" when "1100110",
      "011010010" when "1100111",
      "011010100" when "1101000",
      "011010101" when "1101001",
      "011010111" when "1101010",
      "011011001" when "1101011",
      "011011010" when "1101100",
      "011011100" when "1101101",
      "011011110" when "1101110",
      "011100000" when "1101111",
      "011100001" when "1110000",
      "011100011" when "1110001",
      "011100101" when "1110010",
      "011100111" when "1110011",
      "011101001" when "1110100",
      "011101010" when "1110101",
      "011101100" when "1110110",
      "011101110" when "1110111",
      "011110000" when "1111000",
      "011110010" when "1111001",
      "011110100" when "1111010",
      "011110110" when "1111011",
      "011111000" when "1111100",
      "011111010" when "1111101",
      "011111100" when "1111110",
      "011111110" when "1111111",
      "---------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                      FixFunctionByTable_Freq800_uid44
-- Evaluator for exp(x*1b-10)-1-x*1b-10 on [0,1) for lsbIn=-7 (wIn=7), msbout=-22, lsbOut=-27 (wOut=6). Out interval: [0; 4.69567e-07]. Output is unsigned

-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq800_uid44 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq800_uid44 is
signal Y0 :  std_logic_vector(5 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(5 downto 0);
begin
   with X  select  Y0 <= 
      "000000" when "0000000",
      "000000" when "0000001",
      "000000" when "0000010",
      "000000" when "0000011",
      "000000" when "0000100",
      "000000" when "0000101",
      "000000" when "0000110",
      "000000" when "0000111",
      "000000" when "0001000",
      "000000" when "0001001",
      "000000" when "0001010",
      "000000" when "0001011",
      "000001" when "0001100",
      "000001" when "0001101",
      "000001" when "0001110",
      "000001" when "0001111",
      "000001" when "0010000",
      "000001" when "0010001",
      "000001" when "0010010",
      "000001" when "0010011",
      "000010" when "0010100",
      "000010" when "0010101",
      "000010" when "0010110",
      "000010" when "0010111",
      "000010" when "0011000",
      "000010" when "0011001",
      "000011" when "0011010",
      "000011" when "0011011",
      "000011" when "0011100",
      "000011" when "0011101",
      "000100" when "0011110",
      "000100" when "0011111",
      "000100" when "0100000",
      "000100" when "0100001",
      "000101" when "0100010",
      "000101" when "0100011",
      "000101" when "0100100",
      "000101" when "0100101",
      "000110" when "0100110",
      "000110" when "0100111",
      "000110" when "0101000",
      "000111" when "0101001",
      "000111" when "0101010",
      "000111" when "0101011",
      "001000" when "0101100",
      "001000" when "0101101",
      "001000" when "0101110",
      "001001" when "0101111",
      "001001" when "0110000",
      "001001" when "0110001",
      "001010" when "0110010",
      "001010" when "0110011",
      "001011" when "0110100",
      "001011" when "0110101",
      "001011" when "0110110",
      "001100" when "0110111",
      "001100" when "0111000",
      "001101" when "0111001",
      "001101" when "0111010",
      "001110" when "0111011",
      "001110" when "0111100",
      "001111" when "0111101",
      "001111" when "0111110",
      "010000" when "0111111",
      "010000" when "1000000",
      "010001" when "1000001",
      "010001" when "1000010",
      "010010" when "1000011",
      "010010" when "1000100",
      "010011" when "1000101",
      "010011" when "1000110",
      "010100" when "1000111",
      "010100" when "1001000",
      "010101" when "1001001",
      "010101" when "1001010",
      "010110" when "1001011",
      "010111" when "1001100",
      "010111" when "1001101",
      "011000" when "1001110",
      "011000" when "1001111",
      "011001" when "1010000",
      "011010" when "1010001",
      "011010" when "1010010",
      "011011" when "1010011",
      "011100" when "1010100",
      "011100" when "1010101",
      "011101" when "1010110",
      "011110" when "1010111",
      "011110" when "1011000",
      "011111" when "1011001",
      "100000" when "1011010",
      "100000" when "1011011",
      "100001" when "1011100",
      "100010" when "1011101",
      "100011" when "1011110",
      "100011" when "1011111",
      "100100" when "1100000",
      "100101" when "1100001",
      "100110" when "1100010",
      "100110" when "1100011",
      "100111" when "1100100",
      "101000" when "1100101",
      "101001" when "1100110",
      "101001" when "1100111",
      "101010" when "1101000",
      "101011" when "1101001",
      "101100" when "1101010",
      "101101" when "1101011",
      "101110" when "1101100",
      "101110" when "1101101",
      "101111" when "1101110",
      "110000" when "1101111",
      "110001" when "1110000",
      "110010" when "1110001",
      "110011" when "1110010",
      "110100" when "1110011",
      "110101" when "1110100",
      "110101" when "1110101",
      "110110" when "1110110",
      "110111" when "1110111",
      "111000" when "1111000",
      "111001" when "1111001",
      "111010" when "1111010",
      "111011" when "1111011",
      "111100" when "1111100",
      "111101" when "1111101",
      "111110" when "1111110",
      "111111" when "1111111",
      "------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid62
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid62 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid62 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid67
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid67 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid67 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid76
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid76 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid76 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid81
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid81 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid81 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid88
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid88 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid88 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid93
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid93 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid93 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid98
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid98 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid98 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid105
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid105 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid105 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid110
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid110 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid110 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid115
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid115 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid115 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid120
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid120 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid120 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid129
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid129 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid129 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid134
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid134 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid134 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid139
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid139 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid139 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid144
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid144 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid144 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid151
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid151 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid151 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid156
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid156 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid156 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid161
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid161 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid161 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid166
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid166 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid166 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid171
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid171 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid171 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid176
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid176 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid176 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid181
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid181 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid181 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid186
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid186 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid186 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid191
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid191 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid191 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid196
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid196 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid196 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid201
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid201 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid201 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid206
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid206 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid206 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid211
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid211 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid211 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid216
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid216 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid216 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid221
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid221 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid221 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid226
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid226 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid226 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid231
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid231 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid231 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid236
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid236 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid236 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid241
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid241 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid241 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid246
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid246 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid246 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid251
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid251 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid251 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid256
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid256 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid256 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid261
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid261 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid261 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq800_uid265
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq800_uid265 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq800_uid265 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq800_uid271
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq800_uid271 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq800_uid271 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq800_uid277
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq800_uid277 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq800_uid277 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq800_uid289
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq800_uid289 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq800_uid289 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                    LeftShifter24_by_max_33_Freq800_uid4
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X S
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter24_by_max_33_Freq800_uid4 is
    port (clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          S : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of LeftShifter24_by_max_33_Freq800_uid4 is
signal ps_c1, ps_c2, ps_c3, ps_c4 :  std_logic_vector(5 downto 0);
signal level0_c0, level0_c1 :  std_logic_vector(23 downto 0);
signal level1_c1 :  std_logic_vector(24 downto 0);
signal level2_c1 :  std_logic_vector(26 downto 0);
signal level3_c1, level3_c2, level3_c3 :  std_logic_vector(30 downto 0);
signal level4_c3 :  std_logic_vector(38 downto 0);
signal level5_c3, level5_c4 :  std_logic_vector(54 downto 0);
signal level6_c4 :  std_logic_vector(86 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               level0_c1 <= level0_c0;
            end if;
            if ce_2 = '1' then
               ps_c2 <= ps_c1;
               level3_c2 <= level3_c1;
            end if;
            if ce_3 = '1' then
               ps_c3 <= ps_c2;
               level3_c3 <= level3_c2;
            end if;
            if ce_4 = '1' then
               ps_c4 <= ps_c3;
               level5_c4 <= level5_c3;
            end if;
         end if;
      end process;
   ps_c1<= S;
   level0_c0<= X;
   level1_c1<= level0_c1 & (0 downto 0 => '0') when ps_c1(0)= '1' else     (0 downto 0 => '0') & level0_c1;
   level2_c1<= level1_c1 & (1 downto 0 => '0') when ps_c1(1)= '1' else     (1 downto 0 => '0') & level1_c1;
   level3_c1<= level2_c1 & (3 downto 0 => '0') when ps_c1(2)= '1' else     (3 downto 0 => '0') & level2_c1;
   level4_c3<= level3_c3 & (7 downto 0 => '0') when ps_c3(3)= '1' else     (7 downto 0 => '0') & level3_c3;
   level5_c3<= level4_c3 & (15 downto 0 => '0') when ps_c3(4)= '1' else     (15 downto 0 => '0') & level4_c3;
   level6_c4<= level5_c4 & (31 downto 0 => '0') when ps_c4(5)= '1' else     (31 downto 0 => '0') & level5_c4;
   R <= level6_c4(56 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_13_Freq800_uid18
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_13_Freq800_uid18 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10 : in std_logic;
          X : in  std_logic_vector(12 downto 0);
          Y : in  std_logic_vector(12 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(12 downto 0)   );
end entity;

architecture arch of IntAdder_13_Freq800_uid18 is
signal Cin_1_c0, Cin_1_c1, Cin_1_c2, Cin_1_c3, Cin_1_c4, Cin_1_c5, Cin_1_c6 :  std_logic;
signal X_1_c5, X_1_c6 :  std_logic_vector(3 downto 0);
signal Y_1_c5, Y_1_c6 :  std_logic_vector(3 downto 0);
signal S_1_c6 :  std_logic_vector(3 downto 0);
signal R_1_c6, R_1_c7, R_1_c8, R_1_c9, R_1_c10 :  std_logic_vector(2 downto 0);
signal Cin_2_c6, Cin_2_c7 :  std_logic;
signal X_2_c5, X_2_c6, X_2_c7 :  std_logic_vector(3 downto 0);
signal Y_2_c5, Y_2_c6, Y_2_c7 :  std_logic_vector(3 downto 0);
signal S_2_c7 :  std_logic_vector(3 downto 0);
signal R_2_c7, R_2_c8, R_2_c9, R_2_c10 :  std_logic_vector(2 downto 0);
signal Cin_3_c7, Cin_3_c8 :  std_logic;
signal X_3_c5, X_3_c6, X_3_c7, X_3_c8 :  std_logic_vector(3 downto 0);
signal Y_3_c5, Y_3_c6, Y_3_c7, Y_3_c8 :  std_logic_vector(3 downto 0);
signal S_3_c8 :  std_logic_vector(3 downto 0);
signal R_3_c8, R_3_c9, R_3_c10 :  std_logic_vector(2 downto 0);
signal Cin_4_c8, Cin_4_c9 :  std_logic;
signal X_4_c5, X_4_c6, X_4_c7, X_4_c8, X_4_c9 :  std_logic_vector(3 downto 0);
signal Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8, Y_4_c9 :  std_logic_vector(3 downto 0);
signal S_4_c9 :  std_logic_vector(3 downto 0);
signal R_4_c9, R_4_c10 :  std_logic_vector(2 downto 0);
signal Cin_5_c9, Cin_5_c10 :  std_logic;
signal X_5_c5, X_5_c6, X_5_c7, X_5_c8, X_5_c9, X_5_c10 :  std_logic_vector(1 downto 0);
signal Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9, Y_5_c10 :  std_logic_vector(1 downto 0);
signal S_5_c10 :  std_logic_vector(1 downto 0);
signal R_5_c10 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_1_c1 <= Cin_1_c0;
            end if;
            if ce_2 = '1' then
               Cin_1_c2 <= Cin_1_c1;
            end if;
            if ce_3 = '1' then
               Cin_1_c3 <= Cin_1_c2;
            end if;
            if ce_4 = '1' then
               Cin_1_c4 <= Cin_1_c3;
            end if;
            if ce_5 = '1' then
               Cin_1_c5 <= Cin_1_c4;
            end if;
            if ce_6 = '1' then
               Cin_1_c6 <= Cin_1_c5;
               X_1_c6 <= X_1_c5;
               Y_1_c6 <= Y_1_c5;
               X_2_c6 <= X_2_c5;
               Y_2_c6 <= Y_2_c5;
               X_3_c6 <= X_3_c5;
               Y_3_c6 <= Y_3_c5;
               X_4_c6 <= X_4_c5;
               Y_4_c6 <= Y_4_c5;
               X_5_c6 <= X_5_c5;
               Y_5_c6 <= Y_5_c5;
            end if;
            if ce_7 = '1' then
               R_1_c7 <= R_1_c6;
               Cin_2_c7 <= Cin_2_c6;
               X_2_c7 <= X_2_c6;
               Y_2_c7 <= Y_2_c6;
               X_3_c7 <= X_3_c6;
               Y_3_c7 <= Y_3_c6;
               X_4_c7 <= X_4_c6;
               Y_4_c7 <= Y_4_c6;
               X_5_c7 <= X_5_c6;
               Y_5_c7 <= Y_5_c6;
            end if;
            if ce_8 = '1' then
               R_1_c8 <= R_1_c7;
               R_2_c8 <= R_2_c7;
               Cin_3_c8 <= Cin_3_c7;
               X_3_c8 <= X_3_c7;
               Y_3_c8 <= Y_3_c7;
               X_4_c8 <= X_4_c7;
               Y_4_c8 <= Y_4_c7;
               X_5_c8 <= X_5_c7;
               Y_5_c8 <= Y_5_c7;
            end if;
            if ce_9 = '1' then
               R_1_c9 <= R_1_c8;
               R_2_c9 <= R_2_c8;
               R_3_c9 <= R_3_c8;
               Cin_4_c9 <= Cin_4_c8;
               X_4_c9 <= X_4_c8;
               Y_4_c9 <= Y_4_c8;
               X_5_c9 <= X_5_c8;
               Y_5_c9 <= Y_5_c8;
            end if;
            if ce_10 = '1' then
               R_1_c10 <= R_1_c9;
               R_2_c10 <= R_2_c9;
               R_3_c10 <= R_3_c9;
               R_4_c10 <= R_4_c9;
               Cin_5_c10 <= Cin_5_c9;
               X_5_c10 <= X_5_c9;
               Y_5_c10 <= Y_5_c9;
            end if;
         end if;
      end process;
   Cin_1_c0 <= Cin;
   X_1_c5 <= '0' & X(2 downto 0);
   Y_1_c5 <= '0' & Y(2 downto 0);
   S_1_c6 <= X_1_c6 + Y_1_c6 + Cin_1_c6;
   R_1_c6 <= S_1_c6(2 downto 0);
   Cin_2_c6 <= S_1_c6(3);
   X_2_c5 <= '0' & X(5 downto 3);
   Y_2_c5 <= '0' & Y(5 downto 3);
   S_2_c7 <= X_2_c7 + Y_2_c7 + Cin_2_c7;
   R_2_c7 <= S_2_c7(2 downto 0);
   Cin_3_c7 <= S_2_c7(3);
   X_3_c5 <= '0' & X(8 downto 6);
   Y_3_c5 <= '0' & Y(8 downto 6);
   S_3_c8 <= X_3_c8 + Y_3_c8 + Cin_3_c8;
   R_3_c8 <= S_3_c8(2 downto 0);
   Cin_4_c8 <= S_3_c8(3);
   X_4_c5 <= '0' & X(11 downto 9);
   Y_4_c5 <= '0' & Y(11 downto 9);
   S_4_c9 <= X_4_c9 + Y_4_c9 + Cin_4_c9;
   R_4_c9 <= S_4_c9(2 downto 0);
   Cin_5_c9 <= S_4_c9(3);
   X_5_c5 <= '0' & X(12 downto 12);
   Y_5_c5 <= '0' & Y(12 downto 12);
   S_5_c10 <= X_5_c10 + Y_5_c10 + Cin_5_c10;
   R_5_c10 <= S_5_c10(0 downto 0);
   R <= R_5_c10 & R_4_c10 & R_3_c10 & R_2_c10 & R_1_c10 ;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq800_uid8
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq800_uid8 is
    port (clk, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10 : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          R : out  std_logic_vector(7 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq800_uid8 is
   component FixRealKCM_Freq800_uid8_T0_Freq800_uid11 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(11 downto 0)   );
   end component;

   component FixRealKCM_Freq800_uid8_T1_Freq800_uid14 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(6 downto 0)   );
   end component;

   component IntAdder_13_Freq800_uid18 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10 : in std_logic;
             X : in  std_logic_vector(12 downto 0);
             Y : in  std_logic_vector(12 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(12 downto 0)   );
   end component;

signal FixRealKCM_Freq800_uid8_A0_c4 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq800_uid8_T0_c5 :  std_logic_vector(11 downto 0);
signal FixRealKCM_Freq800_uid8_T0_copy12_c4, FixRealKCM_Freq800_uid8_T0_copy12_c5 :  std_logic_vector(11 downto 0);
signal bh9_w0_0_c5 :  std_logic;
signal bh9_w1_0_c5 :  std_logic;
signal bh9_w2_0_c5 :  std_logic;
signal bh9_w3_0_c5 :  std_logic;
signal bh9_w4_0_c5 :  std_logic;
signal bh9_w5_0_c5 :  std_logic;
signal bh9_w6_0_c5 :  std_logic;
signal bh9_w7_0_c5 :  std_logic;
signal bh9_w8_0_c5 :  std_logic;
signal bh9_w9_0_c5 :  std_logic;
signal bh9_w10_0_c5 :  std_logic;
signal bh9_w11_0_c5 :  std_logic;
signal FixRealKCM_Freq800_uid8_A1_c4 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq800_uid8_T1_c5 :  std_logic_vector(6 downto 0);
signal FixRealKCM_Freq800_uid8_T1_copy15_c4, FixRealKCM_Freq800_uid8_T1_copy15_c5 :  std_logic_vector(6 downto 0);
signal bh9_w0_1_c5 :  std_logic;
signal bh9_w1_1_c5 :  std_logic;
signal bh9_w2_1_c5 :  std_logic;
signal bh9_w3_1_c5 :  std_logic;
signal bh9_w4_1_c5 :  std_logic;
signal bh9_w5_1_c5 :  std_logic;
signal bh9_w6_1_c5 :  std_logic;
signal bitheapFinalAdd_bh9_In0_c5 :  std_logic_vector(12 downto 0);
signal bitheapFinalAdd_bh9_In1_c5 :  std_logic_vector(12 downto 0);
signal bitheapFinalAdd_bh9_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh9_Out_c10 :  std_logic_vector(12 downto 0);
signal bitheapResult_bh9_c10 :  std_logic_vector(11 downto 0);
signal OutRes_c10 :  std_logic_vector(11 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_5 = '1' then
               FixRealKCM_Freq800_uid8_T0_copy12_c5 <= FixRealKCM_Freq800_uid8_T0_copy12_c4;
               FixRealKCM_Freq800_uid8_T1_copy15_c5 <= FixRealKCM_Freq800_uid8_T1_copy15_c4;
            end if;
            if ce_6 = '1' then
            end if;
            if ce_7 = '1' then
            end if;
            if ce_8 = '1' then
            end if;
            if ce_9 = '1' then
            end if;
            if ce_10 = '1' then
            end if;
         end if;
      end process;
-- This operator multiplies by 1/log(2)
   FixRealKCM_Freq800_uid8_A0_c4 <= X(9 downto 5);-- input address  m=6  l=2
   FixRealKCM_Freq800_uid8_Table0: FixRealKCM_Freq800_uid8_T0_Freq800_uid11
      port map ( X => FixRealKCM_Freq800_uid8_A0_c4,
                 Y => FixRealKCM_Freq800_uid8_T0_copy12_c4);
   FixRealKCM_Freq800_uid8_T0_c5 <= FixRealKCM_Freq800_uid8_T0_copy12_c5; -- output copy to hold a pipeline register if needed
   bh9_w0_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(0);
   bh9_w1_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(1);
   bh9_w2_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(2);
   bh9_w3_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(3);
   bh9_w4_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(4);
   bh9_w5_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(5);
   bh9_w6_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(6);
   bh9_w7_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(7);
   bh9_w8_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(8);
   bh9_w9_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(9);
   bh9_w10_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(10);
   bh9_w11_0_c5 <= FixRealKCM_Freq800_uid8_T0_c5(11);
   FixRealKCM_Freq800_uid8_A1_c4 <= X(4 downto 0);-- input address  m=1  l=-3
   FixRealKCM_Freq800_uid8_Table1: FixRealKCM_Freq800_uid8_T1_Freq800_uid14
      port map ( X => FixRealKCM_Freq800_uid8_A1_c4,
                 Y => FixRealKCM_Freq800_uid8_T1_copy15_c4);
   FixRealKCM_Freq800_uid8_T1_c5 <= FixRealKCM_Freq800_uid8_T1_copy15_c5; -- output copy to hold a pipeline register if needed
   bh9_w0_1_c5 <= FixRealKCM_Freq800_uid8_T1_c5(0);
   bh9_w1_1_c5 <= FixRealKCM_Freq800_uid8_T1_c5(1);
   bh9_w2_1_c5 <= FixRealKCM_Freq800_uid8_T1_c5(2);
   bh9_w3_1_c5 <= FixRealKCM_Freq800_uid8_T1_c5(3);
   bh9_w4_1_c5 <= FixRealKCM_Freq800_uid8_T1_c5(4);
   bh9_w5_1_c5 <= FixRealKCM_Freq800_uid8_T1_c5(5);
   bh9_w6_1_c5 <= FixRealKCM_Freq800_uid8_T1_c5(6);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh9_In0_c5 <= "0" & bh9_w11_0_c5 & bh9_w10_0_c5 & bh9_w9_0_c5 & bh9_w8_0_c5 & bh9_w7_0_c5 & bh9_w6_1_c5 & bh9_w5_1_c5 & bh9_w4_1_c5 & bh9_w3_1_c5 & bh9_w2_1_c5 & bh9_w1_1_c5 & bh9_w0_1_c5;
   bitheapFinalAdd_bh9_In1_c5 <= "0" & "0" & "0" & "0" & "0" & "0" & bh9_w6_0_c5 & bh9_w5_0_c5 & bh9_w4_0_c5 & bh9_w3_0_c5 & bh9_w2_0_c5 & bh9_w1_0_c5 & bh9_w0_0_c5;
   bitheapFinalAdd_bh9_Cin_c0 <= '0';

   bitheapFinalAdd_bh9: IntAdder_13_Freq800_uid18
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 Cin => bitheapFinalAdd_bh9_Cin_c0,
                 X => bitheapFinalAdd_bh9_In0_c5,
                 Y => bitheapFinalAdd_bh9_In1_c5,
                 R => bitheapFinalAdd_bh9_Out_c10);
   bitheapResult_bh9_c10 <= bitheapFinalAdd_bh9_Out_c10(11 downto 0);
   OutRes_c10 <= bitheapResult_bh9_c10(11 downto 0);
   R <= OutRes_c10(11 downto 4);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_36_Freq800_uid30
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 23 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_36_Freq800_uid30 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23 : in std_logic;
          X : in  std_logic_vector(35 downto 0);
          Y : in  std_logic_vector(35 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(35 downto 0)   );
end entity;

architecture arch of IntAdder_36_Freq800_uid30 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3, Cin_0_c4, Cin_0_c5, Cin_0_c6, Cin_0_c7, Cin_0_c8, Cin_0_c9, Cin_0_c10, Cin_0_c11 :  std_logic;
signal X_0_c10, X_0_c11 :  std_logic_vector(3 downto 0);
signal Y_0_c10, Y_0_c11 :  std_logic_vector(3 downto 0);
signal S_0_c11 :  std_logic_vector(3 downto 0);
signal R_0_c11, R_0_c12, R_0_c13, R_0_c14, R_0_c15, R_0_c16, R_0_c17, R_0_c18, R_0_c19, R_0_c20, R_0_c21, R_0_c22, R_0_c23 :  std_logic_vector(2 downto 0);
signal Cin_1_c11, Cin_1_c12 :  std_logic;
signal X_1_c10, X_1_c11, X_1_c12 :  std_logic_vector(3 downto 0);
signal Y_1_c10, Y_1_c11, Y_1_c12 :  std_logic_vector(3 downto 0);
signal S_1_c12 :  std_logic_vector(3 downto 0);
signal R_1_c12, R_1_c13, R_1_c14, R_1_c15, R_1_c16, R_1_c17, R_1_c18, R_1_c19, R_1_c20, R_1_c21, R_1_c22, R_1_c23 :  std_logic_vector(2 downto 0);
signal Cin_2_c12, Cin_2_c13 :  std_logic;
signal X_2_c10, X_2_c11, X_2_c12, X_2_c13 :  std_logic_vector(3 downto 0);
signal Y_2_c10, Y_2_c11, Y_2_c12, Y_2_c13 :  std_logic_vector(3 downto 0);
signal S_2_c13 :  std_logic_vector(3 downto 0);
signal R_2_c13, R_2_c14, R_2_c15, R_2_c16, R_2_c17, R_2_c18, R_2_c19, R_2_c20, R_2_c21, R_2_c22, R_2_c23 :  std_logic_vector(2 downto 0);
signal Cin_3_c13, Cin_3_c14 :  std_logic;
signal X_3_c10, X_3_c11, X_3_c12, X_3_c13, X_3_c14 :  std_logic_vector(3 downto 0);
signal Y_3_c10, Y_3_c11, Y_3_c12, Y_3_c13, Y_3_c14 :  std_logic_vector(3 downto 0);
signal S_3_c14 :  std_logic_vector(3 downto 0);
signal R_3_c14, R_3_c15, R_3_c16, R_3_c17, R_3_c18, R_3_c19, R_3_c20, R_3_c21, R_3_c22, R_3_c23 :  std_logic_vector(2 downto 0);
signal Cin_4_c14, Cin_4_c15 :  std_logic;
signal X_4_c10, X_4_c11, X_4_c12, X_4_c13, X_4_c14, X_4_c15 :  std_logic_vector(3 downto 0);
signal Y_4_c10, Y_4_c11, Y_4_c12, Y_4_c13, Y_4_c14, Y_4_c15 :  std_logic_vector(3 downto 0);
signal S_4_c15 :  std_logic_vector(3 downto 0);
signal R_4_c15, R_4_c16, R_4_c17, R_4_c18, R_4_c19, R_4_c20, R_4_c21, R_4_c22, R_4_c23 :  std_logic_vector(2 downto 0);
signal Cin_5_c15, Cin_5_c16, Cin_5_c17 :  std_logic;
signal X_5_c10, X_5_c11, X_5_c12, X_5_c13, X_5_c14, X_5_c15, X_5_c16, X_5_c17 :  std_logic_vector(3 downto 0);
signal Y_5_c10, Y_5_c11, Y_5_c12, Y_5_c13, Y_5_c14, Y_5_c15, Y_5_c16, Y_5_c17 :  std_logic_vector(3 downto 0);
signal S_5_c17 :  std_logic_vector(3 downto 0);
signal R_5_c17, R_5_c18, R_5_c19, R_5_c20, R_5_c21, R_5_c22, R_5_c23 :  std_logic_vector(2 downto 0);
signal Cin_6_c17, Cin_6_c18 :  std_logic;
signal X_6_c10, X_6_c11, X_6_c12, X_6_c13, X_6_c14, X_6_c15, X_6_c16, X_6_c17, X_6_c18 :  std_logic_vector(3 downto 0);
signal Y_6_c10, Y_6_c11, Y_6_c12, Y_6_c13, Y_6_c14, Y_6_c15, Y_6_c16, Y_6_c17, Y_6_c18 :  std_logic_vector(3 downto 0);
signal S_6_c18 :  std_logic_vector(3 downto 0);
signal R_6_c18, R_6_c19, R_6_c20, R_6_c21, R_6_c22, R_6_c23 :  std_logic_vector(2 downto 0);
signal Cin_7_c18, Cin_7_c19 :  std_logic;
signal X_7_c10, X_7_c11, X_7_c12, X_7_c13, X_7_c14, X_7_c15, X_7_c16, X_7_c17, X_7_c18, X_7_c19 :  std_logic_vector(3 downto 0);
signal Y_7_c10, Y_7_c11, Y_7_c12, Y_7_c13, Y_7_c14, Y_7_c15, Y_7_c16, Y_7_c17, Y_7_c18, Y_7_c19 :  std_logic_vector(3 downto 0);
signal S_7_c19 :  std_logic_vector(3 downto 0);
signal R_7_c19, R_7_c20, R_7_c21, R_7_c22, R_7_c23 :  std_logic_vector(2 downto 0);
signal Cin_8_c19, Cin_8_c20 :  std_logic;
signal X_8_c10, X_8_c11, X_8_c12, X_8_c13, X_8_c14, X_8_c15, X_8_c16, X_8_c17, X_8_c18, X_8_c19, X_8_c20 :  std_logic_vector(3 downto 0);
signal Y_8_c10, Y_8_c11, Y_8_c12, Y_8_c13, Y_8_c14, Y_8_c15, Y_8_c16, Y_8_c17, Y_8_c18, Y_8_c19, Y_8_c20 :  std_logic_vector(3 downto 0);
signal S_8_c20 :  std_logic_vector(3 downto 0);
signal R_8_c20, R_8_c21, R_8_c22, R_8_c23 :  std_logic_vector(2 downto 0);
signal Cin_9_c20, Cin_9_c21 :  std_logic;
signal X_9_c10, X_9_c11, X_9_c12, X_9_c13, X_9_c14, X_9_c15, X_9_c16, X_9_c17, X_9_c18, X_9_c19, X_9_c20, X_9_c21 :  std_logic_vector(3 downto 0);
signal Y_9_c10, Y_9_c11, Y_9_c12, Y_9_c13, Y_9_c14, Y_9_c15, Y_9_c16, Y_9_c17, Y_9_c18, Y_9_c19, Y_9_c20, Y_9_c21 :  std_logic_vector(3 downto 0);
signal S_9_c21 :  std_logic_vector(3 downto 0);
signal R_9_c21, R_9_c22, R_9_c23 :  std_logic_vector(2 downto 0);
signal Cin_10_c21, Cin_10_c22 :  std_logic;
signal X_10_c10, X_10_c11, X_10_c12, X_10_c13, X_10_c14, X_10_c15, X_10_c16, X_10_c17, X_10_c18, X_10_c19, X_10_c20, X_10_c21, X_10_c22 :  std_logic_vector(3 downto 0);
signal Y_10_c10, Y_10_c11, Y_10_c12, Y_10_c13, Y_10_c14, Y_10_c15, Y_10_c16, Y_10_c17, Y_10_c18, Y_10_c19, Y_10_c20, Y_10_c21, Y_10_c22 :  std_logic_vector(3 downto 0);
signal S_10_c22 :  std_logic_vector(3 downto 0);
signal R_10_c22, R_10_c23 :  std_logic_vector(2 downto 0);
signal Cin_11_c22, Cin_11_c23 :  std_logic;
signal X_11_c10, X_11_c11, X_11_c12, X_11_c13, X_11_c14, X_11_c15, X_11_c16, X_11_c17, X_11_c18, X_11_c19, X_11_c20, X_11_c21, X_11_c22, X_11_c23 :  std_logic_vector(3 downto 0);
signal Y_11_c10, Y_11_c11, Y_11_c12, Y_11_c13, Y_11_c14, Y_11_c15, Y_11_c16, Y_11_c17, Y_11_c18, Y_11_c19, Y_11_c20, Y_11_c21, Y_11_c22, Y_11_c23 :  std_logic_vector(3 downto 0);
signal S_11_c23 :  std_logic_vector(3 downto 0);
signal R_11_c23 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
            end if;
            if ce_4 = '1' then
               Cin_0_c4 <= Cin_0_c3;
            end if;
            if ce_5 = '1' then
               Cin_0_c5 <= Cin_0_c4;
            end if;
            if ce_6 = '1' then
               Cin_0_c6 <= Cin_0_c5;
            end if;
            if ce_7 = '1' then
               Cin_0_c7 <= Cin_0_c6;
            end if;
            if ce_8 = '1' then
               Cin_0_c8 <= Cin_0_c7;
            end if;
            if ce_9 = '1' then
               Cin_0_c9 <= Cin_0_c8;
            end if;
            if ce_10 = '1' then
               Cin_0_c10 <= Cin_0_c9;
            end if;
            if ce_11 = '1' then
               Cin_0_c11 <= Cin_0_c10;
               X_0_c11 <= X_0_c10;
               Y_0_c11 <= Y_0_c10;
               X_1_c11 <= X_1_c10;
               Y_1_c11 <= Y_1_c10;
               X_2_c11 <= X_2_c10;
               Y_2_c11 <= Y_2_c10;
               X_3_c11 <= X_3_c10;
               Y_3_c11 <= Y_3_c10;
               X_4_c11 <= X_4_c10;
               Y_4_c11 <= Y_4_c10;
               X_5_c11 <= X_5_c10;
               Y_5_c11 <= Y_5_c10;
               X_6_c11 <= X_6_c10;
               Y_6_c11 <= Y_6_c10;
               X_7_c11 <= X_7_c10;
               Y_7_c11 <= Y_7_c10;
               X_8_c11 <= X_8_c10;
               Y_8_c11 <= Y_8_c10;
               X_9_c11 <= X_9_c10;
               Y_9_c11 <= Y_9_c10;
               X_10_c11 <= X_10_c10;
               Y_10_c11 <= Y_10_c10;
               X_11_c11 <= X_11_c10;
               Y_11_c11 <= Y_11_c10;
            end if;
            if ce_12 = '1' then
               R_0_c12 <= R_0_c11;
               Cin_1_c12 <= Cin_1_c11;
               X_1_c12 <= X_1_c11;
               Y_1_c12 <= Y_1_c11;
               X_2_c12 <= X_2_c11;
               Y_2_c12 <= Y_2_c11;
               X_3_c12 <= X_3_c11;
               Y_3_c12 <= Y_3_c11;
               X_4_c12 <= X_4_c11;
               Y_4_c12 <= Y_4_c11;
               X_5_c12 <= X_5_c11;
               Y_5_c12 <= Y_5_c11;
               X_6_c12 <= X_6_c11;
               Y_6_c12 <= Y_6_c11;
               X_7_c12 <= X_7_c11;
               Y_7_c12 <= Y_7_c11;
               X_8_c12 <= X_8_c11;
               Y_8_c12 <= Y_8_c11;
               X_9_c12 <= X_9_c11;
               Y_9_c12 <= Y_9_c11;
               X_10_c12 <= X_10_c11;
               Y_10_c12 <= Y_10_c11;
               X_11_c12 <= X_11_c11;
               Y_11_c12 <= Y_11_c11;
            end if;
            if ce_13 = '1' then
               R_0_c13 <= R_0_c12;
               R_1_c13 <= R_1_c12;
               Cin_2_c13 <= Cin_2_c12;
               X_2_c13 <= X_2_c12;
               Y_2_c13 <= Y_2_c12;
               X_3_c13 <= X_3_c12;
               Y_3_c13 <= Y_3_c12;
               X_4_c13 <= X_4_c12;
               Y_4_c13 <= Y_4_c12;
               X_5_c13 <= X_5_c12;
               Y_5_c13 <= Y_5_c12;
               X_6_c13 <= X_6_c12;
               Y_6_c13 <= Y_6_c12;
               X_7_c13 <= X_7_c12;
               Y_7_c13 <= Y_7_c12;
               X_8_c13 <= X_8_c12;
               Y_8_c13 <= Y_8_c12;
               X_9_c13 <= X_9_c12;
               Y_9_c13 <= Y_9_c12;
               X_10_c13 <= X_10_c12;
               Y_10_c13 <= Y_10_c12;
               X_11_c13 <= X_11_c12;
               Y_11_c13 <= Y_11_c12;
            end if;
            if ce_14 = '1' then
               R_0_c14 <= R_0_c13;
               R_1_c14 <= R_1_c13;
               R_2_c14 <= R_2_c13;
               Cin_3_c14 <= Cin_3_c13;
               X_3_c14 <= X_3_c13;
               Y_3_c14 <= Y_3_c13;
               X_4_c14 <= X_4_c13;
               Y_4_c14 <= Y_4_c13;
               X_5_c14 <= X_5_c13;
               Y_5_c14 <= Y_5_c13;
               X_6_c14 <= X_6_c13;
               Y_6_c14 <= Y_6_c13;
               X_7_c14 <= X_7_c13;
               Y_7_c14 <= Y_7_c13;
               X_8_c14 <= X_8_c13;
               Y_8_c14 <= Y_8_c13;
               X_9_c14 <= X_9_c13;
               Y_9_c14 <= Y_9_c13;
               X_10_c14 <= X_10_c13;
               Y_10_c14 <= Y_10_c13;
               X_11_c14 <= X_11_c13;
               Y_11_c14 <= Y_11_c13;
            end if;
            if ce_15 = '1' then
               R_0_c15 <= R_0_c14;
               R_1_c15 <= R_1_c14;
               R_2_c15 <= R_2_c14;
               R_3_c15 <= R_3_c14;
               Cin_4_c15 <= Cin_4_c14;
               X_4_c15 <= X_4_c14;
               Y_4_c15 <= Y_4_c14;
               X_5_c15 <= X_5_c14;
               Y_5_c15 <= Y_5_c14;
               X_6_c15 <= X_6_c14;
               Y_6_c15 <= Y_6_c14;
               X_7_c15 <= X_7_c14;
               Y_7_c15 <= Y_7_c14;
               X_8_c15 <= X_8_c14;
               Y_8_c15 <= Y_8_c14;
               X_9_c15 <= X_9_c14;
               Y_9_c15 <= Y_9_c14;
               X_10_c15 <= X_10_c14;
               Y_10_c15 <= Y_10_c14;
               X_11_c15 <= X_11_c14;
               Y_11_c15 <= Y_11_c14;
            end if;
            if ce_16 = '1' then
               R_0_c16 <= R_0_c15;
               R_1_c16 <= R_1_c15;
               R_2_c16 <= R_2_c15;
               R_3_c16 <= R_3_c15;
               R_4_c16 <= R_4_c15;
               Cin_5_c16 <= Cin_5_c15;
               X_5_c16 <= X_5_c15;
               Y_5_c16 <= Y_5_c15;
               X_6_c16 <= X_6_c15;
               Y_6_c16 <= Y_6_c15;
               X_7_c16 <= X_7_c15;
               Y_7_c16 <= Y_7_c15;
               X_8_c16 <= X_8_c15;
               Y_8_c16 <= Y_8_c15;
               X_9_c16 <= X_9_c15;
               Y_9_c16 <= Y_9_c15;
               X_10_c16 <= X_10_c15;
               Y_10_c16 <= Y_10_c15;
               X_11_c16 <= X_11_c15;
               Y_11_c16 <= Y_11_c15;
            end if;
            if ce_17 = '1' then
               R_0_c17 <= R_0_c16;
               R_1_c17 <= R_1_c16;
               R_2_c17 <= R_2_c16;
               R_3_c17 <= R_3_c16;
               R_4_c17 <= R_4_c16;
               Cin_5_c17 <= Cin_5_c16;
               X_5_c17 <= X_5_c16;
               Y_5_c17 <= Y_5_c16;
               X_6_c17 <= X_6_c16;
               Y_6_c17 <= Y_6_c16;
               X_7_c17 <= X_7_c16;
               Y_7_c17 <= Y_7_c16;
               X_8_c17 <= X_8_c16;
               Y_8_c17 <= Y_8_c16;
               X_9_c17 <= X_9_c16;
               Y_9_c17 <= Y_9_c16;
               X_10_c17 <= X_10_c16;
               Y_10_c17 <= Y_10_c16;
               X_11_c17 <= X_11_c16;
               Y_11_c17 <= Y_11_c16;
            end if;
            if ce_18 = '1' then
               R_0_c18 <= R_0_c17;
               R_1_c18 <= R_1_c17;
               R_2_c18 <= R_2_c17;
               R_3_c18 <= R_3_c17;
               R_4_c18 <= R_4_c17;
               R_5_c18 <= R_5_c17;
               Cin_6_c18 <= Cin_6_c17;
               X_6_c18 <= X_6_c17;
               Y_6_c18 <= Y_6_c17;
               X_7_c18 <= X_7_c17;
               Y_7_c18 <= Y_7_c17;
               X_8_c18 <= X_8_c17;
               Y_8_c18 <= Y_8_c17;
               X_9_c18 <= X_9_c17;
               Y_9_c18 <= Y_9_c17;
               X_10_c18 <= X_10_c17;
               Y_10_c18 <= Y_10_c17;
               X_11_c18 <= X_11_c17;
               Y_11_c18 <= Y_11_c17;
            end if;
            if ce_19 = '1' then
               R_0_c19 <= R_0_c18;
               R_1_c19 <= R_1_c18;
               R_2_c19 <= R_2_c18;
               R_3_c19 <= R_3_c18;
               R_4_c19 <= R_4_c18;
               R_5_c19 <= R_5_c18;
               R_6_c19 <= R_6_c18;
               Cin_7_c19 <= Cin_7_c18;
               X_7_c19 <= X_7_c18;
               Y_7_c19 <= Y_7_c18;
               X_8_c19 <= X_8_c18;
               Y_8_c19 <= Y_8_c18;
               X_9_c19 <= X_9_c18;
               Y_9_c19 <= Y_9_c18;
               X_10_c19 <= X_10_c18;
               Y_10_c19 <= Y_10_c18;
               X_11_c19 <= X_11_c18;
               Y_11_c19 <= Y_11_c18;
            end if;
            if ce_20 = '1' then
               R_0_c20 <= R_0_c19;
               R_1_c20 <= R_1_c19;
               R_2_c20 <= R_2_c19;
               R_3_c20 <= R_3_c19;
               R_4_c20 <= R_4_c19;
               R_5_c20 <= R_5_c19;
               R_6_c20 <= R_6_c19;
               R_7_c20 <= R_7_c19;
               Cin_8_c20 <= Cin_8_c19;
               X_8_c20 <= X_8_c19;
               Y_8_c20 <= Y_8_c19;
               X_9_c20 <= X_9_c19;
               Y_9_c20 <= Y_9_c19;
               X_10_c20 <= X_10_c19;
               Y_10_c20 <= Y_10_c19;
               X_11_c20 <= X_11_c19;
               Y_11_c20 <= Y_11_c19;
            end if;
            if ce_21 = '1' then
               R_0_c21 <= R_0_c20;
               R_1_c21 <= R_1_c20;
               R_2_c21 <= R_2_c20;
               R_3_c21 <= R_3_c20;
               R_4_c21 <= R_4_c20;
               R_5_c21 <= R_5_c20;
               R_6_c21 <= R_6_c20;
               R_7_c21 <= R_7_c20;
               R_8_c21 <= R_8_c20;
               Cin_9_c21 <= Cin_9_c20;
               X_9_c21 <= X_9_c20;
               Y_9_c21 <= Y_9_c20;
               X_10_c21 <= X_10_c20;
               Y_10_c21 <= Y_10_c20;
               X_11_c21 <= X_11_c20;
               Y_11_c21 <= Y_11_c20;
            end if;
            if ce_22 = '1' then
               R_0_c22 <= R_0_c21;
               R_1_c22 <= R_1_c21;
               R_2_c22 <= R_2_c21;
               R_3_c22 <= R_3_c21;
               R_4_c22 <= R_4_c21;
               R_5_c22 <= R_5_c21;
               R_6_c22 <= R_6_c21;
               R_7_c22 <= R_7_c21;
               R_8_c22 <= R_8_c21;
               R_9_c22 <= R_9_c21;
               Cin_10_c22 <= Cin_10_c21;
               X_10_c22 <= X_10_c21;
               Y_10_c22 <= Y_10_c21;
               X_11_c22 <= X_11_c21;
               Y_11_c22 <= Y_11_c21;
            end if;
            if ce_23 = '1' then
               R_0_c23 <= R_0_c22;
               R_1_c23 <= R_1_c22;
               R_2_c23 <= R_2_c22;
               R_3_c23 <= R_3_c22;
               R_4_c23 <= R_4_c22;
               R_5_c23 <= R_5_c22;
               R_6_c23 <= R_6_c22;
               R_7_c23 <= R_7_c22;
               R_8_c23 <= R_8_c22;
               R_9_c23 <= R_9_c22;
               R_10_c23 <= R_10_c22;
               Cin_11_c23 <= Cin_11_c22;
               X_11_c23 <= X_11_c22;
               Y_11_c23 <= Y_11_c22;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c10 <= '0' & X(2 downto 0);
   Y_0_c10 <= '0' & Y(2 downto 0);
   S_0_c11 <= X_0_c11 + Y_0_c11 + Cin_0_c11;
   R_0_c11 <= S_0_c11(2 downto 0);
   Cin_1_c11 <= S_0_c11(3);
   X_1_c10 <= '0' & X(5 downto 3);
   Y_1_c10 <= '0' & Y(5 downto 3);
   S_1_c12 <= X_1_c12 + Y_1_c12 + Cin_1_c12;
   R_1_c12 <= S_1_c12(2 downto 0);
   Cin_2_c12 <= S_1_c12(3);
   X_2_c10 <= '0' & X(8 downto 6);
   Y_2_c10 <= '0' & Y(8 downto 6);
   S_2_c13 <= X_2_c13 + Y_2_c13 + Cin_2_c13;
   R_2_c13 <= S_2_c13(2 downto 0);
   Cin_3_c13 <= S_2_c13(3);
   X_3_c10 <= '0' & X(11 downto 9);
   Y_3_c10 <= '0' & Y(11 downto 9);
   S_3_c14 <= X_3_c14 + Y_3_c14 + Cin_3_c14;
   R_3_c14 <= S_3_c14(2 downto 0);
   Cin_4_c14 <= S_3_c14(3);
   X_4_c10 <= '0' & X(14 downto 12);
   Y_4_c10 <= '0' & Y(14 downto 12);
   S_4_c15 <= X_4_c15 + Y_4_c15 + Cin_4_c15;
   R_4_c15 <= S_4_c15(2 downto 0);
   Cin_5_c15 <= S_4_c15(3);
   X_5_c10 <= '0' & X(17 downto 15);
   Y_5_c10 <= '0' & Y(17 downto 15);
   S_5_c17 <= X_5_c17 + Y_5_c17 + Cin_5_c17;
   R_5_c17 <= S_5_c17(2 downto 0);
   Cin_6_c17 <= S_5_c17(3);
   X_6_c10 <= '0' & X(20 downto 18);
   Y_6_c10 <= '0' & Y(20 downto 18);
   S_6_c18 <= X_6_c18 + Y_6_c18 + Cin_6_c18;
   R_6_c18 <= S_6_c18(2 downto 0);
   Cin_7_c18 <= S_6_c18(3);
   X_7_c10 <= '0' & X(23 downto 21);
   Y_7_c10 <= '0' & Y(23 downto 21);
   S_7_c19 <= X_7_c19 + Y_7_c19 + Cin_7_c19;
   R_7_c19 <= S_7_c19(2 downto 0);
   Cin_8_c19 <= S_7_c19(3);
   X_8_c10 <= '0' & X(26 downto 24);
   Y_8_c10 <= '0' & Y(26 downto 24);
   S_8_c20 <= X_8_c20 + Y_8_c20 + Cin_8_c20;
   R_8_c20 <= S_8_c20(2 downto 0);
   Cin_9_c20 <= S_8_c20(3);
   X_9_c10 <= '0' & X(29 downto 27);
   Y_9_c10 <= '0' & Y(29 downto 27);
   S_9_c21 <= X_9_c21 + Y_9_c21 + Cin_9_c21;
   R_9_c21 <= S_9_c21(2 downto 0);
   Cin_10_c21 <= S_9_c21(3);
   X_10_c10 <= '0' & X(32 downto 30);
   Y_10_c10 <= '0' & Y(32 downto 30);
   S_10_c22 <= X_10_c22 + Y_10_c22 + Cin_10_c22;
   R_10_c22 <= S_10_c22(2 downto 0);
   Cin_11_c22 <= S_10_c22(3);
   X_11_c10 <= '0' & X(35 downto 33);
   Y_11_c10 <= '0' & Y(35 downto 33);
   S_11_c23 <= X_11_c23 + Y_11_c23 + Cin_11_c23;
   R_11_c23 <= S_11_c23(2 downto 0);
   R <= R_11_c23 & R_10_c23 & R_9_c23 & R_8_c23 & R_7_c23 & R_6_c23 & R_5_c23 & R_4_c23 & R_3_c23 & R_2_c23 & R_1_c23 & R_0_c23 ;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq800_uid20
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq800_uid20 is
    port (clk, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23 : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          R : out  std_logic_vector(34 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq800_uid20 is
   component FixRealKCM_Freq800_uid20_T0_Freq800_uid23 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(34 downto 0)   );
   end component;

   component FixRealKCM_Freq800_uid20_T1_Freq800_uid26 is
      port ( X : in  std_logic_vector(2 downto 0);
             Y : out  std_logic_vector(29 downto 0)   );
   end component;

   component IntAdder_36_Freq800_uid30 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23 : in std_logic;
             X : in  std_logic_vector(35 downto 0);
             Y : in  std_logic_vector(35 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(35 downto 0)   );
   end component;

signal FixRealKCM_Freq800_uid20_A0_c10 :  std_logic_vector(4 downto 0);
signal FixRealKCM_Freq800_uid20_T0_c10 :  std_logic_vector(34 downto 0);
signal FixRealKCM_Freq800_uid20_T0_copy24_c10 :  std_logic_vector(34 downto 0);
signal bh21_w0_0_c10 :  std_logic;
signal bh21_w1_0_c10 :  std_logic;
signal bh21_w2_0_c10 :  std_logic;
signal bh21_w3_0_c10 :  std_logic;
signal bh21_w4_0_c10 :  std_logic;
signal bh21_w5_0_c10 :  std_logic;
signal bh21_w6_0_c10 :  std_logic;
signal bh21_w7_0_c10 :  std_logic;
signal bh21_w8_0_c10 :  std_logic;
signal bh21_w9_0_c10 :  std_logic;
signal bh21_w10_0_c10 :  std_logic;
signal bh21_w11_0_c10 :  std_logic;
signal bh21_w12_0_c10 :  std_logic;
signal bh21_w13_0_c10 :  std_logic;
signal bh21_w14_0_c10 :  std_logic;
signal bh21_w15_0_c10 :  std_logic;
signal bh21_w16_0_c10 :  std_logic;
signal bh21_w17_0_c10 :  std_logic;
signal bh21_w18_0_c10 :  std_logic;
signal bh21_w19_0_c10 :  std_logic;
signal bh21_w20_0_c10 :  std_logic;
signal bh21_w21_0_c10 :  std_logic;
signal bh21_w22_0_c10 :  std_logic;
signal bh21_w23_0_c10 :  std_logic;
signal bh21_w24_0_c10 :  std_logic;
signal bh21_w25_0_c10 :  std_logic;
signal bh21_w26_0_c10 :  std_logic;
signal bh21_w27_0_c10 :  std_logic;
signal bh21_w28_0_c10 :  std_logic;
signal bh21_w29_0_c10 :  std_logic;
signal bh21_w30_0_c10 :  std_logic;
signal bh21_w31_0_c10 :  std_logic;
signal bh21_w32_0_c10 :  std_logic;
signal bh21_w33_0_c10 :  std_logic;
signal bh21_w34_0_c10 :  std_logic;
signal FixRealKCM_Freq800_uid20_A1_c10 :  std_logic_vector(2 downto 0);
signal FixRealKCM_Freq800_uid20_T1_c10 :  std_logic_vector(29 downto 0);
signal FixRealKCM_Freq800_uid20_T1_copy27_c10 :  std_logic_vector(29 downto 0);
signal bh21_w0_1_c10 :  std_logic;
signal bh21_w1_1_c10 :  std_logic;
signal bh21_w2_1_c10 :  std_logic;
signal bh21_w3_1_c10 :  std_logic;
signal bh21_w4_1_c10 :  std_logic;
signal bh21_w5_1_c10 :  std_logic;
signal bh21_w6_1_c10 :  std_logic;
signal bh21_w7_1_c10 :  std_logic;
signal bh21_w8_1_c10 :  std_logic;
signal bh21_w9_1_c10 :  std_logic;
signal bh21_w10_1_c10 :  std_logic;
signal bh21_w11_1_c10 :  std_logic;
signal bh21_w12_1_c10 :  std_logic;
signal bh21_w13_1_c10 :  std_logic;
signal bh21_w14_1_c10 :  std_logic;
signal bh21_w15_1_c10 :  std_logic;
signal bh21_w16_1_c10 :  std_logic;
signal bh21_w17_1_c10 :  std_logic;
signal bh21_w18_1_c10 :  std_logic;
signal bh21_w19_1_c10 :  std_logic;
signal bh21_w20_1_c10 :  std_logic;
signal bh21_w21_1_c10 :  std_logic;
signal bh21_w22_1_c10 :  std_logic;
signal bh21_w23_1_c10 :  std_logic;
signal bh21_w24_1_c10 :  std_logic;
signal bh21_w25_1_c10 :  std_logic;
signal bh21_w26_1_c10 :  std_logic;
signal bh21_w27_1_c10 :  std_logic;
signal bh21_w28_1_c10 :  std_logic;
signal bh21_w29_1_c10 :  std_logic;
signal bitheapFinalAdd_bh21_In0_c10 :  std_logic_vector(35 downto 0);
signal bitheapFinalAdd_bh21_In1_c10 :  std_logic_vector(35 downto 0);
signal bitheapFinalAdd_bh21_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh21_Out_c23 :  std_logic_vector(35 downto 0);
signal bitheapResult_bh21_c23 :  std_logic_vector(34 downto 0);
signal OutRes_c23 :  std_logic_vector(34 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_11 = '1' then
            end if;
            if ce_12 = '1' then
            end if;
            if ce_13 = '1' then
            end if;
            if ce_14 = '1' then
            end if;
            if ce_15 = '1' then
            end if;
            if ce_16 = '1' then
            end if;
            if ce_17 = '1' then
            end if;
            if ce_18 = '1' then
            end if;
            if ce_19 = '1' then
            end if;
            if ce_20 = '1' then
            end if;
            if ce_21 = '1' then
            end if;
            if ce_22 = '1' then
            end if;
            if ce_23 = '1' then
            end if;
         end if;
      end process;
-- This operator multiplies by log(2)
   FixRealKCM_Freq800_uid20_A0_c10 <= X(7 downto 3);-- input address  m=7  l=3
   FixRealKCM_Freq800_uid20_Table0: FixRealKCM_Freq800_uid20_T0_Freq800_uid23
      port map ( X => FixRealKCM_Freq800_uid20_A0_c10,
                 Y => FixRealKCM_Freq800_uid20_T0_copy24_c10);
   FixRealKCM_Freq800_uid20_T0_c10 <= FixRealKCM_Freq800_uid20_T0_copy24_c10; -- output copy to hold a pipeline register if needed
   bh21_w0_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(0);
   bh21_w1_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(1);
   bh21_w2_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(2);
   bh21_w3_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(3);
   bh21_w4_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(4);
   bh21_w5_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(5);
   bh21_w6_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(6);
   bh21_w7_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(7);
   bh21_w8_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(8);
   bh21_w9_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(9);
   bh21_w10_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(10);
   bh21_w11_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(11);
   bh21_w12_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(12);
   bh21_w13_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(13);
   bh21_w14_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(14);
   bh21_w15_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(15);
   bh21_w16_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(16);
   bh21_w17_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(17);
   bh21_w18_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(18);
   bh21_w19_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(19);
   bh21_w20_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(20);
   bh21_w21_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(21);
   bh21_w22_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(22);
   bh21_w23_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(23);
   bh21_w24_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(24);
   bh21_w25_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(25);
   bh21_w26_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(26);
   bh21_w27_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(27);
   bh21_w28_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(28);
   bh21_w29_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(29);
   bh21_w30_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(30);
   bh21_w31_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(31);
   bh21_w32_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(32);
   bh21_w33_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(33);
   bh21_w34_0_c10 <= FixRealKCM_Freq800_uid20_T0_c10(34);
   FixRealKCM_Freq800_uid20_A1_c10 <= X(2 downto 0);-- input address  m=2  l=0
   FixRealKCM_Freq800_uid20_Table1: FixRealKCM_Freq800_uid20_T1_Freq800_uid26
      port map ( X => FixRealKCM_Freq800_uid20_A1_c10,
                 Y => FixRealKCM_Freq800_uid20_T1_copy27_c10);
   FixRealKCM_Freq800_uid20_T1_c10 <= FixRealKCM_Freq800_uid20_T1_copy27_c10; -- output copy to hold a pipeline register if needed
   bh21_w0_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(0);
   bh21_w1_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(1);
   bh21_w2_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(2);
   bh21_w3_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(3);
   bh21_w4_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(4);
   bh21_w5_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(5);
   bh21_w6_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(6);
   bh21_w7_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(7);
   bh21_w8_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(8);
   bh21_w9_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(9);
   bh21_w10_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(10);
   bh21_w11_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(11);
   bh21_w12_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(12);
   bh21_w13_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(13);
   bh21_w14_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(14);
   bh21_w15_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(15);
   bh21_w16_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(16);
   bh21_w17_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(17);
   bh21_w18_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(18);
   bh21_w19_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(19);
   bh21_w20_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(20);
   bh21_w21_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(21);
   bh21_w22_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(22);
   bh21_w23_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(23);
   bh21_w24_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(24);
   bh21_w25_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(25);
   bh21_w26_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(26);
   bh21_w27_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(27);
   bh21_w28_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(28);
   bh21_w29_1_c10 <= FixRealKCM_Freq800_uid20_T1_c10(29);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   bitheapFinalAdd_bh21_In0_c10 <= "0" & bh21_w34_0_c10 & bh21_w33_0_c10 & bh21_w32_0_c10 & bh21_w31_0_c10 & bh21_w30_0_c10 & bh21_w29_0_c10 & bh21_w28_0_c10 & bh21_w27_0_c10 & bh21_w26_0_c10 & bh21_w25_0_c10 & bh21_w24_0_c10 & bh21_w23_0_c10 & bh21_w22_0_c10 & bh21_w21_0_c10 & bh21_w20_0_c10 & bh21_w19_0_c10 & bh21_w18_0_c10 & bh21_w17_0_c10 & bh21_w16_0_c10 & bh21_w15_0_c10 & bh21_w14_0_c10 & bh21_w13_0_c10 & bh21_w12_0_c10 & bh21_w11_0_c10 & bh21_w10_0_c10 & bh21_w9_0_c10 & bh21_w8_0_c10 & bh21_w7_0_c10 & bh21_w6_0_c10 & bh21_w5_0_c10 & bh21_w4_0_c10 & bh21_w3_0_c10 & bh21_w2_0_c10 & bh21_w1_0_c10 & bh21_w0_0_c10;
   bitheapFinalAdd_bh21_In1_c10 <= "0" & "0" & "0" & "0" & "0" & "0" & bh21_w29_1_c10 & bh21_w28_1_c10 & bh21_w27_1_c10 & bh21_w26_1_c10 & bh21_w25_1_c10 & bh21_w24_1_c10 & bh21_w23_1_c10 & bh21_w22_1_c10 & bh21_w21_1_c10 & bh21_w20_1_c10 & bh21_w19_1_c10 & bh21_w18_1_c10 & bh21_w17_1_c10 & bh21_w16_1_c10 & bh21_w15_1_c10 & bh21_w14_1_c10 & bh21_w13_1_c10 & bh21_w12_1_c10 & bh21_w11_1_c10 & bh21_w10_1_c10 & bh21_w9_1_c10 & bh21_w8_1_c10 & bh21_w7_1_c10 & bh21_w6_1_c10 & bh21_w5_1_c10 & bh21_w4_1_c10 & bh21_w3_1_c10 & bh21_w2_1_c10 & bh21_w1_1_c10 & bh21_w0_1_c10;
   bitheapFinalAdd_bh21_Cin_c0 <= '0';

   bitheapFinalAdd_bh21: IntAdder_36_Freq800_uid30
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 Cin => bitheapFinalAdd_bh21_Cin_c0,
                 X => bitheapFinalAdd_bh21_In0_c10,
                 Y => bitheapFinalAdd_bh21_In1_c10,
                 R => bitheapFinalAdd_bh21_Out_c23);
   bitheapResult_bh21_c23 <= bitheapFinalAdd_bh21_Out_c23(34 downto 0);
   OutRes_c23 <= bitheapResult_bh21_c23(34 downto 0);
   R <= OutRes_c23(34 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_27_Freq800_uid33
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 32 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_Freq800_uid33 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32 : in std_logic;
          X : in  std_logic_vector(26 downto 0);
          Y : in  std_logic_vector(26 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_Freq800_uid33 is
signal Cin_1_c0, Cin_1_c1, Cin_1_c2, Cin_1_c3, Cin_1_c4, Cin_1_c5, Cin_1_c6, Cin_1_c7, Cin_1_c8, Cin_1_c9, Cin_1_c10, Cin_1_c11, Cin_1_c12, Cin_1_c13, Cin_1_c14, Cin_1_c15, Cin_1_c16, Cin_1_c17, Cin_1_c18, Cin_1_c19, Cin_1_c20, Cin_1_c21, Cin_1_c22, Cin_1_c23, Cin_1_c24 :  std_logic;
signal X_1_c5, X_1_c6, X_1_c7, X_1_c8, X_1_c9, X_1_c10, X_1_c11, X_1_c12, X_1_c13, X_1_c14, X_1_c15, X_1_c16, X_1_c17, X_1_c18, X_1_c19, X_1_c20, X_1_c21, X_1_c22, X_1_c23, X_1_c24 :  std_logic_vector(3 downto 0);
signal Y_1_c23, Y_1_c24 :  std_logic_vector(3 downto 0);
signal S_1_c24 :  std_logic_vector(3 downto 0);
signal R_1_c24, R_1_c25, R_1_c26, R_1_c27, R_1_c28, R_1_c29, R_1_c30, R_1_c31, R_1_c32 :  std_logic_vector(2 downto 0);
signal Cin_2_c24, Cin_2_c25 :  std_logic;
signal X_2_c5, X_2_c6, X_2_c7, X_2_c8, X_2_c9, X_2_c10, X_2_c11, X_2_c12, X_2_c13, X_2_c14, X_2_c15, X_2_c16, X_2_c17, X_2_c18, X_2_c19, X_2_c20, X_2_c21, X_2_c22, X_2_c23, X_2_c24, X_2_c25 :  std_logic_vector(3 downto 0);
signal Y_2_c23, Y_2_c24, Y_2_c25 :  std_logic_vector(3 downto 0);
signal S_2_c25 :  std_logic_vector(3 downto 0);
signal R_2_c25, R_2_c26, R_2_c27, R_2_c28, R_2_c29, R_2_c30, R_2_c31, R_2_c32 :  std_logic_vector(2 downto 0);
signal Cin_3_c25, Cin_3_c26 :  std_logic;
signal X_3_c5, X_3_c6, X_3_c7, X_3_c8, X_3_c9, X_3_c10, X_3_c11, X_3_c12, X_3_c13, X_3_c14, X_3_c15, X_3_c16, X_3_c17, X_3_c18, X_3_c19, X_3_c20, X_3_c21, X_3_c22, X_3_c23, X_3_c24, X_3_c25, X_3_c26 :  std_logic_vector(3 downto 0);
signal Y_3_c23, Y_3_c24, Y_3_c25, Y_3_c26 :  std_logic_vector(3 downto 0);
signal S_3_c26 :  std_logic_vector(3 downto 0);
signal R_3_c26, R_3_c27, R_3_c28, R_3_c29, R_3_c30, R_3_c31, R_3_c32 :  std_logic_vector(2 downto 0);
signal Cin_4_c26, Cin_4_c27 :  std_logic;
signal X_4_c5, X_4_c6, X_4_c7, X_4_c8, X_4_c9, X_4_c10, X_4_c11, X_4_c12, X_4_c13, X_4_c14, X_4_c15, X_4_c16, X_4_c17, X_4_c18, X_4_c19, X_4_c20, X_4_c21, X_4_c22, X_4_c23, X_4_c24, X_4_c25, X_4_c26, X_4_c27 :  std_logic_vector(3 downto 0);
signal Y_4_c23, Y_4_c24, Y_4_c25, Y_4_c26, Y_4_c27 :  std_logic_vector(3 downto 0);
signal S_4_c27 :  std_logic_vector(3 downto 0);
signal R_4_c27, R_4_c28, R_4_c29, R_4_c30, R_4_c31, R_4_c32 :  std_logic_vector(2 downto 0);
signal Cin_5_c27, Cin_5_c28 :  std_logic;
signal X_5_c5, X_5_c6, X_5_c7, X_5_c8, X_5_c9, X_5_c10, X_5_c11, X_5_c12, X_5_c13, X_5_c14, X_5_c15, X_5_c16, X_5_c17, X_5_c18, X_5_c19, X_5_c20, X_5_c21, X_5_c22, X_5_c23, X_5_c24, X_5_c25, X_5_c26, X_5_c27, X_5_c28 :  std_logic_vector(3 downto 0);
signal Y_5_c23, Y_5_c24, Y_5_c25, Y_5_c26, Y_5_c27, Y_5_c28 :  std_logic_vector(3 downto 0);
signal S_5_c28 :  std_logic_vector(3 downto 0);
signal R_5_c28, R_5_c29, R_5_c30, R_5_c31, R_5_c32 :  std_logic_vector(2 downto 0);
signal Cin_6_c28, Cin_6_c29 :  std_logic;
signal X_6_c5, X_6_c6, X_6_c7, X_6_c8, X_6_c9, X_6_c10, X_6_c11, X_6_c12, X_6_c13, X_6_c14, X_6_c15, X_6_c16, X_6_c17, X_6_c18, X_6_c19, X_6_c20, X_6_c21, X_6_c22, X_6_c23, X_6_c24, X_6_c25, X_6_c26, X_6_c27, X_6_c28, X_6_c29 :  std_logic_vector(3 downto 0);
signal Y_6_c23, Y_6_c24, Y_6_c25, Y_6_c26, Y_6_c27, Y_6_c28, Y_6_c29 :  std_logic_vector(3 downto 0);
signal S_6_c29 :  std_logic_vector(3 downto 0);
signal R_6_c29, R_6_c30, R_6_c31, R_6_c32 :  std_logic_vector(2 downto 0);
signal Cin_7_c29, Cin_7_c30 :  std_logic;
signal X_7_c5, X_7_c6, X_7_c7, X_7_c8, X_7_c9, X_7_c10, X_7_c11, X_7_c12, X_7_c13, X_7_c14, X_7_c15, X_7_c16, X_7_c17, X_7_c18, X_7_c19, X_7_c20, X_7_c21, X_7_c22, X_7_c23, X_7_c24, X_7_c25, X_7_c26, X_7_c27, X_7_c28, X_7_c29, X_7_c30 :  std_logic_vector(3 downto 0);
signal Y_7_c23, Y_7_c24, Y_7_c25, Y_7_c26, Y_7_c27, Y_7_c28, Y_7_c29, Y_7_c30 :  std_logic_vector(3 downto 0);
signal S_7_c30 :  std_logic_vector(3 downto 0);
signal R_7_c30, R_7_c31, R_7_c32 :  std_logic_vector(2 downto 0);
signal Cin_8_c30, Cin_8_c31 :  std_logic;
signal X_8_c5, X_8_c6, X_8_c7, X_8_c8, X_8_c9, X_8_c10, X_8_c11, X_8_c12, X_8_c13, X_8_c14, X_8_c15, X_8_c16, X_8_c17, X_8_c18, X_8_c19, X_8_c20, X_8_c21, X_8_c22, X_8_c23, X_8_c24, X_8_c25, X_8_c26, X_8_c27, X_8_c28, X_8_c29, X_8_c30, X_8_c31 :  std_logic_vector(3 downto 0);
signal Y_8_c23, Y_8_c24, Y_8_c25, Y_8_c26, Y_8_c27, Y_8_c28, Y_8_c29, Y_8_c30, Y_8_c31 :  std_logic_vector(3 downto 0);
signal S_8_c31 :  std_logic_vector(3 downto 0);
signal R_8_c31, R_8_c32 :  std_logic_vector(2 downto 0);
signal Cin_9_c31, Cin_9_c32 :  std_logic;
signal X_9_c5, X_9_c6, X_9_c7, X_9_c8, X_9_c9, X_9_c10, X_9_c11, X_9_c12, X_9_c13, X_9_c14, X_9_c15, X_9_c16, X_9_c17, X_9_c18, X_9_c19, X_9_c20, X_9_c21, X_9_c22, X_9_c23, X_9_c24, X_9_c25, X_9_c26, X_9_c27, X_9_c28, X_9_c29, X_9_c30, X_9_c31, X_9_c32 :  std_logic_vector(3 downto 0);
signal Y_9_c23, Y_9_c24, Y_9_c25, Y_9_c26, Y_9_c27, Y_9_c28, Y_9_c29, Y_9_c30, Y_9_c31, Y_9_c32 :  std_logic_vector(3 downto 0);
signal S_9_c32 :  std_logic_vector(3 downto 0);
signal R_9_c32 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_1_c1 <= Cin_1_c0;
            end if;
            if ce_2 = '1' then
               Cin_1_c2 <= Cin_1_c1;
            end if;
            if ce_3 = '1' then
               Cin_1_c3 <= Cin_1_c2;
            end if;
            if ce_4 = '1' then
               Cin_1_c4 <= Cin_1_c3;
            end if;
            if ce_5 = '1' then
               Cin_1_c5 <= Cin_1_c4;
            end if;
            if ce_6 = '1' then
               Cin_1_c6 <= Cin_1_c5;
               X_1_c6 <= X_1_c5;
               X_2_c6 <= X_2_c5;
               X_3_c6 <= X_3_c5;
               X_4_c6 <= X_4_c5;
               X_5_c6 <= X_5_c5;
               X_6_c6 <= X_6_c5;
               X_7_c6 <= X_7_c5;
               X_8_c6 <= X_8_c5;
               X_9_c6 <= X_9_c5;
            end if;
            if ce_7 = '1' then
               Cin_1_c7 <= Cin_1_c6;
               X_1_c7 <= X_1_c6;
               X_2_c7 <= X_2_c6;
               X_3_c7 <= X_3_c6;
               X_4_c7 <= X_4_c6;
               X_5_c7 <= X_5_c6;
               X_6_c7 <= X_6_c6;
               X_7_c7 <= X_7_c6;
               X_8_c7 <= X_8_c6;
               X_9_c7 <= X_9_c6;
            end if;
            if ce_8 = '1' then
               Cin_1_c8 <= Cin_1_c7;
               X_1_c8 <= X_1_c7;
               X_2_c8 <= X_2_c7;
               X_3_c8 <= X_3_c7;
               X_4_c8 <= X_4_c7;
               X_5_c8 <= X_5_c7;
               X_6_c8 <= X_6_c7;
               X_7_c8 <= X_7_c7;
               X_8_c8 <= X_8_c7;
               X_9_c8 <= X_9_c7;
            end if;
            if ce_9 = '1' then
               Cin_1_c9 <= Cin_1_c8;
               X_1_c9 <= X_1_c8;
               X_2_c9 <= X_2_c8;
               X_3_c9 <= X_3_c8;
               X_4_c9 <= X_4_c8;
               X_5_c9 <= X_5_c8;
               X_6_c9 <= X_6_c8;
               X_7_c9 <= X_7_c8;
               X_8_c9 <= X_8_c8;
               X_9_c9 <= X_9_c8;
            end if;
            if ce_10 = '1' then
               Cin_1_c10 <= Cin_1_c9;
               X_1_c10 <= X_1_c9;
               X_2_c10 <= X_2_c9;
               X_3_c10 <= X_3_c9;
               X_4_c10 <= X_4_c9;
               X_5_c10 <= X_5_c9;
               X_6_c10 <= X_6_c9;
               X_7_c10 <= X_7_c9;
               X_8_c10 <= X_8_c9;
               X_9_c10 <= X_9_c9;
            end if;
            if ce_11 = '1' then
               Cin_1_c11 <= Cin_1_c10;
               X_1_c11 <= X_1_c10;
               X_2_c11 <= X_2_c10;
               X_3_c11 <= X_3_c10;
               X_4_c11 <= X_4_c10;
               X_5_c11 <= X_5_c10;
               X_6_c11 <= X_6_c10;
               X_7_c11 <= X_7_c10;
               X_8_c11 <= X_8_c10;
               X_9_c11 <= X_9_c10;
            end if;
            if ce_12 = '1' then
               Cin_1_c12 <= Cin_1_c11;
               X_1_c12 <= X_1_c11;
               X_2_c12 <= X_2_c11;
               X_3_c12 <= X_3_c11;
               X_4_c12 <= X_4_c11;
               X_5_c12 <= X_5_c11;
               X_6_c12 <= X_6_c11;
               X_7_c12 <= X_7_c11;
               X_8_c12 <= X_8_c11;
               X_9_c12 <= X_9_c11;
            end if;
            if ce_13 = '1' then
               Cin_1_c13 <= Cin_1_c12;
               X_1_c13 <= X_1_c12;
               X_2_c13 <= X_2_c12;
               X_3_c13 <= X_3_c12;
               X_4_c13 <= X_4_c12;
               X_5_c13 <= X_5_c12;
               X_6_c13 <= X_6_c12;
               X_7_c13 <= X_7_c12;
               X_8_c13 <= X_8_c12;
               X_9_c13 <= X_9_c12;
            end if;
            if ce_14 = '1' then
               Cin_1_c14 <= Cin_1_c13;
               X_1_c14 <= X_1_c13;
               X_2_c14 <= X_2_c13;
               X_3_c14 <= X_3_c13;
               X_4_c14 <= X_4_c13;
               X_5_c14 <= X_5_c13;
               X_6_c14 <= X_6_c13;
               X_7_c14 <= X_7_c13;
               X_8_c14 <= X_8_c13;
               X_9_c14 <= X_9_c13;
            end if;
            if ce_15 = '1' then
               Cin_1_c15 <= Cin_1_c14;
               X_1_c15 <= X_1_c14;
               X_2_c15 <= X_2_c14;
               X_3_c15 <= X_3_c14;
               X_4_c15 <= X_4_c14;
               X_5_c15 <= X_5_c14;
               X_6_c15 <= X_6_c14;
               X_7_c15 <= X_7_c14;
               X_8_c15 <= X_8_c14;
               X_9_c15 <= X_9_c14;
            end if;
            if ce_16 = '1' then
               Cin_1_c16 <= Cin_1_c15;
               X_1_c16 <= X_1_c15;
               X_2_c16 <= X_2_c15;
               X_3_c16 <= X_3_c15;
               X_4_c16 <= X_4_c15;
               X_5_c16 <= X_5_c15;
               X_6_c16 <= X_6_c15;
               X_7_c16 <= X_7_c15;
               X_8_c16 <= X_8_c15;
               X_9_c16 <= X_9_c15;
            end if;
            if ce_17 = '1' then
               Cin_1_c17 <= Cin_1_c16;
               X_1_c17 <= X_1_c16;
               X_2_c17 <= X_2_c16;
               X_3_c17 <= X_3_c16;
               X_4_c17 <= X_4_c16;
               X_5_c17 <= X_5_c16;
               X_6_c17 <= X_6_c16;
               X_7_c17 <= X_7_c16;
               X_8_c17 <= X_8_c16;
               X_9_c17 <= X_9_c16;
            end if;
            if ce_18 = '1' then
               Cin_1_c18 <= Cin_1_c17;
               X_1_c18 <= X_1_c17;
               X_2_c18 <= X_2_c17;
               X_3_c18 <= X_3_c17;
               X_4_c18 <= X_4_c17;
               X_5_c18 <= X_5_c17;
               X_6_c18 <= X_6_c17;
               X_7_c18 <= X_7_c17;
               X_8_c18 <= X_8_c17;
               X_9_c18 <= X_9_c17;
            end if;
            if ce_19 = '1' then
               Cin_1_c19 <= Cin_1_c18;
               X_1_c19 <= X_1_c18;
               X_2_c19 <= X_2_c18;
               X_3_c19 <= X_3_c18;
               X_4_c19 <= X_4_c18;
               X_5_c19 <= X_5_c18;
               X_6_c19 <= X_6_c18;
               X_7_c19 <= X_7_c18;
               X_8_c19 <= X_8_c18;
               X_9_c19 <= X_9_c18;
            end if;
            if ce_20 = '1' then
               Cin_1_c20 <= Cin_1_c19;
               X_1_c20 <= X_1_c19;
               X_2_c20 <= X_2_c19;
               X_3_c20 <= X_3_c19;
               X_4_c20 <= X_4_c19;
               X_5_c20 <= X_5_c19;
               X_6_c20 <= X_6_c19;
               X_7_c20 <= X_7_c19;
               X_8_c20 <= X_8_c19;
               X_9_c20 <= X_9_c19;
            end if;
            if ce_21 = '1' then
               Cin_1_c21 <= Cin_1_c20;
               X_1_c21 <= X_1_c20;
               X_2_c21 <= X_2_c20;
               X_3_c21 <= X_3_c20;
               X_4_c21 <= X_4_c20;
               X_5_c21 <= X_5_c20;
               X_6_c21 <= X_6_c20;
               X_7_c21 <= X_7_c20;
               X_8_c21 <= X_8_c20;
               X_9_c21 <= X_9_c20;
            end if;
            if ce_22 = '1' then
               Cin_1_c22 <= Cin_1_c21;
               X_1_c22 <= X_1_c21;
               X_2_c22 <= X_2_c21;
               X_3_c22 <= X_3_c21;
               X_4_c22 <= X_4_c21;
               X_5_c22 <= X_5_c21;
               X_6_c22 <= X_6_c21;
               X_7_c22 <= X_7_c21;
               X_8_c22 <= X_8_c21;
               X_9_c22 <= X_9_c21;
            end if;
            if ce_23 = '1' then
               Cin_1_c23 <= Cin_1_c22;
               X_1_c23 <= X_1_c22;
               X_2_c23 <= X_2_c22;
               X_3_c23 <= X_3_c22;
               X_4_c23 <= X_4_c22;
               X_5_c23 <= X_5_c22;
               X_6_c23 <= X_6_c22;
               X_7_c23 <= X_7_c22;
               X_8_c23 <= X_8_c22;
               X_9_c23 <= X_9_c22;
            end if;
            if ce_24 = '1' then
               Cin_1_c24 <= Cin_1_c23;
               X_1_c24 <= X_1_c23;
               Y_1_c24 <= Y_1_c23;
               X_2_c24 <= X_2_c23;
               Y_2_c24 <= Y_2_c23;
               X_3_c24 <= X_3_c23;
               Y_3_c24 <= Y_3_c23;
               X_4_c24 <= X_4_c23;
               Y_4_c24 <= Y_4_c23;
               X_5_c24 <= X_5_c23;
               Y_5_c24 <= Y_5_c23;
               X_6_c24 <= X_6_c23;
               Y_6_c24 <= Y_6_c23;
               X_7_c24 <= X_7_c23;
               Y_7_c24 <= Y_7_c23;
               X_8_c24 <= X_8_c23;
               Y_8_c24 <= Y_8_c23;
               X_9_c24 <= X_9_c23;
               Y_9_c24 <= Y_9_c23;
            end if;
            if ce_25 = '1' then
               R_1_c25 <= R_1_c24;
               Cin_2_c25 <= Cin_2_c24;
               X_2_c25 <= X_2_c24;
               Y_2_c25 <= Y_2_c24;
               X_3_c25 <= X_3_c24;
               Y_3_c25 <= Y_3_c24;
               X_4_c25 <= X_4_c24;
               Y_4_c25 <= Y_4_c24;
               X_5_c25 <= X_5_c24;
               Y_5_c25 <= Y_5_c24;
               X_6_c25 <= X_6_c24;
               Y_6_c25 <= Y_6_c24;
               X_7_c25 <= X_7_c24;
               Y_7_c25 <= Y_7_c24;
               X_8_c25 <= X_8_c24;
               Y_8_c25 <= Y_8_c24;
               X_9_c25 <= X_9_c24;
               Y_9_c25 <= Y_9_c24;
            end if;
            if ce_26 = '1' then
               R_1_c26 <= R_1_c25;
               R_2_c26 <= R_2_c25;
               Cin_3_c26 <= Cin_3_c25;
               X_3_c26 <= X_3_c25;
               Y_3_c26 <= Y_3_c25;
               X_4_c26 <= X_4_c25;
               Y_4_c26 <= Y_4_c25;
               X_5_c26 <= X_5_c25;
               Y_5_c26 <= Y_5_c25;
               X_6_c26 <= X_6_c25;
               Y_6_c26 <= Y_6_c25;
               X_7_c26 <= X_7_c25;
               Y_7_c26 <= Y_7_c25;
               X_8_c26 <= X_8_c25;
               Y_8_c26 <= Y_8_c25;
               X_9_c26 <= X_9_c25;
               Y_9_c26 <= Y_9_c25;
            end if;
            if ce_27 = '1' then
               R_1_c27 <= R_1_c26;
               R_2_c27 <= R_2_c26;
               R_3_c27 <= R_3_c26;
               Cin_4_c27 <= Cin_4_c26;
               X_4_c27 <= X_4_c26;
               Y_4_c27 <= Y_4_c26;
               X_5_c27 <= X_5_c26;
               Y_5_c27 <= Y_5_c26;
               X_6_c27 <= X_6_c26;
               Y_6_c27 <= Y_6_c26;
               X_7_c27 <= X_7_c26;
               Y_7_c27 <= Y_7_c26;
               X_8_c27 <= X_8_c26;
               Y_8_c27 <= Y_8_c26;
               X_9_c27 <= X_9_c26;
               Y_9_c27 <= Y_9_c26;
            end if;
            if ce_28 = '1' then
               R_1_c28 <= R_1_c27;
               R_2_c28 <= R_2_c27;
               R_3_c28 <= R_3_c27;
               R_4_c28 <= R_4_c27;
               Cin_5_c28 <= Cin_5_c27;
               X_5_c28 <= X_5_c27;
               Y_5_c28 <= Y_5_c27;
               X_6_c28 <= X_6_c27;
               Y_6_c28 <= Y_6_c27;
               X_7_c28 <= X_7_c27;
               Y_7_c28 <= Y_7_c27;
               X_8_c28 <= X_8_c27;
               Y_8_c28 <= Y_8_c27;
               X_9_c28 <= X_9_c27;
               Y_9_c28 <= Y_9_c27;
            end if;
            if ce_29 = '1' then
               R_1_c29 <= R_1_c28;
               R_2_c29 <= R_2_c28;
               R_3_c29 <= R_3_c28;
               R_4_c29 <= R_4_c28;
               R_5_c29 <= R_5_c28;
               Cin_6_c29 <= Cin_6_c28;
               X_6_c29 <= X_6_c28;
               Y_6_c29 <= Y_6_c28;
               X_7_c29 <= X_7_c28;
               Y_7_c29 <= Y_7_c28;
               X_8_c29 <= X_8_c28;
               Y_8_c29 <= Y_8_c28;
               X_9_c29 <= X_9_c28;
               Y_9_c29 <= Y_9_c28;
            end if;
            if ce_30 = '1' then
               R_1_c30 <= R_1_c29;
               R_2_c30 <= R_2_c29;
               R_3_c30 <= R_3_c29;
               R_4_c30 <= R_4_c29;
               R_5_c30 <= R_5_c29;
               R_6_c30 <= R_6_c29;
               Cin_7_c30 <= Cin_7_c29;
               X_7_c30 <= X_7_c29;
               Y_7_c30 <= Y_7_c29;
               X_8_c30 <= X_8_c29;
               Y_8_c30 <= Y_8_c29;
               X_9_c30 <= X_9_c29;
               Y_9_c30 <= Y_9_c29;
            end if;
            if ce_31 = '1' then
               R_1_c31 <= R_1_c30;
               R_2_c31 <= R_2_c30;
               R_3_c31 <= R_3_c30;
               R_4_c31 <= R_4_c30;
               R_5_c31 <= R_5_c30;
               R_6_c31 <= R_6_c30;
               R_7_c31 <= R_7_c30;
               Cin_8_c31 <= Cin_8_c30;
               X_8_c31 <= X_8_c30;
               Y_8_c31 <= Y_8_c30;
               X_9_c31 <= X_9_c30;
               Y_9_c31 <= Y_9_c30;
            end if;
            if ce_32 = '1' then
               R_1_c32 <= R_1_c31;
               R_2_c32 <= R_2_c31;
               R_3_c32 <= R_3_c31;
               R_4_c32 <= R_4_c31;
               R_5_c32 <= R_5_c31;
               R_6_c32 <= R_6_c31;
               R_7_c32 <= R_7_c31;
               R_8_c32 <= R_8_c31;
               Cin_9_c32 <= Cin_9_c31;
               X_9_c32 <= X_9_c31;
               Y_9_c32 <= Y_9_c31;
            end if;
         end if;
      end process;
   Cin_1_c0 <= Cin;
   X_1_c5 <= '0' & X(2 downto 0);
   Y_1_c23 <= '0' & Y(2 downto 0);
   S_1_c24 <= X_1_c24 + Y_1_c24 + Cin_1_c24;
   R_1_c24 <= S_1_c24(2 downto 0);
   Cin_2_c24 <= S_1_c24(3);
   X_2_c5 <= '0' & X(5 downto 3);
   Y_2_c23 <= '0' & Y(5 downto 3);
   S_2_c25 <= X_2_c25 + Y_2_c25 + Cin_2_c25;
   R_2_c25 <= S_2_c25(2 downto 0);
   Cin_3_c25 <= S_2_c25(3);
   X_3_c5 <= '0' & X(8 downto 6);
   Y_3_c23 <= '0' & Y(8 downto 6);
   S_3_c26 <= X_3_c26 + Y_3_c26 + Cin_3_c26;
   R_3_c26 <= S_3_c26(2 downto 0);
   Cin_4_c26 <= S_3_c26(3);
   X_4_c5 <= '0' & X(11 downto 9);
   Y_4_c23 <= '0' & Y(11 downto 9);
   S_4_c27 <= X_4_c27 + Y_4_c27 + Cin_4_c27;
   R_4_c27 <= S_4_c27(2 downto 0);
   Cin_5_c27 <= S_4_c27(3);
   X_5_c5 <= '0' & X(14 downto 12);
   Y_5_c23 <= '0' & Y(14 downto 12);
   S_5_c28 <= X_5_c28 + Y_5_c28 + Cin_5_c28;
   R_5_c28 <= S_5_c28(2 downto 0);
   Cin_6_c28 <= S_5_c28(3);
   X_6_c5 <= '0' & X(17 downto 15);
   Y_6_c23 <= '0' & Y(17 downto 15);
   S_6_c29 <= X_6_c29 + Y_6_c29 + Cin_6_c29;
   R_6_c29 <= S_6_c29(2 downto 0);
   Cin_7_c29 <= S_6_c29(3);
   X_7_c5 <= '0' & X(20 downto 18);
   Y_7_c23 <= '0' & Y(20 downto 18);
   S_7_c30 <= X_7_c30 + Y_7_c30 + Cin_7_c30;
   R_7_c30 <= S_7_c30(2 downto 0);
   Cin_8_c30 <= S_7_c30(3);
   X_8_c5 <= '0' & X(23 downto 21);
   Y_8_c23 <= '0' & Y(23 downto 21);
   S_8_c31 <= X_8_c31 + Y_8_c31 + Cin_8_c31;
   R_8_c31 <= S_8_c31(2 downto 0);
   Cin_9_c31 <= S_8_c31(3);
   X_9_c5 <= '0' & X(26 downto 24);
   Y_9_c23 <= '0' & Y(26 downto 24);
   S_9_c32 <= X_9_c32 + Y_9_c32 + Cin_9_c32;
   R_9_c32 <= S_9_c32(2 downto 0);
   R <= R_9_c32 & R_8_c32 & R_7_c32 & R_6_c32 & R_5_c32 & R_4_c32 & R_3_c32 & R_2_c32 & R_1_c32 ;
end architecture;

--------------------------------------------------------------------------------
--              compressedTable_Freq800_uid37_diff_Freq800_uid42
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity compressedTable_Freq800_uid37_diff_Freq800_uid42 is
    port (clk, ce_33, ce_34 : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(20 downto 0)   );
end entity;

architecture arch of compressedTable_Freq800_uid37_diff_Freq800_uid42 is
signal Y0_c34 :  std_logic_vector(20 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "block";
signal Y1_c34 :  std_logic_vector(20 downto 0);
signal X_c33, X_c34 :  std_logic_vector(9 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_33 = '1' then
               X_c33 <= X;
            end if;
            if ce_34 = '1' then
               X_c34 <= X_c33;
            end if;
         end if;
      end process;
   with X_c34  select  Y0_c34 <= 
      "000000000000000000000" when "0000000000",
      "000100000000001000000" when "0000000001",
      "001000000000100000000" when "0000000010",
      "001100000001001000001" when "0000000011",
      "010000000010000000001" when "0000000100",
      "010100000011001000011" when "0000000101",
      "011000000100100000101" when "0000000110",
      "011100000110001000111" when "0000000111",
      "000000001000000001011" when "0000001000",
      "000100001010001001111" when "0000001001",
      "001000001100100010101" when "0000001010",
      "001100001111001011100" when "0000001011",
      "010000010010000100100" when "0000001100",
      "010100010101001101110" when "0000001101",
      "011000011000100111001" when "0000001110",
      "011100011100010000111" when "0000001111",
      "000000100000001010110" when "0000010000",
      "000100100100010100111" when "0000010001",
      "001000101000101111010" when "0000010010",
      "001100101101011010000" when "0000010011",
      "010000110010010100111" when "0000010100",
      "010100110111100000010" when "0000010101",
      "011000111100111011111" when "0000010110",
      "011101000010100111111" when "0000010111",
      "000001001000100100010" when "0000011000",
      "000101001110110001000" when "0000011001",
      "001001010101001110001" when "0000011010",
      "001101011011111011101" when "0000011011",
      "010001100010111001100" when "0000011100",
      "010101101010001000000" when "0000011101",
      "011001110001100110111" when "0000011110",
      "011101111001010110001" when "0000011111",
      "000010000001010110000" when "0000100000",
      "000110001001100110011" when "0000100001",
      "001010010010000111010" when "0000100010",
      "001110011010111000101" when "0000100011",
      "010010100011111010101" when "0000100100",
      "010110101101001101001" when "0000100101",
      "011010110110110000010" when "0000100110",
      "011111000000100100000" when "0000100111",
      "000011001010101000010" when "0000101000",
      "000111010100111101010" when "0000101001",
      "001011011111100010111" when "0000101010",
      "001111101010011001010" when "0000101011",
      "010011110101100000010" when "0000101100",
      "011000000000110111111" when "0000101101",
      "011100001100100000011" when "0000101110",
      "100000011000011001100" when "0000101111",
      "000100100100100011011" when "0000110000",
      "001000110000111110001" when "0000110001",
      "001100111101101001100" when "0000110010",
      "010001001010100101110" when "0000110011",
      "010101010111110010111" when "0000110100",
      "011001100101010000110" when "0000110101",
      "011101110010111111100" when "0000110110",
      "100010000000111111001" when "0000110111",
      "000110001111001111101" when "0000111000",
      "001010011101110001000" when "0000111001",
      "001110101100100011011" when "0000111010",
      "010010111011100110101" when "0000111011",
      "010111001010111010111" when "0000111100",
      "011011011010100000000" when "0000111101",
      "011111101010010110001" when "0000111110",
      "100011111010011101010" when "0000111111",
      "001000001010110101100" when "0001000000",
      "001100011011011110101" when "0001000001",
      "010000101100011000111" when "0001000010",
      "010100111101100100010" when "0001000011",
      "011001001111000000101" when "0001000100",
      "011101100000101110001" when "0001000101",
      "100001110010101100110" when "0001000110",
      "100110000100111100100" when "0001000111",
      "001010010111011101011" when "0001001000",
      "001110101010001111011" when "0001001001",
      "010010111101010010101" when "0001001010",
      "010111010000100111000" when "0001001011",
      "011011100100001100110" when "0001001100",
      "011111111000000011101" when "0001001101",
      "100100001100001011110" when "0001001110",
      "101000100000100101001" when "0001001111",
      "001100110101001111110" when "0001010000",
      "010001001010001011110" when "0001010001",
      "010101011111011001001" when "0001010010",
      "011001110100110111110" when "0001010011",
      "011110001010100111101" when "0001010100",
      "100010100000101001000" when "0001010101",
      "100110110110111011110" when "0001010110",
      "101011001101011111111" when "0001010111",
      "001111100100010101100" when "0001011000",
      "010011111011011100100" when "0001011001",
      "011000010010110100111" when "0001011010",
      "011100101010011110110" when "0001011011",
      "100001000010011010010" when "0001011100",
      "100101011010100111001" when "0001011101",
      "101001110011000101100" when "0001011110",
      "101110001011110101100" when "0001011111",
      "000010100100110111000" when "0001100000",
      "000110111110001010001" when "0001100001",
      "001011010111101110110" when "0001100010",
      "001111110001100101001" when "0001100011",
      "010100001011101101000" when "0001100100",
      "011000100110000110100" when "0001100101",
      "011101000000110001110" when "0001100110",
      "100001011011101110101" when "0001100111",
      "000101110110111101010" when "0001101000",
      "001010010010011101100" when "0001101001",
      "001110101110001111100" when "0001101010",
      "010011001010010011011" when "0001101011",
      "010111100110101000111" when "0001101100",
      "011100000011010000001" when "0001101101",
      "100000100000001001010" when "0001101110",
      "100100111101010100001" when "0001101111",
      "001001011010110000111" when "0001110000",
      "001101111000011111100" when "0001110001",
      "010010010110100000000" when "0001110010",
      "010110110100110010011" when "0001110011",
      "011011010011010110101" when "0001110100",
      "011111110010001100110" when "0001110101",
      "100100010001010100111" when "0001110110",
      "101000110000101111000" when "0001110111",
      "001101010000011011000" when "0001111000",
      "010001110000011001000" when "0001111001",
      "010110010000101001000" when "0001111010",
      "011010110001001011001" when "0001111011",
      "011111010001111111010" when "0001111100",
      "100011110011000101011" when "0001111101",
      "101000010100011101101" when "0001111110",
      "101100110110000111111" when "0001111111",
      "000001011000000100011" when "0010000000",
      "000101111010010010111" when "0010000001",
      "001010011100110011101" when "0010000010",
      "001110111111100110100" when "0010000011",
      "010011100010101011101" when "0010000100",
      "011000000110000010111" when "0010000101",
      "011100101001101100011" when "0010000110",
      "100001001101101000001" when "0010000111",
      "000101110001110110001" when "0010001000",
      "001010010110010110011" when "0010001001",
      "001110111011001000111" when "0010001010",
      "010011100000001101110" when "0010001011",
      "011000000101100100111" when "0010001100",
      "011100101011001110011" when "0010001101",
      "100001010001001010011" when "0010001110",
      "100101110111011000101" when "0010001111",
      "001010011101111001010" when "0010010000",
      "001111000100101100011" when "0010010001",
      "010011101011110001111" when "0010010010",
      "011000010011001001110" when "0010010011",
      "011100111010110100010" when "0010010100",
      "100001100010110001001" when "0010010101",
      "100110001011000000101" when "0010010110",
      "101010110011100010100" when "0010010111",
      "001111011100010111000" when "0010011000",
      "010100000101011110001" when "0010011001",
      "011000101110110111110" when "0010011010",
      "011101011000100100000" when "0010011011",
      "100010000010100010110" when "0010011100",
      "100110101100110100010" when "0010011101",
      "101011010111011000011" when "0010011110",
      "110000000010001111010" when "0010011111",
      "000100101101011000110" when "0010100000",
      "001001011000110100111" when "0010100001",
      "001110000100100011110" when "0010100010",
      "010010110000100101100" when "0010100011",
      "010111011100111001111" when "0010100100",
      "011100001001100001001" when "0010100101",
      "100000110110011011001" when "0010100110",
      "100101100011100111111" when "0010100111",
      "001010010001000111100" when "0010101000",
      "001110111110111010000" when "0010101001",
      "010011101100111111011" when "0010101010",
      "011000011011010111101" when "0010101011",
      "011101001010000010111" when "0010101100",
      "100001111001000000111" when "0010101101",
      "100110101000010010000" when "0010101110",
      "101011010111110110000" when "0010101111",
      "000000000111101101000" when "0010110000",
      "000100110111110111000" when "0010110001",
      "001001101000010100000" when "0010110010",
      "001110011001000100000" when "0010110011",
      "010011001010000111001" when "0010110100",
      "010111111011011101010" when "0010110101",
      "011100101101000110100" when "0010110110",
      "100001011111000010111" when "0010110111",
      "000110010001010010011" when "0010111000",
      "001011000011110101001" when "0010111001",
      "001111110110101010111" when "0010111010",
      "010100101001110011111" when "0010111011",
      "011001011101010000001" when "0010111100",
      "011110010000111111101" when "0010111101",
      "100011000101000010010" when "0010111110",
      "100111111001011000010" when "0010111111",
      "001100101110000001100" when "0011000000",
      "010001100010111110000" when "0011000001",
      "010110011000001101111" when "0011000010",
      "011011001101110001000" when "0011000011",
      "100000000011100111100" when "0011000100",
      "100100111001110001100" when "0011000101",
      "101001110000001110110" when "0011000110",
      "101110100110111111100" when "0011000111",
      "000011011110000011101" when "0011001000",
      "001000010101011011010" when "0011001001",
      "001101001101000110011" when "0011001010",
      "010010000101000100111" when "0011001011",
      "010110111101010111000" when "0011001100",
      "011011110101111100101" when "0011001101",
      "100000101110110101110" when "0011001110",
      "100101101000000010100" when "0011001111",
      "001010100001100010110" when "0011010000",
      "001111011011010110101" when "0011010001",
      "010100010101011110001" when "0011010010",
      "011001001111111001011" when "0011010011",
      "011110001010101000001" when "0011010100",
      "100011000101101010101" when "0011010101",
      "101000000001000000111" when "0011010110",
      "101100111100101010110" when "0011010111",
      "000001111000101000100" when "0011011000",
      "000110110100111001111" when "0011011001",
      "001011110001011111001" when "0011011010",
      "010000101110011000001" when "0011011011",
      "010101101011100100111" when "0011011100",
      "011010101001000101100" when "0011011101",
      "011111100110111010000" when "0011011110",
      "100100100101000010011" when "0011011111",
      "001001100011011110101" when "0011100000",
      "001110100010001110111" when "0011100001",
      "010011100001010011000" when "0011100010",
      "011000100000101011000" when "0011100011",
      "011101100000010111000" when "0011100100",
      "100010100000010111000" when "0011100101",
      "100111100000101011001" when "0011100110",
      "101100100001010011001" when "0011100111",
      "000001100010001111010" when "0011101000",
      "000110100011011111100" when "0011101001",
      "001011100101000011110" when "0011101010",
      "010000100110111100001" when "0011101011",
      "010101101001001000101" when "0011101100",
      "011010101011101001010" when "0011101101",
      "011111101110011110000" when "0011101110",
      "100100110001100111000" when "0011101111",
      "001001110101000100010" when "0011110000",
      "001110111000110101101" when "0011110001",
      "010011111100111011011" when "0011110010",
      "011001000001010101010" when "0011110011",
      "011110000110000011100" when "0011110100",
      "100011001011000110001" when "0011110101",
      "101000010000011100111" when "0011110110",
      "101101010110001000001" when "0011110111",
      "000010011100000111110" when "0011111000",
      "000111100010011011101" when "0011111001",
      "001100101001000100000" when "0011111010",
      "010001110000000000110" when "0011111011",
      "010110110111010010000" when "0011111100",
      "011011111110110111110" when "0011111101",
      "100001000110110001111" when "0011111110",
      "100110001111000000100" when "0011111111",
      "001011010111100011110" when "0100000000",
      "010000100000011011100" when "0100000001",
      "010101101001100111111" when "0100000010",
      "011010110011001000110" when "0100000011",
      "011111111100111110010" when "0100000100",
      "100101000111001000011" when "0100000101",
      "101010010001100111001" when "0100000110",
      "101111011100011010100" when "0100000111",
      "000100100111100010101" when "0100001000",
      "001001110010111111100" when "0100001001",
      "001110111110110001000" when "0100001010",
      "010100001010110111011" when "0100001011",
      "011001010111010010011" when "0100001100",
      "011110100100000010010" when "0100001101",
      "100011110001000111000" when "0100001110",
      "101000111110100000011" when "0100001111",
      "001110001100001110110" when "0100010000",
      "010011011010010010000" when "0100010001",
      "011000101000101010000" when "0100010010",
      "011101110111010111000" when "0100010011",
      "100011000110011001000" when "0100010100",
      "101000010101101111111" when "0100010101",
      "101101100101011011110" when "0100010110",
      "110010110101011100100" when "0100010111",
      "001000000101110010011" when "0100011000",
      "001101010110011101010" when "0100011001",
      "010010100111011101010" when "0100011010",
      "010111111000110010010" when "0100011011",
      "011101001010011100010" when "0100011100",
      "100010011100011011100" when "0100011101",
      "100111101110101111111" when "0100011110",
      "101101000001011001011" when "0100011111",
      "000010010100011000000" when "0100100000",
      "000111100111101011111" when "0100100001",
      "001100111011010101000" when "0100100010",
      "010010001111010011011" when "0100100011",
      "010111100011100111000" when "0100100100",
      "011100111000001111110" when "0100100101",
      "100010001101001110000" when "0100100110",
      "100111100010100001100" when "0100100111",
      "001100111000001010010" when "0100101000",
      "010010001110001000100" when "0100101001",
      "010111100100011100001" when "0100101010",
      "011100111011000101000" when "0100101011",
      "100010010010000011100" when "0100101100",
      "100111101001010111011" when "0100101101",
      "101101000001000000101" when "0100101110",
      "110010011000111111100" when "0100101111",
      "000111110001010011110" when "0100110000",
      "001101001001111101101" when "0100110001",
      "010010100010111101000" when "0100110010",
      "010111111100010010000" when "0100110011",
      "011101010101111100101" when "0100110100",
      "100010101111111100110" when "0100110101",
      "101000001010010010101" when "0100110110",
      "101101100100111110000" when "0100110111",
      "000010111111111111010" when "0100111000",
      "001000011011010110000" when "0100111001",
      "001101110111000010101" when "0100111010",
      "010011010011000100111" when "0100111011",
      "011000101111011101000" when "0100111100",
      "011110001100001010111" when "0100111101",
      "100011101001001110100" when "0100111110",
      "101001000110101000000" when "0100111111",
      "001110100100010111011" when "0101000000",
      "010100000010011100101" when "0101000001",
      "011001100000110111110" when "0101000010",
      "011110111111101000110" when "0101000011",
      "100100011110101111101" when "0101000100",
      "101001111110001100100" when "0101000101",
      "101111011101111111011" when "0101000110",
      "110100111110001000010" when "0101000111",
      "001010011110100111010" when "0101001000",
      "001111111111011100001" when "0101001001",
      "010101100000100111001" when "0101001010",
      "011011000010001000010" when "0101001011",
      "100000100011111111011" when "0101001100",
      "100110000110001100110" when "0101001101",
      "101011101000110000010" when "0101001110",
      "110001001011101001111" when "0101001111",
      "000110101110111001101" when "0101010000",
      "001100010010011111110" when "0101010001",
      "010001110110011100000" when "0101010010",
      "010111011010101110100" when "0101010011",
      "011100111111010111011" when "0101010100",
      "100010100100010110100" when "0101010101",
      "101000001001101011111" when "0101010110",
      "101101101111010111101" when "0101010111",
      "000011010101011001110" when "0101011000",
      "001000111011110010011" when "0101011001",
      "001110100010100001010" when "0101011010",
      "010100001001100110101" when "0101011011",
      "011001110001000010100" when "0101011100",
      "011111011000110100110" when "0101011101",
      "100101000000111101101" when "0101011110",
      "101010101001011100111" when "0101011111",
      "000000010010010010110" when "0101100000",
      "000101111011011111010" when "0101100001",
      "001011100101000010010" when "0101100010",
      "010001001110111011111" when "0101100011",
      "010110111001001100001" when "0101100100",
      "011100100011110011000" when "0101100101",
      "100010001110110000101" when "0101100110",
      "100111111010000100111" when "0101100111",
      "001101100101101111111" when "0101101000",
      "010011010001110001101" when "0101101001",
      "011000111110001010001" when "0101101010",
      "011110101010111001011" when "0101101011",
      "100100010111111111100" when "0101101100",
      "101010000101011100011" when "0101101101",
      "101111110011010000001" when "0101101110",
      "110101100001011010110" when "0101101111",
      "001011001111111100011" when "0101110000",
      "010000111110110100110" when "0101110001",
      "010110101110000100010" when "0101110010",
      "011100011101101010100" when "0101110011",
      "100010001101100111111" when "0101110100",
      "100111111101111100010" when "0101110101",
      "101101101110100111101" when "0101110110",
      "110011011111101010001" when "0101110111",
      "001001010001000011101" when "0101111000",
      "001111000010110100010" when "0101111001",
      "010100110100111100000" when "0101111010",
      "011010100111011010111" when "0101111011",
      "100000011010010000111" when "0101111100",
      "100110001101011110001" when "0101111101",
      "101100000001000010101" when "0101111110",
      "110001110100111110010" when "0101111111",
      "000111101001010001010" when "0110000000",
      "001101011101111011100" when "0110000001",
      "010011010010111101000" when "0110000010",
      "011001001000010101111" when "0110000011",
      "011110111110000110000" when "0110000100",
      "100100110100001101101" when "0110000101",
      "101010101010101100101" when "0110000110",
      "110000100001100011000" when "0110000111",
      "000110011000110000110" when "0110001000",
      "001100010000010110000" when "0110001001",
      "010010001000010010111" when "0110001010",
      "011000000000100111001" when "0110001011",
      "011101111001010010111" when "0110001100",
      "100011110010010110010" when "0110001101",
      "101001101011110001010" when "0110001110",
      "101111100101100011110" when "0110001111",
      "000101011111101101111" when "0110010000",
      "001011011010001111110" when "0110010001",
      "010001010101001001010" when "0110010010",
      "010111010000011010011" when "0110010011",
      "011101001100000011010" when "0110010100",
      "100011001000000011111" when "0110010101",
      "101001000100011100010" when "0110010110",
      "101111000001001100100" when "0110010111",
      "000100111110010100011" when "0110011000",
      "001010111011110100010" when "0110011001",
      "010000111001101011111" when "0110011010",
      "010110110111111011100" when "0110011011",
      "011100110110100010111" when "0110011100",
      "100010110101100010010" when "0110011101",
      "101000110100111001101" when "0110011110",
      "101110110100101000111" when "0110011111",
      "000100110100110000010" when "0110100000",
      "001010110101001111100" when "0110100001",
      "010000110110000110111" when "0110100010",
      "010110110111010110010" when "0110100011",
      "011100111000111101110" when "0110100100",
      "100010111010111101011" when "0110100101",
      "101000111101010101001" when "0110100110",
      "101111000000000101001" when "0110100111",
      "000101000011001101010" when "0110101000",
      "001011000110101101100" when "0110101001",
      "010001001010100110000" when "0110101010",
      "010111001110110110111" when "0110101011",
      "011101010011011111111" when "0110101100",
      "100011011000100001010" when "0110101101",
      "101001011101111011000" when "0110101110",
      "101111100011101101000" when "0110101111",
      "000101101001110111100" when "0110110000",
      "001011110000011010010" when "0110110001",
      "010001110111010101100" when "0110110010",
      "010111111110101001010" when "0110110011",
      "011110000110010101011" when "0110110100",
      "100100001110011010000" when "0110110101",
      "101010010110110111001" when "0110110110",
      "110000011111101100111" when "0110110111",
      "000110101000111011001" when "0110111000",
      "001100110010100010000" when "0110111001",
      "010010111100100001100" when "0110111010",
      "011001000110111001100" when "0110111011",
      "011111010001101010011" when "0110111100",
      "100101011100110011110" when "0110111101",
      "101011101000010101111" when "0110111110",
      "110001110100010000111" when "0110111111",
      "001000000000100100100" when "0111000000",
      "001110001101010000111" when "0111000001",
      "010100011010010110001" when "0111000010",
      "011010100111110100010" when "0111000011",
      "100000110101101011001" when "0111000100",
      "100111000011111010111" when "0111000101",
      "101101010010100011101" when "0111000110",
      "110011100001100101010" when "0111000111",
      "001001110000111111111" when "0111001000",
      "010000000000110011011" when "0111001001",
      "010110010000111111111" when "0111001010",
      "011100100001100101100" when "0111001011",
      "100010110010100100001" when "0111001100",
      "101001000011111011111" when "0111001101",
      "101111010101101100101" when "0111001110",
      "110101100111110110100" when "0111001111",
      "001011111010011001101" when "0111010000",
      "010010001101010101111" when "0111010001",
      "011000100000101011010" when "0111010010",
      "011110110100011010000" when "0111010011",
      "100101001000100001111" when "0111010100",
      "101011011101000011000" when "0111010101",
      "110001110001111101100" when "0111010110",
      "111000000111010001010" when "0111010111",
      "001110011100111110011" when "0111011000",
      "010100110011000100111" when "0111011001",
      "011011001001100100110" when "0111011010",
      "100001100000011110001" when "0111011011",
      "100111110111110000111" when "0111011100",
      "101110001111011101001" when "0111011101",
      "110100100111100010111" when "0111011110",
      "111011000000000010000" when "0111011111",
      "000001011000111010111" when "0111100000",
      "000111110010001101001" when "0111100001",
      "001110001011111001001" when "0111100010",
      "010100100101111110101" when "0111100011",
      "011011000000011101111" when "0111100100",
      "100001011011010110110" when "0111100101",
      "100111110110101001010" when "0111100110",
      "101110010010010101101" when "0111100111",
      "000100101110011011101" when "0111101000",
      "001011001010111011011" when "0111101001",
      "010001100111110101000" when "0111101010",
      "011000000101001000011" when "0111101011",
      "011110100010110101101" when "0111101100",
      "100101000000111100110" when "0111101101",
      "101011011111011101110" when "0111101110",
      "110001111110011000101" when "0111101111",
      "001000011101101101100" when "0111110000",
      "001110111101011100011" when "0111110001",
      "010101011101100101010" when "0111110010",
      "011011111110001000001" when "0111110011",
      "100010011111000101000" when "0111110100",
      "101001000000011100000" when "0111110101",
      "101111100010001101001" when "0111110110",
      "110110000100011000010" when "0111110111",
      "001100100110111101101" when "0111111000",
      "010011001001111101001" when "0111111001",
      "011001101101010110111" when "0111111010",
      "100000010001001010111" when "0111111011",
      "100110110101011001000" when "0111111100",
      "101101011010000001100" when "0111111101",
      "110011111111000100010" when "0111111110",
      "111010100100100001011" when "0111111111",
      "000100010110010111111" when "1000000000",
      "000110110001101110001" when "1000000001",
      "001001001101001110001" when "1000000010",
      "001011101000110111110" when "1000000011",
      "001110000100101011010" when "1000000100",
      "010000100000101000011" when "1000000101",
      "010010111100101111010" when "1000000110",
      "010101011001000000000" when "1000000111",
      "000111110101011010011" when "1000001000",
      "001010010001111110101" when "1000001001",
      "001100101110101100101" when "1000001010",
      "001111001011100100100" when "1000001011",
      "010001101000100110001" when "1000001100",
      "010100000101110001101" when "1000001101",
      "010110100011000110111" when "1000001110",
      "011001000000100110000" when "1000001111",
      "001011011110001110111" when "1000010000",
      "001101111100000001110" when "1000010001",
      "010000011001111110100" when "1000010010",
      "010010111000000101000" when "1000010011",
      "010101010110010101100" when "1000010100",
      "010111110100101111110" when "1000010101",
      "011010010011010100000" when "1000010110",
      "011100110010000010010" when "1000010111",
      "001111010000111010010" when "1000011000",
      "010001101111111100011" when "1000011001",
      "010100001111001000010" when "1000011010",
      "010110101110011110010" when "1000011011",
      "011001001101111110001" when "1000011100",
      "011011101101101000000" when "1000011101",
      "011110001101011011111" when "1000011110",
      "100000101101011001101" when "1000011111",
      "000011001101100001100" when "1000100000",
      "000101101101110011011" when "1000100001",
      "001000001110001111010" when "1000100010",
      "001010101110110101001" when "1000100011",
      "001101001111100101001" when "1000100100",
      "001111110000011111001" when "1000100101",
      "010010010001100011001" when "1000100110",
      "010100110010110001010" when "1000100111",
      "000111010100001001100" when "1000101000",
      "001001110101101011110" when "1000101001",
      "001100010111011000010" when "1000101010",
      "001110111001001110110" when "1000101011",
      "010001011011001111011" when "1000101100",
      "010011111101011010001" when "1000101101",
      "010110011111101111000" when "1000101110",
      "011001000010001110001" when "1000101111",
      "001011100100110111011" when "1000110000",
      "001110000111101010110" when "1000110001",
      "010000101010101000010" when "1000110010",
      "010011001101110000000" when "1000110011",
      "010101110001000010000" when "1000110100",
      "011000010100011110001" when "1000110101",
      "011010111000000100101" when "1000110110",
      "011101011011110101010" when "1000110111",
      "001111111111110000000" when "1000111000",
      "010010100011110101001" when "1000111001",
      "010101001000000100100" when "1000111010",
      "010111101100011110001" when "1000111011",
      "011010010001000010001" when "1000111100",
      "011100110101110000011" when "1000111101",
      "011111011010101000111" when "1000111110",
      "100001111111101011101" when "1000111111",
      "000100100100111000110" when "1001000000",
      "000111001010010000010" when "1001000001",
      "001001101111110010001" when "1001000010",
      "001100010101011110010" when "1001000011",
      "001110111011010100110" when "1001000100",
      "010001100001010101101" when "1001000101",
      "010100000111100000111" when "1001000110",
      "010110101101110110101" when "1001000111",
      "001001010100010110101" when "1001001000",
      "001011111011000001001" when "1001001001",
      "001110100001110110000" when "1001001010",
      "010001001000110101011" when "1001001011",
      "010011101111111111001" when "1001001100",
      "010110010111010011011" when "1001001101",
      "011000111110110010001" when "1001001110",
      "011011100110011011010" when "1001001111",
      "001110001110001110111" when "1001010000",
      "010000110110001101000" when "1001010001",
      "010011011110010101101" when "1001010010",
      "010110000110101000110" when "1001010011",
      "011000101111000110100" when "1001010100",
      "011011010111101110110" when "1001010101",
      "011110000000100001100" when "1001010110",
      "100000101001011110110" when "1001010111",
      "000011010010100110101" when "1001011000",
      "000101111011111001001" when "1001011001",
      "001000100101010110001" when "1001011010",
      "001011001110111101110" when "1001011011",
      "001101111000110000000" when "1001011100",
      "010000100010101100111" when "1001011101",
      "010011001100110100011" when "1001011110",
      "010101110111000110100" when "1001011111",
      "001000100001100011010" when "1001100000",
      "001011001100001010101" when "1001100001",
      "001101110110111100110" when "1001100010",
      "010000100001111001100" when "1001100011",
      "010011001101000001000" when "1001100100",
      "010101111000010011001" when "1001100101",
      "011000100011110000000" when "1001100110",
      "011011001111010111101" when "1001100111",
      "001101111011001010000" when "1001101000",
      "010000100111000111000" when "1001101001",
      "010011010011001110111" when "1001101010",
      "010101111111100001100" when "1001101011",
      "011000101011111110110" when "1001101100",
      "011011011000100111000" when "1001101101",
      "011110000101011001111" when "1001101110",
      "100000110010010111101" when "1001101111",
      "000011011111100000010" when "1001110000",
      "000110001100110011101" when "1001110001",
      "001000111010010001110" when "1001110010",
      "001011100111111010111" when "1001110011",
      "001110010101101110110" when "1001110100",
      "010001000011101101101" when "1001110101",
      "010011110001110111010" when "1001110110",
      "010110100000001011111" when "1001110111",
      "001001001110101011010" when "1001111000",
      "001011111101010101101" when "1001111001",
      "001110101100001011000" when "1001111010",
      "010001011011001011001" when "1001111011",
      "010100001010010110011" when "1001111100",
      "010110111001101100100" when "1001111101",
      "011001101001001101101" when "1001111110",
      "011100011000111001101" when "1001111111",
      "001111001000110000101" when "1010000000",
      "010001111000110010110" when "1010000001",
      "010100101000111111110" when "1010000010",
      "010111011001010111111" when "1010000011",
      "011010001001111011000" when "1010000100",
      "011100111010101001001" when "1010000101",
      "011111101011100010010" when "1010000110",
      "100010011100100110100" when "1010000111",
      "000101001101110101111" when "1010001000",
      "000111111111010000010" when "1010001001",
      "001010110000110101110" when "1010001010",
      "001101100010100110011" when "1010001011",
      "010000010100100010001" when "1010001100",
      "010011000110101001000" when "1010001101",
      "010101111000111011000" when "1010001110",
      "011000101011011000001" when "1010001111",
      "001011011110000000011" when "1010010000",
      "001110010000110011111" when "1010010001",
      "010001000011110010100" when "1010010010",
      "010011110110111100011" when "1010010011",
      "010110101010010001011" when "1010010100",
      "011001011101110001101" when "1010010101",
      "011100010001011101001" when "1010010110",
      "011111000101010011110" when "1010010111",
      "000001111001010101110" when "1010011000",
      "000100101101100011000" when "1010011001",
      "000111100001111011100" when "1010011010",
      "001010010110011111010" when "1010011011",
      "001101001011001110010" when "1010011100",
      "010000000000001000101" when "1010011101",
      "010010110101001110010" when "1010011110",
      "010101101010011111010" when "1010011111",
      "001000011111111011101" when "1010100000",
      "001011010101100011010" when "1010100001",
      "001110001011010110010" when "1010100010",
      "010001000001010100101" when "1010100011",
      "010011110111011110100" when "1010100100",
      "010110101101110011101" when "1010100101",
      "011001100100010100001" when "1010100110",
      "011100011011000000001" when "1010100111",
      "001111010001110111101" when "1010101000",
      "010010001000111010011" when "1010101001",
      "010101000000001000101" when "1010101010",
      "010111110111100010011" when "1010101011",
      "011010101111000111101" when "1010101100",
      "011101100110111000011" when "1010101101",
      "100000011110110100100" when "1010101110",
      "100011010110111100001" when "1010101111",
      "000110001111001111011" when "1010110000",
      "001001000111101110001" when "1010110001",
      "001100000000011000011" when "1010110010",
      "001110111001001110001" when "1010110011",
      "010001110010001111100" when "1010110100",
      "010100101011011100011" when "1010110101",
      "010111100100110100111" when "1010110110",
      "011010011110011001000" when "1010110111",
      "001101011000001000110" when "1010111000",
      "010000010010000100000" when "1010111001",
      "010011001100001011000" when "1010111010",
      "010110000110011101101" when "1010111011",
      "011001000000111011110" when "1010111100",
      "011011111011100101110" when "1010111101",
      "011110110110011011010" when "1010111110",
      "100001110001011100100" when "1010111111",
      "000100101100101001011" when "1011000000",
      "000111101000000010001" when "1011000001",
      "001010100011100110100" when "1011000010",
      "001101011111010110100" when "1011000011",
      "010000011011010010011" when "1011000100",
      "010011010111011010000" when "1011000101",
      "010110010011101101010" when "1011000110",
      "011001010000001100011" when "1011000111",
      "001100001100110111011" when "1011001000",
      "001111001001101110000" when "1011001001",
      "010010000110110000100" when "1011001010",
      "010101000011111110111" when "1011001011",
      "011000000001011001000" when "1011001100",
      "011010111110111111000" when "1011001101",
      "011101111100110000111" when "1011001110",
      "100000111010101110101" when "1011001111",
      "000011111000111000010" when "1011010000",
      "000110110111001101110" when "1011010001",
      "001001110101101111001" when "1011010010",
      "001100110100011100100" when "1011010011",
      "001111110011010101110" when "1011010100",
      "010010110010011010111" when "1011010101",
      "010101110001101100000" when "1011010110",
      "011000110001001001001" when "1011010111",
      "001011110000110010001" when "1011011000",
      "001110110000100111010" when "1011011001",
      "010001110000101000010" when "1011011010",
      "010100110000110101010" when "1011011011",
      "010111110001001110011" when "1011011100",
      "011010110001110011100" when "1011011101",
      "011101110010100100101" when "1011011110",
      "100000110011100001110" when "1011011111",
      "000011110100101011000" when "1011100000",
      "000110110110000000011" when "1011100001",
      "001001110111100001110" when "1011100010",
      "001100111001001111011" when "1011100011",
      "001111111011001001000" when "1011100100",
      "010010111101001110110" when "1011100101",
      "010101111111100000101" when "1011100110",
      "011001000001111110101" when "1011100111",
      "001100000100101000111" when "1011101000",
      "001111000111011111010" when "1011101001",
      "010010001010100001110" when "1011101010",
      "010101001101110000101" when "1011101011",
      "011000010001001011100" when "1011101100",
      "011011010100110010110" when "1011101101",
      "011110011000100110001" when "1011101110",
      "100001011100100101110" when "1011101111",
      "000100100000110001110" when "1011110000",
      "000111100101001001111" when "1011110001",
      "001010101001101110011" when "1011110010",
      "001101101110011111001" when "1011110011",
      "010000110011011100001" when "1011110100",
      "010011111000100101100" when "1011110101",
      "010110111101111011010" when "1011110110",
      "011010000011011101010" when "1011110111",
      "001101001001001011110" when "1011111000",
      "010000001111000110100" when "1011111001",
      "010011010101001101101" when "1011111010",
      "010110011011100001001" when "1011111011",
      "011001100010000001000" when "1011111100",
      "011100101000101101011" when "1011111101",
      "011111101111100110001" when "1011111110",
      "100010110110101011011" when "1011111111",
      "000101111101111101000" when "1100000000",
      "001001000101011011001" when "1100000001",
      "001100001101000101101" when "1100000010",
      "001111010100111100110" when "1100000011",
      "010010011101000000010" when "1100000100",
      "010101100101010000011" when "1100000101",
      "011000101101101100111" when "1100000110",
      "011011110110010110000" when "1100000111",
      "001110111111001011110" when "1100001000",
      "010010001000001110000" when "1100001001",
      "010101010001011100110" when "1100001010",
      "011000011010111000001" when "1100001011",
      "011011100100100000001" when "1100001100",
      "011110101110010100110" when "1100001101",
      "100001111000010101111" when "1100001110",
      "100101000010100011110" when "1100001111",
      "001000001100111110010" when "1100010000",
      "001011010111100101011" when "1100010001",
      "001110100010011001001" when "1100010010",
      "010001101101011001101" when "1100010011",
      "010100111000100110111" when "1100010100",
      "011000000100000000110" when "1100010101",
      "011011001111100111011" when "1100010110",
      "011110011011011010110" when "1100010111",
      "000001100111011010110" when "1100011000",
      "000100110011100111101" when "1100011001",
      "001000000000000001010" when "1100011010",
      "001011001100100111101" when "1100011011",
      "001110011001011010111" when "1100011100",
      "010001100110011010111" when "1100011101",
      "010100110011100111101" when "1100011110",
      "011000000001000001010" when "1100011111",
      "001011001110100111110" when "1100100000",
      "001110011100011011001" when "1100100001",
      "010001101010011011011" when "1100100010",
      "010100111000101000011" when "1100100011",
      "011000000111000010011" when "1100100100",
      "011011010101101001011" when "1100100101",
      "011110100100011101001" when "1100100110",
      "100001110011011101111" when "1100100111",
      "000101000010101011101" when "1100101000",
      "001000010010000110010" when "1100101001",
      "001011100001101101111" when "1100101010",
      "001110110001100010011" when "1100101011",
      "010010000001100100000" when "1100101100",
      "010101010001110010101" when "1100101101",
      "011000100010001110010" when "1100101110",
      "011011110010110110111" when "1100101111",
      "001111000011101100101" when "1100110000",
      "010010010100101111011" when "1100110001",
      "010101100101111111010" when "1100110010",
      "011000110111011100001" when "1100110011",
      "011100001001000110001" when "1100110100",
      "011111011010111101010" when "1100110101",
      "100010101101000001100" when "1100110110",
      "100101111111010010111" when "1100110111",
      "001001010001110001100" when "1100111000",
      "001100100100011101001" when "1100111001",
      "001111110111010110000" when "1100111010",
      "010011001010011100000" when "1100111011",
      "010110011101101111010" when "1100111100",
      "011001110001001111110" when "1100111101",
      "011101000100111101100" when "1100111110",
      "100000011000111000011" when "1100111111",
      "000011101101000000101" when "1101000000",
      "000111000001010110000" when "1101000001",
      "001010010101111000110" when "1101000010",
      "001101101010101000110" when "1101000011",
      "010000111111100110001" when "1101000100",
      "010100010100110000110" when "1101000101",
      "010111101010001000110" when "1101000110",
      "011010111111101110000" when "1101000111",
      "001110010101100000101" when "1101001000",
      "010001101011100000110" when "1101001001",
      "010101000001101110001" when "1101001010",
      "011000011000001000111" when "1101001011",
      "011011101110110001001" when "1101001100",
      "011111000101100110110" when "1101001101",
      "100010011100101001111" when "1101001110",
      "100101110011111010011" when "1101001111",
      "001001001011011000011" when "1101010000",
      "001100100011000011110" when "1101010001",
      "001111111010111100110" when "1101010010",
      "010011010011000011001" when "1101010011",
      "010110101011010111001" when "1101010100",
      "011010000011111000101" when "1101010101",
      "011101011100100111101" when "1101010110",
      "100000110101100100001" when "1101010111",
      "000100001110101110010" when "1101011000",
      "000111101000000110000" when "1101011001",
      "001011000001101011010" when "1101011010",
      "001110011011011110010" when "1101011011",
      "010001110101011110110" when "1101011100",
      "010101001111101100111" when "1101011101",
      "011000101010001000110" when "1101011110",
      "011100000100110010001" when "1101011111",
      "001111011111101001010" when "1101100000",
      "010010111010101110001" when "1101100001",
      "010110010110000000101" when "1101100010",
      "011001110001100000111" when "1101100011",
      "011101001101001110111" when "1101100100",
      "100000101001001010100" when "1101100101",
      "100100000101010100000" when "1101100110",
      "100111100001101011010" when "1101100111",
      "001010111110010000010" when "1101101000",
      "001110011011000011000" when "1101101001",
      "010001111000000011101" when "1101101010",
      "010101010101010010000" when "1101101011",
      "011000110010101110010" when "1101101100",
      "011100010000011000011" when "1101101101",
      "011111101110010000011" when "1101101110",
      "100011001100010110001" when "1101101111",
      "000110101010101001111" when "1101110000",
      "001010001001001011100" when "1101110001",
      "001101100111111011000" when "1101110010",
      "010001000110111000100" when "1101110011",
      "010100100110000011111" when "1101110100",
      "011000000101011101010" when "1101110101",
      "011011100101000100101" when "1101110110",
      "011111000100111001111" when "1101110111",
      "000010100100111101001" when "1101111000",
      "000110000101001110100" when "1101111001",
      "001001100101101101111" when "1101111010",
      "001101000110011011010" when "1101111011",
      "010000100111010110101" when "1101111100",
      "010100001000100000001" when "1101111101",
      "010111101001110111110" when "1101111110",
      "011011001011011101011" when "1101111111",
      "001110101101010001001" when "1110000000",
      "010010001111010011000" when "1110000001",
      "010101110001100011001" when "1110000010",
      "011001010100000001010" when "1110000011",
      "011100110110101101101" when "1110000100",
      "100000011001101000001" when "1110000101",
      "100011111100110000110" when "1110000110",
      "100111100000000111101" when "1110000111",
      "001011000011101100110" when "1110001000",
      "001110100111100000001" when "1110001001",
      "010010001011100001110" when "1110001010",
      "010101101111110001101" when "1110001011",
      "011001010100001111110" when "1110001100",
      "011100111000111100001" when "1110001101",
      "100000011101110110111" when "1110001110",
      "100100000010111111111" when "1110001111",
      "000111101000010111010" when "1110010000",
      "001011001101111100111" when "1110010001",
      "001110110011110001000" when "1110010010",
      "010010011001110011011" when "1110010011",
      "010110000000000100010" when "1110010100",
      "011001100110100011011" when "1110010101",
      "011101001101010001000" when "1110010110",
      "100000110100001101001" when "1110010111",
      "000100011011010111100" when "1110011000",
      "001000000010110000100" when "1110011001",
      "001011101010010111111" when "1110011010",
      "001111010010001101110" when "1110011011",
      "010010111010010010010" when "1110011100",
      "010110100010100101001" when "1110011101",
      "011010001011000110100" when "1110011110",
      "011101110011110110100" when "1110011111",
      "000001011100110101000" when "1110100000",
      "000101000110000010001" when "1110100001",
      "001000101111011101110" when "1110100010",
      "001100011001001000000" when "1110100011",
      "010000000011000000111" when "1110100100",
      "010011101101001000011" when "1110100101",
      "010111010111011110100" when "1110100110",
      "011011000010000011011" when "1110100111",
      "001110101100110110111" when "1110101000",
      "010010010111111001000" when "1110101001",
      "010110000011001001110" when "1110101010",
      "011001101110101001011" when "1110101011",
      "011101011010010111101" when "1110101100",
      "100001000110010100101" when "1110101101",
      "100100110010100000011" when "1110101110",
      "101000011110111011000" when "1110101111",
      "001100001011100100010" when "1110110000",
      "001111111000011100011" when "1110110001",
      "010011100101100011011" when "1110110010",
      "010111010010111001001" when "1110110011",
      "011011000000011101110" when "1110110100",
      "011110101110010001010" when "1110110101",
      "100010011100010011100" when "1110110110",
      "100110001010100100110" when "1110110111",
      "001001111001000100111" when "1110111000",
      "001101100111110011111" when "1110111001",
      "010001010110110001111" when "1110111010",
      "010101000101111110110" when "1110111011",
      "011000110101011010101" when "1110111100",
      "011100100101000101011" when "1110111101",
      "100000010100111111010" when "1110111110",
      "100100000101001000000" when "1110111111",
      "000111110101011111111" when "1111000000",
      "001011100110000110110" when "1111000001",
      "001111010110111100101" when "1111000010",
      "010011001000000001101" when "1111000011",
      "010110111001010101101" when "1111000100",
      "011010101010111000110" when "1111000101",
      "011110011100101011000" when "1111000110",
      "100010001110101100011" when "1111000111",
      "000110000000111100111" when "1111001000",
      "001001110011011100100" when "1111001001",
      "001101100110001011010" when "1111001010",
      "010001011001001001010" when "1111001011",
      "010101001100010110011" when "1111001100",
      "011000111111110010111" when "1111001101",
      "011100110011011110011" when "1111001110",
      "100000100111011001010" when "1111001111",
      "000100011011100011011" when "1111010000",
      "001000001111111100110" when "1111010001",
      "001100000100100101011" when "1111010010",
      "001111111001011101010" when "1111010011",
      "010011101110100100100" when "1111010100",
      "010111100011111011001" when "1111010101",
      "011011011001100001000" when "1111010110",
      "011111001111010110010" when "1111010111",
      "000011000101011011000" when "1111011000",
      "000110111011101111000" when "1111011001",
      "001010110010010010011" when "1111011010",
      "001110101001000101010" when "1111011011",
      "010010100000000111100" when "1111011100",
      "010110010111011001010" when "1111011101",
      "011010001110111010100" when "1111011110",
      "011110000110101011001" when "1111011111",
      "000001111110101011011" when "1111100000",
      "000101110110111011000" when "1111100001",
      "001001101111011010010" when "1111100010",
      "001101101000001000111" when "1111100011",
      "010001100001000111010" when "1111100100",
      "010101011010010101001" when "1111100101",
      "011001010011110010100" when "1111100110",
      "011101001101011111100" when "1111100111",
      "000001000111011100010" when "1111101000",
      "000101000001101000100" when "1111101001",
      "001000111100000100011" when "1111101010",
      "001100110110110000000" when "1111101011",
      "010000110001101011010" when "1111101100",
      "010100101100110110010" when "1111101101",
      "011000101000010000111" when "1111101110",
      "011100100011111011010" when "1111101111",
      "000000011111110101011" when "1111110000",
      "000100011011111111010" when "1111110001",
      "001000011000011000111" when "1111110010",
      "001100010101000010010" when "1111110011",
      "010000010001111011100" when "1111110100",
      "010100001111000100100" when "1111110101",
      "011000001100011101011" when "1111110110",
      "011100001010000110001" when "1111110111",
      "000000000111111110101" when "1111111000",
      "000100000110000111001" when "1111111001",
      "001000000100011111100" when "1111111010",
      "001100000011000111101" when "1111111011",
      "010000000001111111111" when "1111111100",
      "010100000001000111111" when "1111111101",
      "011000000000100000000" when "1111111110",
      "011100000000001000000" when "1111111111",
      "---------------------" when others;
   Y1_c34 <= Y0_c34; -- for the possible blockram register
   Y <= Y1_c34;
end architecture;

--------------------------------------------------------------------------------
--                       compressedTable_Freq800_uid37
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Luc Forget, Maxime Christ (2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity compressedTable_Freq800_uid37 is
    port (clk, ce_33, ce_34, ce_35 : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of compressedTable_Freq800_uid37 is
   component compressedTable_Freq800_uid37_subsampling_Freq800_uid39 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(8 downto 0)   );
   end component;

   component compressedTable_Freq800_uid37_diff_Freq800_uid42 is
      port ( clk, ce_33, ce_34 : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(20 downto 0)   );
   end component;

signal X_subsampling_c32 :  std_logic_vector(6 downto 0);
signal Y_subsampling_c32, Y_subsampling_c33, Y_subsampling_c34, Y_subsampling_c35 :  std_logic_vector(8 downto 0);
signal Y_subsampling_copy40_c32 :  std_logic_vector(8 downto 0);
signal Y_diff_c34, Y_diff_c35 :  std_logic_vector(20 downto 0);
signal fullOut_topbits_c35 :  std_logic_vector(8 downto 0);
signal fullOut_c35 :  std_logic_vector(27 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_33 = '1' then
               Y_subsampling_c33 <= Y_subsampling_c32;
            end if;
            if ce_34 = '1' then
               Y_subsampling_c34 <= Y_subsampling_c33;
            end if;
            if ce_35 = '1' then
               Y_subsampling_c35 <= Y_subsampling_c34;
               Y_diff_c35 <= Y_diff_c34;
            end if;
         end if;
      end process;
   X_subsampling_c32 <= X(9 downto 3);
   compressedTable_Freq800_uid37_subsampling: compressedTable_Freq800_uid37_subsampling_Freq800_uid39
      port map ( X => X_subsampling_c32,
                 Y => Y_subsampling_copy40_c32);
   Y_subsampling_c32 <= Y_subsampling_copy40_c32; -- output copy to hold a pipeline register if needed
   compressedTable_Freq800_uid37_diff: compressedTable_Freq800_uid37_diff_Freq800_uid42
      port map ( clk  => clk,
                 ce_33 => ce_33,
                 ce_34=> ce_34,
                 X => X,
                 Y => Y_diff_c34);
   fullOut_topbits_c35 <= Y_subsampling_c35 + ("0000000"& (Y_diff_c35(20 downto 19)));
   fullOut_c35 <= fullOut_topbits_c35 & (Y_diff_c35(18 downto 0));
   Y <= fullOut_c35;
end architecture;

--------------------------------------------------------------------------------
--                      FixFunctionByTable_Freq800_uid35
-- Evaluator for exp(x*1b-1) on [-1,1) for lsbIn=-9 (wIn=10), msbout=0, lsbOut=-27 (wOut=28). Out interval: [0.606531; 1.64711]. Output is unsigned

-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq800_uid35 is
    port (clk, ce_33, ce_34, ce_35 : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq800_uid35 is
   component compressedTable_Freq800_uid37 is
      port ( clk, ce_33, ce_34, ce_35 : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(27 downto 0)   );
   end component;

begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_33 = '1' then
            end if;
            if ce_34 = '1' then
            end if;
            if ce_35 = '1' then
            end if;
         end if;
      end process;
   compressedTable: compressedTable_Freq800_uid37
      port map ( clk  => clk,
                 ce_33 => ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 X => X,
                 Y => Y);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_18_Freq800_uid48
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 38 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_18_Freq800_uid48 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38 : in std_logic;
          X : in  std_logic_vector(17 downto 0);
          Y : in  std_logic_vector(17 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of IntAdder_18_Freq800_uid48 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3, Cin_0_c4, Cin_0_c5, Cin_0_c6, Cin_0_c7, Cin_0_c8, Cin_0_c9, Cin_0_c10, Cin_0_c11, Cin_0_c12, Cin_0_c13, Cin_0_c14, Cin_0_c15, Cin_0_c16, Cin_0_c17, Cin_0_c18, Cin_0_c19, Cin_0_c20, Cin_0_c21, Cin_0_c22, Cin_0_c23, Cin_0_c24, Cin_0_c25, Cin_0_c26, Cin_0_c27, Cin_0_c28, Cin_0_c29, Cin_0_c30, Cin_0_c31, Cin_0_c32, Cin_0_c33 :  std_logic;
signal X_0_c32, X_0_c33 :  std_logic_vector(3 downto 0);
signal Y_0_c32, Y_0_c33 :  std_logic_vector(3 downto 0);
signal S_0_c33 :  std_logic_vector(3 downto 0);
signal R_0_c33, R_0_c34, R_0_c35, R_0_c36, R_0_c37, R_0_c38 :  std_logic_vector(2 downto 0);
signal Cin_1_c33, Cin_1_c34 :  std_logic;
signal X_1_c32, X_1_c33, X_1_c34 :  std_logic_vector(3 downto 0);
signal Y_1_c32, Y_1_c33, Y_1_c34 :  std_logic_vector(3 downto 0);
signal S_1_c34 :  std_logic_vector(3 downto 0);
signal R_1_c34, R_1_c35, R_1_c36, R_1_c37, R_1_c38 :  std_logic_vector(2 downto 0);
signal Cin_2_c34, Cin_2_c35 :  std_logic;
signal X_2_c32, X_2_c33, X_2_c34, X_2_c35 :  std_logic_vector(3 downto 0);
signal Y_2_c32, Y_2_c33, Y_2_c34, Y_2_c35 :  std_logic_vector(3 downto 0);
signal S_2_c35 :  std_logic_vector(3 downto 0);
signal R_2_c35, R_2_c36, R_2_c37, R_2_c38 :  std_logic_vector(2 downto 0);
signal Cin_3_c35, Cin_3_c36 :  std_logic;
signal X_3_c32, X_3_c33, X_3_c34, X_3_c35, X_3_c36 :  std_logic_vector(3 downto 0);
signal Y_3_c32, Y_3_c33, Y_3_c34, Y_3_c35, Y_3_c36 :  std_logic_vector(3 downto 0);
signal S_3_c36 :  std_logic_vector(3 downto 0);
signal R_3_c36, R_3_c37, R_3_c38 :  std_logic_vector(2 downto 0);
signal Cin_4_c36, Cin_4_c37 :  std_logic;
signal X_4_c32, X_4_c33, X_4_c34, X_4_c35, X_4_c36, X_4_c37 :  std_logic_vector(3 downto 0);
signal Y_4_c32, Y_4_c33, Y_4_c34, Y_4_c35, Y_4_c36, Y_4_c37 :  std_logic_vector(3 downto 0);
signal S_4_c37 :  std_logic_vector(3 downto 0);
signal R_4_c37, R_4_c38 :  std_logic_vector(2 downto 0);
signal Cin_5_c37, Cin_5_c38 :  std_logic;
signal X_5_c32, X_5_c33, X_5_c34, X_5_c35, X_5_c36, X_5_c37, X_5_c38 :  std_logic_vector(3 downto 0);
signal Y_5_c32, Y_5_c33, Y_5_c34, Y_5_c35, Y_5_c36, Y_5_c37, Y_5_c38 :  std_logic_vector(3 downto 0);
signal S_5_c38 :  std_logic_vector(3 downto 0);
signal R_5_c38 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
            end if;
            if ce_4 = '1' then
               Cin_0_c4 <= Cin_0_c3;
            end if;
            if ce_5 = '1' then
               Cin_0_c5 <= Cin_0_c4;
            end if;
            if ce_6 = '1' then
               Cin_0_c6 <= Cin_0_c5;
            end if;
            if ce_7 = '1' then
               Cin_0_c7 <= Cin_0_c6;
            end if;
            if ce_8 = '1' then
               Cin_0_c8 <= Cin_0_c7;
            end if;
            if ce_9 = '1' then
               Cin_0_c9 <= Cin_0_c8;
            end if;
            if ce_10 = '1' then
               Cin_0_c10 <= Cin_0_c9;
            end if;
            if ce_11 = '1' then
               Cin_0_c11 <= Cin_0_c10;
            end if;
            if ce_12 = '1' then
               Cin_0_c12 <= Cin_0_c11;
            end if;
            if ce_13 = '1' then
               Cin_0_c13 <= Cin_0_c12;
            end if;
            if ce_14 = '1' then
               Cin_0_c14 <= Cin_0_c13;
            end if;
            if ce_15 = '1' then
               Cin_0_c15 <= Cin_0_c14;
            end if;
            if ce_16 = '1' then
               Cin_0_c16 <= Cin_0_c15;
            end if;
            if ce_17 = '1' then
               Cin_0_c17 <= Cin_0_c16;
            end if;
            if ce_18 = '1' then
               Cin_0_c18 <= Cin_0_c17;
            end if;
            if ce_19 = '1' then
               Cin_0_c19 <= Cin_0_c18;
            end if;
            if ce_20 = '1' then
               Cin_0_c20 <= Cin_0_c19;
            end if;
            if ce_21 = '1' then
               Cin_0_c21 <= Cin_0_c20;
            end if;
            if ce_22 = '1' then
               Cin_0_c22 <= Cin_0_c21;
            end if;
            if ce_23 = '1' then
               Cin_0_c23 <= Cin_0_c22;
            end if;
            if ce_24 = '1' then
               Cin_0_c24 <= Cin_0_c23;
            end if;
            if ce_25 = '1' then
               Cin_0_c25 <= Cin_0_c24;
            end if;
            if ce_26 = '1' then
               Cin_0_c26 <= Cin_0_c25;
            end if;
            if ce_27 = '1' then
               Cin_0_c27 <= Cin_0_c26;
            end if;
            if ce_28 = '1' then
               Cin_0_c28 <= Cin_0_c27;
            end if;
            if ce_29 = '1' then
               Cin_0_c29 <= Cin_0_c28;
            end if;
            if ce_30 = '1' then
               Cin_0_c30 <= Cin_0_c29;
            end if;
            if ce_31 = '1' then
               Cin_0_c31 <= Cin_0_c30;
            end if;
            if ce_32 = '1' then
               Cin_0_c32 <= Cin_0_c31;
            end if;
            if ce_33 = '1' then
               Cin_0_c33 <= Cin_0_c32;
               X_0_c33 <= X_0_c32;
               Y_0_c33 <= Y_0_c32;
               X_1_c33 <= X_1_c32;
               Y_1_c33 <= Y_1_c32;
               X_2_c33 <= X_2_c32;
               Y_2_c33 <= Y_2_c32;
               X_3_c33 <= X_3_c32;
               Y_3_c33 <= Y_3_c32;
               X_4_c33 <= X_4_c32;
               Y_4_c33 <= Y_4_c32;
               X_5_c33 <= X_5_c32;
               Y_5_c33 <= Y_5_c32;
            end if;
            if ce_34 = '1' then
               R_0_c34 <= R_0_c33;
               Cin_1_c34 <= Cin_1_c33;
               X_1_c34 <= X_1_c33;
               Y_1_c34 <= Y_1_c33;
               X_2_c34 <= X_2_c33;
               Y_2_c34 <= Y_2_c33;
               X_3_c34 <= X_3_c33;
               Y_3_c34 <= Y_3_c33;
               X_4_c34 <= X_4_c33;
               Y_4_c34 <= Y_4_c33;
               X_5_c34 <= X_5_c33;
               Y_5_c34 <= Y_5_c33;
            end if;
            if ce_35 = '1' then
               R_0_c35 <= R_0_c34;
               R_1_c35 <= R_1_c34;
               Cin_2_c35 <= Cin_2_c34;
               X_2_c35 <= X_2_c34;
               Y_2_c35 <= Y_2_c34;
               X_3_c35 <= X_3_c34;
               Y_3_c35 <= Y_3_c34;
               X_4_c35 <= X_4_c34;
               Y_4_c35 <= Y_4_c34;
               X_5_c35 <= X_5_c34;
               Y_5_c35 <= Y_5_c34;
            end if;
            if ce_36 = '1' then
               R_0_c36 <= R_0_c35;
               R_1_c36 <= R_1_c35;
               R_2_c36 <= R_2_c35;
               Cin_3_c36 <= Cin_3_c35;
               X_3_c36 <= X_3_c35;
               Y_3_c36 <= Y_3_c35;
               X_4_c36 <= X_4_c35;
               Y_4_c36 <= Y_4_c35;
               X_5_c36 <= X_5_c35;
               Y_5_c36 <= Y_5_c35;
            end if;
            if ce_37 = '1' then
               R_0_c37 <= R_0_c36;
               R_1_c37 <= R_1_c36;
               R_2_c37 <= R_2_c36;
               R_3_c37 <= R_3_c36;
               Cin_4_c37 <= Cin_4_c36;
               X_4_c37 <= X_4_c36;
               Y_4_c37 <= Y_4_c36;
               X_5_c37 <= X_5_c36;
               Y_5_c37 <= Y_5_c36;
            end if;
            if ce_38 = '1' then
               R_0_c38 <= R_0_c37;
               R_1_c38 <= R_1_c37;
               R_2_c38 <= R_2_c37;
               R_3_c38 <= R_3_c37;
               R_4_c38 <= R_4_c37;
               Cin_5_c38 <= Cin_5_c37;
               X_5_c38 <= X_5_c37;
               Y_5_c38 <= Y_5_c37;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c32 <= '0' & X(2 downto 0);
   Y_0_c32 <= '0' & Y(2 downto 0);
   S_0_c33 <= X_0_c33 + Y_0_c33 + Cin_0_c33;
   R_0_c33 <= S_0_c33(2 downto 0);
   Cin_1_c33 <= S_0_c33(3);
   X_1_c32 <= '0' & X(5 downto 3);
   Y_1_c32 <= '0' & Y(5 downto 3);
   S_1_c34 <= X_1_c34 + Y_1_c34 + Cin_1_c34;
   R_1_c34 <= S_1_c34(2 downto 0);
   Cin_2_c34 <= S_1_c34(3);
   X_2_c32 <= '0' & X(8 downto 6);
   Y_2_c32 <= '0' & Y(8 downto 6);
   S_2_c35 <= X_2_c35 + Y_2_c35 + Cin_2_c35;
   R_2_c35 <= S_2_c35(2 downto 0);
   Cin_3_c35 <= S_2_c35(3);
   X_3_c32 <= '0' & X(11 downto 9);
   Y_3_c32 <= '0' & Y(11 downto 9);
   S_3_c36 <= X_3_c36 + Y_3_c36 + Cin_3_c36;
   R_3_c36 <= S_3_c36(2 downto 0);
   Cin_4_c36 <= S_3_c36(3);
   X_4_c32 <= '0' & X(14 downto 12);
   Y_4_c32 <= '0' & Y(14 downto 12);
   S_4_c37 <= X_4_c37 + Y_4_c37 + Cin_4_c37;
   R_4_c37 <= S_4_c37(2 downto 0);
   Cin_5_c37 <= S_4_c37(3);
   X_5_c32 <= '0' & X(17 downto 15);
   Y_5_c32 <= '0' & Y(17 downto 15);
   S_5_c38 <= X_5_c38 + Y_5_c38 + Cin_5_c38;
   R_5_c38 <= S_5_c38(2 downto 0);
   R <= R_5_c38 & R_4_c38 & R_3_c38 & R_2_c38 & R_1_c38 & R_0_c38 ;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_18_Freq800_uid52
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 41 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_18_Freq800_uid52 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(17 downto 0);
          Y : in  std_logic_vector(17 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of IntAdder_18_Freq800_uid52 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3, Cin_0_c4, Cin_0_c5, Cin_0_c6, Cin_0_c7, Cin_0_c8, Cin_0_c9, Cin_0_c10, Cin_0_c11, Cin_0_c12, Cin_0_c13, Cin_0_c14, Cin_0_c15, Cin_0_c16, Cin_0_c17, Cin_0_c18, Cin_0_c19, Cin_0_c20, Cin_0_c21, Cin_0_c22, Cin_0_c23, Cin_0_c24, Cin_0_c25, Cin_0_c26, Cin_0_c27, Cin_0_c28, Cin_0_c29, Cin_0_c30, Cin_0_c31, Cin_0_c32, Cin_0_c33, Cin_0_c34, Cin_0_c35, Cin_0_c36 :  std_logic;
signal X_0_c35, X_0_c36 :  std_logic_vector(3 downto 0);
signal Y_0_c0, Y_0_c1, Y_0_c2, Y_0_c3, Y_0_c4, Y_0_c5, Y_0_c6, Y_0_c7, Y_0_c8, Y_0_c9, Y_0_c10, Y_0_c11, Y_0_c12, Y_0_c13, Y_0_c14, Y_0_c15, Y_0_c16, Y_0_c17, Y_0_c18, Y_0_c19, Y_0_c20, Y_0_c21, Y_0_c22, Y_0_c23, Y_0_c24, Y_0_c25, Y_0_c26, Y_0_c27, Y_0_c28, Y_0_c29, Y_0_c30, Y_0_c31, Y_0_c32, Y_0_c33, Y_0_c34, Y_0_c35, Y_0_c36 :  std_logic_vector(3 downto 0);
signal S_0_c36 :  std_logic_vector(3 downto 0);
signal R_0_c36, R_0_c37, R_0_c38, R_0_c39, R_0_c40, R_0_c41 :  std_logic_vector(2 downto 0);
signal Cin_1_c36, Cin_1_c37 :  std_logic;
signal X_1_c35, X_1_c36, X_1_c37 :  std_logic_vector(3 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3, Y_1_c4, Y_1_c5, Y_1_c6, Y_1_c7, Y_1_c8, Y_1_c9, Y_1_c10, Y_1_c11, Y_1_c12, Y_1_c13, Y_1_c14, Y_1_c15, Y_1_c16, Y_1_c17, Y_1_c18, Y_1_c19, Y_1_c20, Y_1_c21, Y_1_c22, Y_1_c23, Y_1_c24, Y_1_c25, Y_1_c26, Y_1_c27, Y_1_c28, Y_1_c29, Y_1_c30, Y_1_c31, Y_1_c32, Y_1_c33, Y_1_c34, Y_1_c35, Y_1_c36, Y_1_c37 :  std_logic_vector(3 downto 0);
signal S_1_c37 :  std_logic_vector(3 downto 0);
signal R_1_c37, R_1_c38, R_1_c39, R_1_c40, R_1_c41 :  std_logic_vector(2 downto 0);
signal Cin_2_c37, Cin_2_c38 :  std_logic;
signal X_2_c35, X_2_c36, X_2_c37, X_2_c38 :  std_logic_vector(3 downto 0);
signal Y_2_c0, Y_2_c1, Y_2_c2, Y_2_c3, Y_2_c4, Y_2_c5, Y_2_c6, Y_2_c7, Y_2_c8, Y_2_c9, Y_2_c10, Y_2_c11, Y_2_c12, Y_2_c13, Y_2_c14, Y_2_c15, Y_2_c16, Y_2_c17, Y_2_c18, Y_2_c19, Y_2_c20, Y_2_c21, Y_2_c22, Y_2_c23, Y_2_c24, Y_2_c25, Y_2_c26, Y_2_c27, Y_2_c28, Y_2_c29, Y_2_c30, Y_2_c31, Y_2_c32, Y_2_c33, Y_2_c34, Y_2_c35, Y_2_c36, Y_2_c37, Y_2_c38 :  std_logic_vector(3 downto 0);
signal S_2_c38 :  std_logic_vector(3 downto 0);
signal R_2_c38, R_2_c39, R_2_c40, R_2_c41 :  std_logic_vector(2 downto 0);
signal Cin_3_c38, Cin_3_c39 :  std_logic;
signal X_3_c35, X_3_c36, X_3_c37, X_3_c38, X_3_c39 :  std_logic_vector(3 downto 0);
signal Y_3_c0, Y_3_c1, Y_3_c2, Y_3_c3, Y_3_c4, Y_3_c5, Y_3_c6, Y_3_c7, Y_3_c8, Y_3_c9, Y_3_c10, Y_3_c11, Y_3_c12, Y_3_c13, Y_3_c14, Y_3_c15, Y_3_c16, Y_3_c17, Y_3_c18, Y_3_c19, Y_3_c20, Y_3_c21, Y_3_c22, Y_3_c23, Y_3_c24, Y_3_c25, Y_3_c26, Y_3_c27, Y_3_c28, Y_3_c29, Y_3_c30, Y_3_c31, Y_3_c32, Y_3_c33, Y_3_c34, Y_3_c35, Y_3_c36, Y_3_c37, Y_3_c38, Y_3_c39 :  std_logic_vector(3 downto 0);
signal S_3_c39 :  std_logic_vector(3 downto 0);
signal R_3_c39, R_3_c40, R_3_c41 :  std_logic_vector(2 downto 0);
signal Cin_4_c39, Cin_4_c40 :  std_logic;
signal X_4_c35, X_4_c36, X_4_c37, X_4_c38, X_4_c39, X_4_c40 :  std_logic_vector(3 downto 0);
signal Y_4_c0, Y_4_c1, Y_4_c2, Y_4_c3, Y_4_c4, Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8, Y_4_c9, Y_4_c10, Y_4_c11, Y_4_c12, Y_4_c13, Y_4_c14, Y_4_c15, Y_4_c16, Y_4_c17, Y_4_c18, Y_4_c19, Y_4_c20, Y_4_c21, Y_4_c22, Y_4_c23, Y_4_c24, Y_4_c25, Y_4_c26, Y_4_c27, Y_4_c28, Y_4_c29, Y_4_c30, Y_4_c31, Y_4_c32, Y_4_c33, Y_4_c34, Y_4_c35, Y_4_c36, Y_4_c37, Y_4_c38, Y_4_c39, Y_4_c40 :  std_logic_vector(3 downto 0);
signal S_4_c40 :  std_logic_vector(3 downto 0);
signal R_4_c40, R_4_c41 :  std_logic_vector(2 downto 0);
signal Cin_5_c40, Cin_5_c41 :  std_logic;
signal X_5_c35, X_5_c36, X_5_c37, X_5_c38, X_5_c39, X_5_c40, X_5_c41 :  std_logic_vector(3 downto 0);
signal Y_5_c0, Y_5_c1, Y_5_c2, Y_5_c3, Y_5_c4, Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9, Y_5_c10, Y_5_c11, Y_5_c12, Y_5_c13, Y_5_c14, Y_5_c15, Y_5_c16, Y_5_c17, Y_5_c18, Y_5_c19, Y_5_c20, Y_5_c21, Y_5_c22, Y_5_c23, Y_5_c24, Y_5_c25, Y_5_c26, Y_5_c27, Y_5_c28, Y_5_c29, Y_5_c30, Y_5_c31, Y_5_c32, Y_5_c33, Y_5_c34, Y_5_c35, Y_5_c36, Y_5_c37, Y_5_c38, Y_5_c39, Y_5_c40, Y_5_c41 :  std_logic_vector(3 downto 0);
signal S_5_c41 :  std_logic_vector(3 downto 0);
signal R_5_c41 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
               Y_0_c1 <= Y_0_c0;
               Y_1_c1 <= Y_1_c0;
               Y_2_c1 <= Y_2_c0;
               Y_3_c1 <= Y_3_c0;
               Y_4_c1 <= Y_4_c0;
               Y_5_c1 <= Y_5_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
               Y_0_c2 <= Y_0_c1;
               Y_1_c2 <= Y_1_c1;
               Y_2_c2 <= Y_2_c1;
               Y_3_c2 <= Y_3_c1;
               Y_4_c2 <= Y_4_c1;
               Y_5_c2 <= Y_5_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
               Y_0_c3 <= Y_0_c2;
               Y_1_c3 <= Y_1_c2;
               Y_2_c3 <= Y_2_c2;
               Y_3_c3 <= Y_3_c2;
               Y_4_c3 <= Y_4_c2;
               Y_5_c3 <= Y_5_c2;
            end if;
            if ce_4 = '1' then
               Cin_0_c4 <= Cin_0_c3;
               Y_0_c4 <= Y_0_c3;
               Y_1_c4 <= Y_1_c3;
               Y_2_c4 <= Y_2_c3;
               Y_3_c4 <= Y_3_c3;
               Y_4_c4 <= Y_4_c3;
               Y_5_c4 <= Y_5_c3;
            end if;
            if ce_5 = '1' then
               Cin_0_c5 <= Cin_0_c4;
               Y_0_c5 <= Y_0_c4;
               Y_1_c5 <= Y_1_c4;
               Y_2_c5 <= Y_2_c4;
               Y_3_c5 <= Y_3_c4;
               Y_4_c5 <= Y_4_c4;
               Y_5_c5 <= Y_5_c4;
            end if;
            if ce_6 = '1' then
               Cin_0_c6 <= Cin_0_c5;
               Y_0_c6 <= Y_0_c5;
               Y_1_c6 <= Y_1_c5;
               Y_2_c6 <= Y_2_c5;
               Y_3_c6 <= Y_3_c5;
               Y_4_c6 <= Y_4_c5;
               Y_5_c6 <= Y_5_c5;
            end if;
            if ce_7 = '1' then
               Cin_0_c7 <= Cin_0_c6;
               Y_0_c7 <= Y_0_c6;
               Y_1_c7 <= Y_1_c6;
               Y_2_c7 <= Y_2_c6;
               Y_3_c7 <= Y_3_c6;
               Y_4_c7 <= Y_4_c6;
               Y_5_c7 <= Y_5_c6;
            end if;
            if ce_8 = '1' then
               Cin_0_c8 <= Cin_0_c7;
               Y_0_c8 <= Y_0_c7;
               Y_1_c8 <= Y_1_c7;
               Y_2_c8 <= Y_2_c7;
               Y_3_c8 <= Y_3_c7;
               Y_4_c8 <= Y_4_c7;
               Y_5_c8 <= Y_5_c7;
            end if;
            if ce_9 = '1' then
               Cin_0_c9 <= Cin_0_c8;
               Y_0_c9 <= Y_0_c8;
               Y_1_c9 <= Y_1_c8;
               Y_2_c9 <= Y_2_c8;
               Y_3_c9 <= Y_3_c8;
               Y_4_c9 <= Y_4_c8;
               Y_5_c9 <= Y_5_c8;
            end if;
            if ce_10 = '1' then
               Cin_0_c10 <= Cin_0_c9;
               Y_0_c10 <= Y_0_c9;
               Y_1_c10 <= Y_1_c9;
               Y_2_c10 <= Y_2_c9;
               Y_3_c10 <= Y_3_c9;
               Y_4_c10 <= Y_4_c9;
               Y_5_c10 <= Y_5_c9;
            end if;
            if ce_11 = '1' then
               Cin_0_c11 <= Cin_0_c10;
               Y_0_c11 <= Y_0_c10;
               Y_1_c11 <= Y_1_c10;
               Y_2_c11 <= Y_2_c10;
               Y_3_c11 <= Y_3_c10;
               Y_4_c11 <= Y_4_c10;
               Y_5_c11 <= Y_5_c10;
            end if;
            if ce_12 = '1' then
               Cin_0_c12 <= Cin_0_c11;
               Y_0_c12 <= Y_0_c11;
               Y_1_c12 <= Y_1_c11;
               Y_2_c12 <= Y_2_c11;
               Y_3_c12 <= Y_3_c11;
               Y_4_c12 <= Y_4_c11;
               Y_5_c12 <= Y_5_c11;
            end if;
            if ce_13 = '1' then
               Cin_0_c13 <= Cin_0_c12;
               Y_0_c13 <= Y_0_c12;
               Y_1_c13 <= Y_1_c12;
               Y_2_c13 <= Y_2_c12;
               Y_3_c13 <= Y_3_c12;
               Y_4_c13 <= Y_4_c12;
               Y_5_c13 <= Y_5_c12;
            end if;
            if ce_14 = '1' then
               Cin_0_c14 <= Cin_0_c13;
               Y_0_c14 <= Y_0_c13;
               Y_1_c14 <= Y_1_c13;
               Y_2_c14 <= Y_2_c13;
               Y_3_c14 <= Y_3_c13;
               Y_4_c14 <= Y_4_c13;
               Y_5_c14 <= Y_5_c13;
            end if;
            if ce_15 = '1' then
               Cin_0_c15 <= Cin_0_c14;
               Y_0_c15 <= Y_0_c14;
               Y_1_c15 <= Y_1_c14;
               Y_2_c15 <= Y_2_c14;
               Y_3_c15 <= Y_3_c14;
               Y_4_c15 <= Y_4_c14;
               Y_5_c15 <= Y_5_c14;
            end if;
            if ce_16 = '1' then
               Cin_0_c16 <= Cin_0_c15;
               Y_0_c16 <= Y_0_c15;
               Y_1_c16 <= Y_1_c15;
               Y_2_c16 <= Y_2_c15;
               Y_3_c16 <= Y_3_c15;
               Y_4_c16 <= Y_4_c15;
               Y_5_c16 <= Y_5_c15;
            end if;
            if ce_17 = '1' then
               Cin_0_c17 <= Cin_0_c16;
               Y_0_c17 <= Y_0_c16;
               Y_1_c17 <= Y_1_c16;
               Y_2_c17 <= Y_2_c16;
               Y_3_c17 <= Y_3_c16;
               Y_4_c17 <= Y_4_c16;
               Y_5_c17 <= Y_5_c16;
            end if;
            if ce_18 = '1' then
               Cin_0_c18 <= Cin_0_c17;
               Y_0_c18 <= Y_0_c17;
               Y_1_c18 <= Y_1_c17;
               Y_2_c18 <= Y_2_c17;
               Y_3_c18 <= Y_3_c17;
               Y_4_c18 <= Y_4_c17;
               Y_5_c18 <= Y_5_c17;
            end if;
            if ce_19 = '1' then
               Cin_0_c19 <= Cin_0_c18;
               Y_0_c19 <= Y_0_c18;
               Y_1_c19 <= Y_1_c18;
               Y_2_c19 <= Y_2_c18;
               Y_3_c19 <= Y_3_c18;
               Y_4_c19 <= Y_4_c18;
               Y_5_c19 <= Y_5_c18;
            end if;
            if ce_20 = '1' then
               Cin_0_c20 <= Cin_0_c19;
               Y_0_c20 <= Y_0_c19;
               Y_1_c20 <= Y_1_c19;
               Y_2_c20 <= Y_2_c19;
               Y_3_c20 <= Y_3_c19;
               Y_4_c20 <= Y_4_c19;
               Y_5_c20 <= Y_5_c19;
            end if;
            if ce_21 = '1' then
               Cin_0_c21 <= Cin_0_c20;
               Y_0_c21 <= Y_0_c20;
               Y_1_c21 <= Y_1_c20;
               Y_2_c21 <= Y_2_c20;
               Y_3_c21 <= Y_3_c20;
               Y_4_c21 <= Y_4_c20;
               Y_5_c21 <= Y_5_c20;
            end if;
            if ce_22 = '1' then
               Cin_0_c22 <= Cin_0_c21;
               Y_0_c22 <= Y_0_c21;
               Y_1_c22 <= Y_1_c21;
               Y_2_c22 <= Y_2_c21;
               Y_3_c22 <= Y_3_c21;
               Y_4_c22 <= Y_4_c21;
               Y_5_c22 <= Y_5_c21;
            end if;
            if ce_23 = '1' then
               Cin_0_c23 <= Cin_0_c22;
               Y_0_c23 <= Y_0_c22;
               Y_1_c23 <= Y_1_c22;
               Y_2_c23 <= Y_2_c22;
               Y_3_c23 <= Y_3_c22;
               Y_4_c23 <= Y_4_c22;
               Y_5_c23 <= Y_5_c22;
            end if;
            if ce_24 = '1' then
               Cin_0_c24 <= Cin_0_c23;
               Y_0_c24 <= Y_0_c23;
               Y_1_c24 <= Y_1_c23;
               Y_2_c24 <= Y_2_c23;
               Y_3_c24 <= Y_3_c23;
               Y_4_c24 <= Y_4_c23;
               Y_5_c24 <= Y_5_c23;
            end if;
            if ce_25 = '1' then
               Cin_0_c25 <= Cin_0_c24;
               Y_0_c25 <= Y_0_c24;
               Y_1_c25 <= Y_1_c24;
               Y_2_c25 <= Y_2_c24;
               Y_3_c25 <= Y_3_c24;
               Y_4_c25 <= Y_4_c24;
               Y_5_c25 <= Y_5_c24;
            end if;
            if ce_26 = '1' then
               Cin_0_c26 <= Cin_0_c25;
               Y_0_c26 <= Y_0_c25;
               Y_1_c26 <= Y_1_c25;
               Y_2_c26 <= Y_2_c25;
               Y_3_c26 <= Y_3_c25;
               Y_4_c26 <= Y_4_c25;
               Y_5_c26 <= Y_5_c25;
            end if;
            if ce_27 = '1' then
               Cin_0_c27 <= Cin_0_c26;
               Y_0_c27 <= Y_0_c26;
               Y_1_c27 <= Y_1_c26;
               Y_2_c27 <= Y_2_c26;
               Y_3_c27 <= Y_3_c26;
               Y_4_c27 <= Y_4_c26;
               Y_5_c27 <= Y_5_c26;
            end if;
            if ce_28 = '1' then
               Cin_0_c28 <= Cin_0_c27;
               Y_0_c28 <= Y_0_c27;
               Y_1_c28 <= Y_1_c27;
               Y_2_c28 <= Y_2_c27;
               Y_3_c28 <= Y_3_c27;
               Y_4_c28 <= Y_4_c27;
               Y_5_c28 <= Y_5_c27;
            end if;
            if ce_29 = '1' then
               Cin_0_c29 <= Cin_0_c28;
               Y_0_c29 <= Y_0_c28;
               Y_1_c29 <= Y_1_c28;
               Y_2_c29 <= Y_2_c28;
               Y_3_c29 <= Y_3_c28;
               Y_4_c29 <= Y_4_c28;
               Y_5_c29 <= Y_5_c28;
            end if;
            if ce_30 = '1' then
               Cin_0_c30 <= Cin_0_c29;
               Y_0_c30 <= Y_0_c29;
               Y_1_c30 <= Y_1_c29;
               Y_2_c30 <= Y_2_c29;
               Y_3_c30 <= Y_3_c29;
               Y_4_c30 <= Y_4_c29;
               Y_5_c30 <= Y_5_c29;
            end if;
            if ce_31 = '1' then
               Cin_0_c31 <= Cin_0_c30;
               Y_0_c31 <= Y_0_c30;
               Y_1_c31 <= Y_1_c30;
               Y_2_c31 <= Y_2_c30;
               Y_3_c31 <= Y_3_c30;
               Y_4_c31 <= Y_4_c30;
               Y_5_c31 <= Y_5_c30;
            end if;
            if ce_32 = '1' then
               Cin_0_c32 <= Cin_0_c31;
               Y_0_c32 <= Y_0_c31;
               Y_1_c32 <= Y_1_c31;
               Y_2_c32 <= Y_2_c31;
               Y_3_c32 <= Y_3_c31;
               Y_4_c32 <= Y_4_c31;
               Y_5_c32 <= Y_5_c31;
            end if;
            if ce_33 = '1' then
               Cin_0_c33 <= Cin_0_c32;
               Y_0_c33 <= Y_0_c32;
               Y_1_c33 <= Y_1_c32;
               Y_2_c33 <= Y_2_c32;
               Y_3_c33 <= Y_3_c32;
               Y_4_c33 <= Y_4_c32;
               Y_5_c33 <= Y_5_c32;
            end if;
            if ce_34 = '1' then
               Cin_0_c34 <= Cin_0_c33;
               Y_0_c34 <= Y_0_c33;
               Y_1_c34 <= Y_1_c33;
               Y_2_c34 <= Y_2_c33;
               Y_3_c34 <= Y_3_c33;
               Y_4_c34 <= Y_4_c33;
               Y_5_c34 <= Y_5_c33;
            end if;
            if ce_35 = '1' then
               Cin_0_c35 <= Cin_0_c34;
               Y_0_c35 <= Y_0_c34;
               Y_1_c35 <= Y_1_c34;
               Y_2_c35 <= Y_2_c34;
               Y_3_c35 <= Y_3_c34;
               Y_4_c35 <= Y_4_c34;
               Y_5_c35 <= Y_5_c34;
            end if;
            if ce_36 = '1' then
               Cin_0_c36 <= Cin_0_c35;
               X_0_c36 <= X_0_c35;
               Y_0_c36 <= Y_0_c35;
               X_1_c36 <= X_1_c35;
               Y_1_c36 <= Y_1_c35;
               X_2_c36 <= X_2_c35;
               Y_2_c36 <= Y_2_c35;
               X_3_c36 <= X_3_c35;
               Y_3_c36 <= Y_3_c35;
               X_4_c36 <= X_4_c35;
               Y_4_c36 <= Y_4_c35;
               X_5_c36 <= X_5_c35;
               Y_5_c36 <= Y_5_c35;
            end if;
            if ce_37 = '1' then
               R_0_c37 <= R_0_c36;
               Cin_1_c37 <= Cin_1_c36;
               X_1_c37 <= X_1_c36;
               Y_1_c37 <= Y_1_c36;
               X_2_c37 <= X_2_c36;
               Y_2_c37 <= Y_2_c36;
               X_3_c37 <= X_3_c36;
               Y_3_c37 <= Y_3_c36;
               X_4_c37 <= X_4_c36;
               Y_4_c37 <= Y_4_c36;
               X_5_c37 <= X_5_c36;
               Y_5_c37 <= Y_5_c36;
            end if;
            if ce_38 = '1' then
               R_0_c38 <= R_0_c37;
               R_1_c38 <= R_1_c37;
               Cin_2_c38 <= Cin_2_c37;
               X_2_c38 <= X_2_c37;
               Y_2_c38 <= Y_2_c37;
               X_3_c38 <= X_3_c37;
               Y_3_c38 <= Y_3_c37;
               X_4_c38 <= X_4_c37;
               Y_4_c38 <= Y_4_c37;
               X_5_c38 <= X_5_c37;
               Y_5_c38 <= Y_5_c37;
            end if;
            if ce_39 = '1' then
               R_0_c39 <= R_0_c38;
               R_1_c39 <= R_1_c38;
               R_2_c39 <= R_2_c38;
               Cin_3_c39 <= Cin_3_c38;
               X_3_c39 <= X_3_c38;
               Y_3_c39 <= Y_3_c38;
               X_4_c39 <= X_4_c38;
               Y_4_c39 <= Y_4_c38;
               X_5_c39 <= X_5_c38;
               Y_5_c39 <= Y_5_c38;
            end if;
            if ce_40 = '1' then
               R_0_c40 <= R_0_c39;
               R_1_c40 <= R_1_c39;
               R_2_c40 <= R_2_c39;
               R_3_c40 <= R_3_c39;
               Cin_4_c40 <= Cin_4_c39;
               X_4_c40 <= X_4_c39;
               Y_4_c40 <= Y_4_c39;
               X_5_c40 <= X_5_c39;
               Y_5_c40 <= Y_5_c39;
            end if;
            if ce_41 = '1' then
               R_0_c41 <= R_0_c40;
               R_1_c41 <= R_1_c40;
               R_2_c41 <= R_2_c40;
               R_3_c41 <= R_3_c40;
               R_4_c41 <= R_4_c40;
               Cin_5_c41 <= Cin_5_c40;
               X_5_c41 <= X_5_c40;
               Y_5_c41 <= Y_5_c40;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c35 <= '0' & X(2 downto 0);
   Y_0_c0 <= '0' & Y(2 downto 0);
   S_0_c36 <= X_0_c36 + Y_0_c36 + Cin_0_c36;
   R_0_c36 <= S_0_c36(2 downto 0);
   Cin_1_c36 <= S_0_c36(3);
   X_1_c35 <= '0' & X(5 downto 3);
   Y_1_c0 <= '0' & Y(5 downto 3);
   S_1_c37 <= X_1_c37 + Y_1_c37 + Cin_1_c37;
   R_1_c37 <= S_1_c37(2 downto 0);
   Cin_2_c37 <= S_1_c37(3);
   X_2_c35 <= '0' & X(8 downto 6);
   Y_2_c0 <= '0' & Y(8 downto 6);
   S_2_c38 <= X_2_c38 + Y_2_c38 + Cin_2_c38;
   R_2_c38 <= S_2_c38(2 downto 0);
   Cin_3_c38 <= S_2_c38(3);
   X_3_c35 <= '0' & X(11 downto 9);
   Y_3_c0 <= '0' & Y(11 downto 9);
   S_3_c39 <= X_3_c39 + Y_3_c39 + Cin_3_c39;
   R_3_c39 <= S_3_c39(2 downto 0);
   Cin_4_c39 <= S_3_c39(3);
   X_4_c35 <= '0' & X(14 downto 12);
   Y_4_c0 <= '0' & Y(14 downto 12);
   S_4_c40 <= X_4_c40 + Y_4_c40 + Cin_4_c40;
   R_4_c40 <= S_4_c40(2 downto 0);
   Cin_5_c40 <= S_4_c40(3);
   X_5_c35 <= '0' & X(17 downto 15);
   Y_5_c0 <= '0' & Y(17 downto 15);
   S_5_c41 <= X_5_c41 + Y_5_c41 + Cin_5_c41;
   R_5_c41 <= S_5_c41(2 downto 0);
   R <= R_5_c41 & R_4_c41 & R_3_c41 & R_2_c41 & R_1_c41 & R_0_c41 ;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x1_Freq800_uid58
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid58 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid58 is
signal replicated_c41 :  std_logic_vector(0 downto 0);
signal prod_c41 :  std_logic_vector(0 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
   replicated_c41 <= (0 downto 0 => X(0));
   prod_c41 <= Y_c41 and replicated_c41;
   R <= prod_c41;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x2_Freq800_uid60
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid60 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid60 is
   component MultTable_Freq800_uid62 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(3 downto 0);
signal Y1_c41 :  std_logic_vector(3 downto 0);
signal Y1_copy63_c41 :  std_logic_vector(3 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid62
      port map ( X => Xtable_c41,
                 Y => Y1_copy63_c41);
   Y1_c41 <= Y1_copy63_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid65
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid65 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid65 is
   component MultTable_Freq800_uid67 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy68_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid67
      port map ( X => Xtable_c41,
                 Y => Y1_copy68_c41);
   Y1_c41 <= Y1_copy68_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x1_Freq800_uid70
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid70 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid70 is
signal replicated_c41 :  std_logic_vector(0 downto 0);
signal prod_c41 :  std_logic_vector(0 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
   replicated_c41 <= (0 downto 0 => X(0));
   prod_c41 <= Y_c41 and replicated_c41;
   R <= prod_c41;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x1_Freq800_uid72
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq800_uid72 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq800_uid72 is
signal replicated_c38, replicated_c39, replicated_c40, replicated_c41 :  std_logic_vector(1 downto 0);
signal prod_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               replicated_c39 <= replicated_c38;
            end if;
            if ce_40 = '1' then
               replicated_c40 <= replicated_c39;
            end if;
            if ce_41 = '1' then
               replicated_c41 <= replicated_c40;
            end if;
         end if;
      end process;
   replicated_c38 <= (1 downto 0 => Y(0));
   prod_c41 <= X and replicated_c41;
   R <= prod_c41;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid74
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid74 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid74 is
   component MultTable_Freq800_uid76 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy77_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid76
      port map ( X => Xtable_c41,
                 Y => Y1_copy77_c41);
   Y1_c41 <= Y1_copy77_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid79
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid79 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid79 is
   component MultTable_Freq800_uid81 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy82_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid81
      port map ( X => Xtable_c41,
                 Y => Y1_copy82_c41);
   Y1_c41 <= Y1_copy82_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x1_Freq800_uid84
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid84 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid84 is
signal replicated_c41 :  std_logic_vector(0 downto 0);
signal prod_c41 :  std_logic_vector(0 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
   replicated_c41 <= (0 downto 0 => X(0));
   prod_c41 <= Y_c41 and replicated_c41;
   R <= prod_c41;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid86
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid86 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid86 is
   component MultTable_Freq800_uid88 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy89_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid88
      port map ( X => Xtable_c41,
                 Y => Y1_copy89_c41);
   Y1_c41 <= Y1_copy89_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid91
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid91 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid91 is
   component MultTable_Freq800_uid93 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy94_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid93
      port map ( X => Xtable_c41,
                 Y => Y1_copy94_c41);
   Y1_c41 <= Y1_copy94_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid96
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid96 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid96 is
   component MultTable_Freq800_uid98 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy99_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid98
      port map ( X => Xtable_c41,
                 Y => Y1_copy99_c41);
   Y1_c41 <= Y1_copy99_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq800_uid101
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid101 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid101 is
signal replicated_c41 :  std_logic_vector(0 downto 0);
signal prod_c41 :  std_logic_vector(0 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
   replicated_c41 <= (0 downto 0 => X(0));
   prod_c41 <= Y_c41 and replicated_c41;
   R <= prod_c41;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid103
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid103 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid103 is
   component MultTable_Freq800_uid105 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(3 downto 0);
signal Y1_c41 :  std_logic_vector(3 downto 0);
signal Y1_copy106_c41 :  std_logic_vector(3 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid105
      port map ( X => Xtable_c41,
                 Y => Y1_copy106_c41);
   Y1_c41 <= Y1_copy106_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid108
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid108 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid108 is
   component MultTable_Freq800_uid110 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy111_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid110
      port map ( X => Xtable_c41,
                 Y => Y1_copy111_c41);
   Y1_c41 <= Y1_copy111_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid113
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid113 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid113 is
   component MultTable_Freq800_uid115 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy116_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid115
      port map ( X => Xtable_c41,
                 Y => Y1_copy116_c41);
   Y1_c41 <= Y1_copy116_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid118
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid118 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid118 is
   component MultTable_Freq800_uid120 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy121_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid120
      port map ( X => Xtable_c41,
                 Y => Y1_copy121_c41);
   Y1_c41 <= Y1_copy121_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq800_uid123
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid123 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid123 is
signal replicated_c41 :  std_logic_vector(0 downto 0);
signal prod_c41 :  std_logic_vector(0 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
   replicated_c41 <= (0 downto 0 => X(0));
   prod_c41 <= Y_c41 and replicated_c41;
   R <= prod_c41;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x1_Freq800_uid125
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x1_Freq800_uid125 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x1_Freq800_uid125 is
signal replicated_c38, replicated_c39, replicated_c40, replicated_c41 :  std_logic_vector(1 downto 0);
signal prod_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               replicated_c39 <= replicated_c38;
            end if;
            if ce_40 = '1' then
               replicated_c40 <= replicated_c39;
            end if;
            if ce_41 = '1' then
               replicated_c41 <= replicated_c40;
            end if;
         end if;
      end process;
   replicated_c38 <= (1 downto 0 => Y(0));
   prod_c41 <= X and replicated_c41;
   R <= prod_c41;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid127
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid127 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid127 is
   component MultTable_Freq800_uid129 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy130_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid129
      port map ( X => Xtable_c41,
                 Y => Y1_copy130_c41);
   Y1_c41 <= Y1_copy130_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid132
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid132 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid132 is
   component MultTable_Freq800_uid134 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy135_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid134
      port map ( X => Xtable_c41,
                 Y => Y1_copy135_c41);
   Y1_c41 <= Y1_copy135_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid137
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid137 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid137 is
   component MultTable_Freq800_uid139 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy140_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid139
      port map ( X => Xtable_c41,
                 Y => Y1_copy140_c41);
   Y1_c41 <= Y1_copy140_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid142
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid142 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid142 is
   component MultTable_Freq800_uid144 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy145_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid144
      port map ( X => Xtable_c41,
                 Y => Y1_copy145_c41);
   Y1_c41 <= Y1_copy145_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq800_uid147
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid147 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid147 is
signal replicated_c41 :  std_logic_vector(0 downto 0);
signal prod_c41 :  std_logic_vector(0 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
   replicated_c41 <= (0 downto 0 => X(0));
   prod_c41 <= Y_c41 and replicated_c41;
   R <= prod_c41;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid149
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid149 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid149 is
   component MultTable_Freq800_uid151 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy152_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid151
      port map ( X => Xtable_c41,
                 Y => Y1_copy152_c41);
   Y1_c41 <= Y1_copy152_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid154
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid154 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid154 is
   component MultTable_Freq800_uid156 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy157_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid156
      port map ( X => Xtable_c41,
                 Y => Y1_copy157_c41);
   Y1_c41 <= Y1_copy157_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid159
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid159 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid159 is
   component MultTable_Freq800_uid161 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy162_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid161
      port map ( X => Xtable_c41,
                 Y => Y1_copy162_c41);
   Y1_c41 <= Y1_copy162_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid164
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid164 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid164 is
   component MultTable_Freq800_uid166 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy167_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid166
      port map ( X => Xtable_c41,
                 Y => Y1_copy167_c41);
   Y1_c41 <= Y1_copy167_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid169
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid169 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid169 is
   component MultTable_Freq800_uid171 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy172_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid171
      port map ( X => Xtable_c41,
                 Y => Y1_copy172_c41);
   Y1_c41 <= Y1_copy172_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid174
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid174 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid174 is
   component MultTable_Freq800_uid176 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(3 downto 0);
signal Y1_c41 :  std_logic_vector(3 downto 0);
signal Y1_copy177_c41 :  std_logic_vector(3 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid176
      port map ( X => Xtable_c41,
                 Y => Y1_copy177_c41);
   Y1_c41 <= Y1_copy177_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid179
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid179 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid179 is
   component MultTable_Freq800_uid181 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy182_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid181
      port map ( X => Xtable_c41,
                 Y => Y1_copy182_c41);
   Y1_c41 <= Y1_copy182_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid184
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid184 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid184 is
   component MultTable_Freq800_uid186 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy187_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid186
      port map ( X => Xtable_c41,
                 Y => Y1_copy187_c41);
   Y1_c41 <= Y1_copy187_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid189
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid189 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid189 is
   component MultTable_Freq800_uid191 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy192_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid191
      port map ( X => Xtable_c41,
                 Y => Y1_copy192_c41);
   Y1_c41 <= Y1_copy192_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid194
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid194 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid194 is
   component MultTable_Freq800_uid196 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy197_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid196
      port map ( X => Xtable_c41,
                 Y => Y1_copy197_c41);
   Y1_c41 <= Y1_copy197_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid199
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid199 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid199 is
   component MultTable_Freq800_uid201 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy202_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid201
      port map ( X => Xtable_c41,
                 Y => Y1_copy202_c41);
   Y1_c41 <= Y1_copy202_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid204
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid204 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid204 is
   component MultTable_Freq800_uid206 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(3 downto 0);
signal Y1_c41 :  std_logic_vector(3 downto 0);
signal Y1_copy207_c41 :  std_logic_vector(3 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid206
      port map ( X => Xtable_c41,
                 Y => Y1_copy207_c41);
   Y1_c41 <= Y1_copy207_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid209
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid209 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid209 is
   component MultTable_Freq800_uid211 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy212_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid211
      port map ( X => Xtable_c41,
                 Y => Y1_copy212_c41);
   Y1_c41 <= Y1_copy212_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid214
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid214 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid214 is
   component MultTable_Freq800_uid216 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy217_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid216
      port map ( X => Xtable_c41,
                 Y => Y1_copy217_c41);
   Y1_c41 <= Y1_copy217_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid219
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid219 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid219 is
   component MultTable_Freq800_uid221 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy222_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid221
      port map ( X => Xtable_c41,
                 Y => Y1_copy222_c41);
   Y1_c41 <= Y1_copy222_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid224
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid224 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid224 is
   component MultTable_Freq800_uid226 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy227_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid226
      port map ( X => Xtable_c41,
                 Y => Y1_copy227_c41);
   Y1_c41 <= Y1_copy227_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid229
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid229 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid229 is
   component MultTable_Freq800_uid231 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy232_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid231
      port map ( X => Xtable_c41,
                 Y => Y1_copy232_c41);
   Y1_c41 <= Y1_copy232_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid234
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid234 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid234 is
   component MultTable_Freq800_uid236 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(3 downto 0);
signal Y1_c41 :  std_logic_vector(3 downto 0);
signal Y1_copy237_c41 :  std_logic_vector(3 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid236
      port map ( X => Xtable_c41,
                 Y => Y1_copy237_c41);
   Y1_c41 <= Y1_copy237_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid239
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid239 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid239 is
   component MultTable_Freq800_uid241 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy242_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid241
      port map ( X => Xtable_c41,
                 Y => Y1_copy242_c41);
   Y1_c41 <= Y1_copy242_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid244
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid244 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid244 is
   component MultTable_Freq800_uid246 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy247_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid246
      port map ( X => Xtable_c41,
                 Y => Y1_copy247_c41);
   Y1_c41 <= Y1_copy247_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid249
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid249 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid249 is
   component MultTable_Freq800_uid251 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy252_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid251
      port map ( X => Xtable_c41,
                 Y => Y1_copy252_c41);
   Y1_c41 <= Y1_copy252_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid254
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid254 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid254 is
   component MultTable_Freq800_uid256 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy257_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid256
      port map ( X => Xtable_c41,
                 Y => Y1_copy257_c41);
   Y1_c41 <= Y1_copy257_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid259
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid259 is
    port (clk, ce_39, ce_40, ce_41 : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid259 is
   component MultTable_Freq800_uid261 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c41 :  std_logic_vector(4 downto 0);
signal Y1_c41 :  std_logic_vector(4 downto 0);
signal Y1_copy262_c41 :  std_logic_vector(4 downto 0);
signal Y_c39, Y_c40, Y_c41 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               Y_c39 <= Y;
            end if;
            if ce_40 = '1' then
               Y_c40 <= Y_c39;
            end if;
            if ce_41 = '1' then
               Y_c41 <= Y_c40;
            end if;
         end if;
      end process;
Xtable_c41 <= Y_c41 & X;
   R <= Y1_c41;
   TableMult: MultTable_Freq800_uid261
      port map ( X => Xtable_c41,
                 Y => Y1_copy262_c41);
   Y1_c41 <= Y1_copy262_c41; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_19_Freq800_uid441
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 50 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_19_Freq800_uid441 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50 : in std_logic;
          X : in  std_logic_vector(18 downto 0);
          Y : in  std_logic_vector(18 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(18 downto 0)   );
end entity;

architecture arch of IntAdder_19_Freq800_uid441 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3, Cin_0_c4, Cin_0_c5, Cin_0_c6, Cin_0_c7, Cin_0_c8, Cin_0_c9, Cin_0_c10, Cin_0_c11, Cin_0_c12, Cin_0_c13, Cin_0_c14, Cin_0_c15, Cin_0_c16, Cin_0_c17, Cin_0_c18, Cin_0_c19, Cin_0_c20, Cin_0_c21, Cin_0_c22, Cin_0_c23, Cin_0_c24, Cin_0_c25, Cin_0_c26, Cin_0_c27, Cin_0_c28, Cin_0_c29, Cin_0_c30, Cin_0_c31, Cin_0_c32, Cin_0_c33, Cin_0_c34, Cin_0_c35, Cin_0_c36, Cin_0_c37, Cin_0_c38, Cin_0_c39, Cin_0_c40, Cin_0_c41, Cin_0_c42, Cin_0_c43, Cin_0_c44 :  std_logic;
signal X_0_c43, X_0_c44 :  std_logic_vector(3 downto 0);
signal Y_0_c43, Y_0_c44 :  std_logic_vector(3 downto 0);
signal S_0_c44 :  std_logic_vector(3 downto 0);
signal R_0_c44, R_0_c45, R_0_c46, R_0_c47, R_0_c48, R_0_c49, R_0_c50 :  std_logic_vector(2 downto 0);
signal Cin_1_c44, Cin_1_c45 :  std_logic;
signal X_1_c43, X_1_c44, X_1_c45 :  std_logic_vector(3 downto 0);
signal Y_1_c43, Y_1_c44, Y_1_c45 :  std_logic_vector(3 downto 0);
signal S_1_c45 :  std_logic_vector(3 downto 0);
signal R_1_c45, R_1_c46, R_1_c47, R_1_c48, R_1_c49, R_1_c50 :  std_logic_vector(2 downto 0);
signal Cin_2_c45, Cin_2_c46 :  std_logic;
signal X_2_c43, X_2_c44, X_2_c45, X_2_c46 :  std_logic_vector(3 downto 0);
signal Y_2_c43, Y_2_c44, Y_2_c45, Y_2_c46 :  std_logic_vector(3 downto 0);
signal S_2_c46 :  std_logic_vector(3 downto 0);
signal R_2_c46, R_2_c47, R_2_c48, R_2_c49, R_2_c50 :  std_logic_vector(2 downto 0);
signal Cin_3_c46, Cin_3_c47 :  std_logic;
signal X_3_c43, X_3_c44, X_3_c45, X_3_c46, X_3_c47 :  std_logic_vector(3 downto 0);
signal Y_3_c43, Y_3_c44, Y_3_c45, Y_3_c46, Y_3_c47 :  std_logic_vector(3 downto 0);
signal S_3_c47 :  std_logic_vector(3 downto 0);
signal R_3_c47, R_3_c48, R_3_c49, R_3_c50 :  std_logic_vector(2 downto 0);
signal Cin_4_c47, Cin_4_c48 :  std_logic;
signal X_4_c43, X_4_c44, X_4_c45, X_4_c46, X_4_c47, X_4_c48 :  std_logic_vector(3 downto 0);
signal Y_4_c43, Y_4_c44, Y_4_c45, Y_4_c46, Y_4_c47, Y_4_c48 :  std_logic_vector(3 downto 0);
signal S_4_c48 :  std_logic_vector(3 downto 0);
signal R_4_c48, R_4_c49, R_4_c50 :  std_logic_vector(2 downto 0);
signal Cin_5_c48, Cin_5_c49, Cin_5_c50 :  std_logic;
signal X_5_c43, X_5_c44, X_5_c45, X_5_c46, X_5_c47, X_5_c48, X_5_c49, X_5_c50 :  std_logic_vector(3 downto 0);
signal Y_5_c43, Y_5_c44, Y_5_c45, Y_5_c46, Y_5_c47, Y_5_c48, Y_5_c49, Y_5_c50 :  std_logic_vector(3 downto 0);
signal S_5_c50 :  std_logic_vector(3 downto 0);
signal R_5_c50 :  std_logic_vector(2 downto 0);
signal Cin_6_c50 :  std_logic;
signal X_6_c43, X_6_c44, X_6_c45, X_6_c46, X_6_c47, X_6_c48, X_6_c49, X_6_c50 :  std_logic_vector(1 downto 0);
signal Y_6_c43, Y_6_c44, Y_6_c45, Y_6_c46, Y_6_c47, Y_6_c48, Y_6_c49, Y_6_c50 :  std_logic_vector(1 downto 0);
signal S_6_c50 :  std_logic_vector(1 downto 0);
signal R_6_c50 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
            end if;
            if ce_4 = '1' then
               Cin_0_c4 <= Cin_0_c3;
            end if;
            if ce_5 = '1' then
               Cin_0_c5 <= Cin_0_c4;
            end if;
            if ce_6 = '1' then
               Cin_0_c6 <= Cin_0_c5;
            end if;
            if ce_7 = '1' then
               Cin_0_c7 <= Cin_0_c6;
            end if;
            if ce_8 = '1' then
               Cin_0_c8 <= Cin_0_c7;
            end if;
            if ce_9 = '1' then
               Cin_0_c9 <= Cin_0_c8;
            end if;
            if ce_10 = '1' then
               Cin_0_c10 <= Cin_0_c9;
            end if;
            if ce_11 = '1' then
               Cin_0_c11 <= Cin_0_c10;
            end if;
            if ce_12 = '1' then
               Cin_0_c12 <= Cin_0_c11;
            end if;
            if ce_13 = '1' then
               Cin_0_c13 <= Cin_0_c12;
            end if;
            if ce_14 = '1' then
               Cin_0_c14 <= Cin_0_c13;
            end if;
            if ce_15 = '1' then
               Cin_0_c15 <= Cin_0_c14;
            end if;
            if ce_16 = '1' then
               Cin_0_c16 <= Cin_0_c15;
            end if;
            if ce_17 = '1' then
               Cin_0_c17 <= Cin_0_c16;
            end if;
            if ce_18 = '1' then
               Cin_0_c18 <= Cin_0_c17;
            end if;
            if ce_19 = '1' then
               Cin_0_c19 <= Cin_0_c18;
            end if;
            if ce_20 = '1' then
               Cin_0_c20 <= Cin_0_c19;
            end if;
            if ce_21 = '1' then
               Cin_0_c21 <= Cin_0_c20;
            end if;
            if ce_22 = '1' then
               Cin_0_c22 <= Cin_0_c21;
            end if;
            if ce_23 = '1' then
               Cin_0_c23 <= Cin_0_c22;
            end if;
            if ce_24 = '1' then
               Cin_0_c24 <= Cin_0_c23;
            end if;
            if ce_25 = '1' then
               Cin_0_c25 <= Cin_0_c24;
            end if;
            if ce_26 = '1' then
               Cin_0_c26 <= Cin_0_c25;
            end if;
            if ce_27 = '1' then
               Cin_0_c27 <= Cin_0_c26;
            end if;
            if ce_28 = '1' then
               Cin_0_c28 <= Cin_0_c27;
            end if;
            if ce_29 = '1' then
               Cin_0_c29 <= Cin_0_c28;
            end if;
            if ce_30 = '1' then
               Cin_0_c30 <= Cin_0_c29;
            end if;
            if ce_31 = '1' then
               Cin_0_c31 <= Cin_0_c30;
            end if;
            if ce_32 = '1' then
               Cin_0_c32 <= Cin_0_c31;
            end if;
            if ce_33 = '1' then
               Cin_0_c33 <= Cin_0_c32;
            end if;
            if ce_34 = '1' then
               Cin_0_c34 <= Cin_0_c33;
            end if;
            if ce_35 = '1' then
               Cin_0_c35 <= Cin_0_c34;
            end if;
            if ce_36 = '1' then
               Cin_0_c36 <= Cin_0_c35;
            end if;
            if ce_37 = '1' then
               Cin_0_c37 <= Cin_0_c36;
            end if;
            if ce_38 = '1' then
               Cin_0_c38 <= Cin_0_c37;
            end if;
            if ce_39 = '1' then
               Cin_0_c39 <= Cin_0_c38;
            end if;
            if ce_40 = '1' then
               Cin_0_c40 <= Cin_0_c39;
            end if;
            if ce_41 = '1' then
               Cin_0_c41 <= Cin_0_c40;
            end if;
            if ce_42 = '1' then
               Cin_0_c42 <= Cin_0_c41;
            end if;
            if ce_43 = '1' then
               Cin_0_c43 <= Cin_0_c42;
            end if;
            if ce_44 = '1' then
               Cin_0_c44 <= Cin_0_c43;
               X_0_c44 <= X_0_c43;
               Y_0_c44 <= Y_0_c43;
               X_1_c44 <= X_1_c43;
               Y_1_c44 <= Y_1_c43;
               X_2_c44 <= X_2_c43;
               Y_2_c44 <= Y_2_c43;
               X_3_c44 <= X_3_c43;
               Y_3_c44 <= Y_3_c43;
               X_4_c44 <= X_4_c43;
               Y_4_c44 <= Y_4_c43;
               X_5_c44 <= X_5_c43;
               Y_5_c44 <= Y_5_c43;
               X_6_c44 <= X_6_c43;
               Y_6_c44 <= Y_6_c43;
            end if;
            if ce_45 = '1' then
               R_0_c45 <= R_0_c44;
               Cin_1_c45 <= Cin_1_c44;
               X_1_c45 <= X_1_c44;
               Y_1_c45 <= Y_1_c44;
               X_2_c45 <= X_2_c44;
               Y_2_c45 <= Y_2_c44;
               X_3_c45 <= X_3_c44;
               Y_3_c45 <= Y_3_c44;
               X_4_c45 <= X_4_c44;
               Y_4_c45 <= Y_4_c44;
               X_5_c45 <= X_5_c44;
               Y_5_c45 <= Y_5_c44;
               X_6_c45 <= X_6_c44;
               Y_6_c45 <= Y_6_c44;
            end if;
            if ce_46 = '1' then
               R_0_c46 <= R_0_c45;
               R_1_c46 <= R_1_c45;
               Cin_2_c46 <= Cin_2_c45;
               X_2_c46 <= X_2_c45;
               Y_2_c46 <= Y_2_c45;
               X_3_c46 <= X_3_c45;
               Y_3_c46 <= Y_3_c45;
               X_4_c46 <= X_4_c45;
               Y_4_c46 <= Y_4_c45;
               X_5_c46 <= X_5_c45;
               Y_5_c46 <= Y_5_c45;
               X_6_c46 <= X_6_c45;
               Y_6_c46 <= Y_6_c45;
            end if;
            if ce_47 = '1' then
               R_0_c47 <= R_0_c46;
               R_1_c47 <= R_1_c46;
               R_2_c47 <= R_2_c46;
               Cin_3_c47 <= Cin_3_c46;
               X_3_c47 <= X_3_c46;
               Y_3_c47 <= Y_3_c46;
               X_4_c47 <= X_4_c46;
               Y_4_c47 <= Y_4_c46;
               X_5_c47 <= X_5_c46;
               Y_5_c47 <= Y_5_c46;
               X_6_c47 <= X_6_c46;
               Y_6_c47 <= Y_6_c46;
            end if;
            if ce_48 = '1' then
               R_0_c48 <= R_0_c47;
               R_1_c48 <= R_1_c47;
               R_2_c48 <= R_2_c47;
               R_3_c48 <= R_3_c47;
               Cin_4_c48 <= Cin_4_c47;
               X_4_c48 <= X_4_c47;
               Y_4_c48 <= Y_4_c47;
               X_5_c48 <= X_5_c47;
               Y_5_c48 <= Y_5_c47;
               X_6_c48 <= X_6_c47;
               Y_6_c48 <= Y_6_c47;
            end if;
            if ce_49 = '1' then
               R_0_c49 <= R_0_c48;
               R_1_c49 <= R_1_c48;
               R_2_c49 <= R_2_c48;
               R_3_c49 <= R_3_c48;
               R_4_c49 <= R_4_c48;
               Cin_5_c49 <= Cin_5_c48;
               X_5_c49 <= X_5_c48;
               Y_5_c49 <= Y_5_c48;
               X_6_c49 <= X_6_c48;
               Y_6_c49 <= Y_6_c48;
            end if;
            if ce_50 = '1' then
               R_0_c50 <= R_0_c49;
               R_1_c50 <= R_1_c49;
               R_2_c50 <= R_2_c49;
               R_3_c50 <= R_3_c49;
               R_4_c50 <= R_4_c49;
               Cin_5_c50 <= Cin_5_c49;
               X_5_c50 <= X_5_c49;
               Y_5_c50 <= Y_5_c49;
               X_6_c50 <= X_6_c49;
               Y_6_c50 <= Y_6_c49;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c43 <= '0' & X(2 downto 0);
   Y_0_c43 <= '0' & Y(2 downto 0);
   S_0_c44 <= X_0_c44 + Y_0_c44 + Cin_0_c44;
   R_0_c44 <= S_0_c44(2 downto 0);
   Cin_1_c44 <= S_0_c44(3);
   X_1_c43 <= '0' & X(5 downto 3);
   Y_1_c43 <= '0' & Y(5 downto 3);
   S_1_c45 <= X_1_c45 + Y_1_c45 + Cin_1_c45;
   R_1_c45 <= S_1_c45(2 downto 0);
   Cin_2_c45 <= S_1_c45(3);
   X_2_c43 <= '0' & X(8 downto 6);
   Y_2_c43 <= '0' & Y(8 downto 6);
   S_2_c46 <= X_2_c46 + Y_2_c46 + Cin_2_c46;
   R_2_c46 <= S_2_c46(2 downto 0);
   Cin_3_c46 <= S_2_c46(3);
   X_3_c43 <= '0' & X(11 downto 9);
   Y_3_c43 <= '0' & Y(11 downto 9);
   S_3_c47 <= X_3_c47 + Y_3_c47 + Cin_3_c47;
   R_3_c47 <= S_3_c47(2 downto 0);
   Cin_4_c47 <= S_3_c47(3);
   X_4_c43 <= '0' & X(14 downto 12);
   Y_4_c43 <= '0' & Y(14 downto 12);
   S_4_c48 <= X_4_c48 + Y_4_c48 + Cin_4_c48;
   R_4_c48 <= S_4_c48(2 downto 0);
   Cin_5_c48 <= S_4_c48(3);
   X_5_c43 <= '0' & X(17 downto 15);
   Y_5_c43 <= '0' & Y(17 downto 15);
   S_5_c50 <= X_5_c50 + Y_5_c50 + Cin_5_c50;
   R_5_c50 <= S_5_c50(2 downto 0);
   Cin_6_c50 <= S_5_c50(3);
   X_6_c43 <= '0' & X(18 downto 18);
   Y_6_c43 <= '0' & Y(18 downto 18);
   S_6_c50 <= X_6_c50 + Y_6_c50 + Cin_6_c50;
   R_6_c50 <= S_6_c50(0 downto 0);
   R <= R_6_c50 & R_5_c50 & R_4_c50 & R_3_c50 & R_2_c50 & R_1_c50 & R_0_c50 ;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_17x18_19_Freq800_uid54
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_17x18_19_Freq800_uid54 is
    port (clk, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(17 downto 0);
          R : out  std_logic_vector(18 downto 0)   );
end entity;

architecture arch of IntMultiplier_17x18_19_Freq800_uid54 is
   component IntMultiplierLUT_1x1_Freq800_uid58 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid60 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid65 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid70 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq800_uid72 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid74 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid79 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid84 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid86 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid91 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid96 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid101 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid103 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid108 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid113 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid118 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid123 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_2x1_Freq800_uid125 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid127 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid132 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid137 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid142 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid147 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid149 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid154 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid159 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid164 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid169 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid174 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid179 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid184 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid189 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid194 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid199 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid204 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid209 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid214 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid219 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid224 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid229 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid234 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid239 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid244 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid249 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid254 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid259 is
      port ( clk, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_6_3_Freq800_uid265 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq800_uid271 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq800_uid277 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_23_3_Freq800_uid289 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_19_Freq800_uid441 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50 : in std_logic;
             X : in  std_logic_vector(18 downto 0);
             Y : in  std_logic_vector(18 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(18 downto 0)   );
   end component;

signal XX_m55_c41 :  std_logic_vector(16 downto 0);
signal YY_m55_c38 :  std_logic_vector(17 downto 0);
signal tile_0_X_c41 :  std_logic_vector(0 downto 0);
signal tile_0_Y_c38 :  std_logic_vector(0 downto 0);
signal tile_0_output_c41 :  std_logic_vector(0 downto 0);
signal tile_0_filtered_output_c41 :  unsigned(0-0 downto 0);
signal bh56_w12_0_c41 :  std_logic;
signal tile_1_X_c41 :  std_logic_vector(1 downto 0);
signal tile_1_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_1_output_c41 :  std_logic_vector(3 downto 0);
signal tile_1_filtered_output_c41 :  unsigned(3-0 downto 0);
signal bh56_w12_1_c41 :  std_logic;
signal bh56_w13_0_c41 :  std_logic;
signal bh56_w14_0_c41 :  std_logic;
signal bh56_w15_0_c41 :  std_logic;
signal tile_2_X_c41 :  std_logic_vector(2 downto 0);
signal tile_2_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_2_output_c41 :  std_logic_vector(4 downto 0);
signal tile_2_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w14_1_c41 :  std_logic;
signal bh56_w15_1_c41 :  std_logic;
signal bh56_w16_0_c41 :  std_logic;
signal bh56_w17_0_c41 :  std_logic;
signal bh56_w18_0_c41 :  std_logic;
signal tile_3_X_c41 :  std_logic_vector(0 downto 0);
signal tile_3_Y_c38 :  std_logic_vector(0 downto 0);
signal tile_3_output_c41 :  std_logic_vector(0 downto 0);
signal tile_3_filtered_output_c41 :  unsigned(0-0 downto 0);
signal bh56_w12_2_c41 :  std_logic;
signal tile_4_X_c41 :  std_logic_vector(1 downto 0);
signal tile_4_Y_c38 :  std_logic_vector(0 downto 0);
signal tile_4_output_c41 :  std_logic_vector(1 downto 0);
signal tile_4_filtered_output_c41 :  unsigned(1-0 downto 0);
signal bh56_w12_3_c41 :  std_logic;
signal bh56_w13_1_c41 :  std_logic;
signal tile_5_X_c41 :  std_logic_vector(2 downto 0);
signal tile_5_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_5_output_c41 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w13_2_c41 :  std_logic;
signal bh56_w14_2_c41 :  std_logic;
signal bh56_w15_2_c41 :  std_logic;
signal bh56_w16_1_c41 :  std_logic;
signal bh56_w17_1_c41 :  std_logic;
signal tile_6_X_c41 :  std_logic_vector(2 downto 0);
signal tile_6_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_6_output_c41 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w16_2_c41 :  std_logic;
signal bh56_w17_2_c41 :  std_logic;
signal bh56_w18_1_c41 :  std_logic;
signal bh56_w19_0_c41 :  std_logic;
signal bh56_w20_0_c41 :  std_logic;
signal tile_7_X_c41 :  std_logic_vector(0 downto 0);
signal tile_7_Y_c38 :  std_logic_vector(0 downto 0);
signal tile_7_output_c41 :  std_logic_vector(0 downto 0);
signal tile_7_filtered_output_c41 :  unsigned(0-0 downto 0);
signal bh56_w12_4_c41 :  std_logic;
signal tile_8_X_c41 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_8_output_c41 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w12_5_c41 :  std_logic;
signal bh56_w13_3_c41 :  std_logic;
signal bh56_w14_3_c41 :  std_logic;
signal bh56_w15_3_c41 :  std_logic;
signal bh56_w16_3_c41 :  std_logic;
signal tile_9_X_c41 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_9_output_c41 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w15_4_c41 :  std_logic;
signal bh56_w16_4_c41 :  std_logic;
signal bh56_w17_3_c41 :  std_logic;
signal bh56_w18_2_c41 :  std_logic;
signal bh56_w19_1_c41 :  std_logic;
signal tile_10_X_c41 :  std_logic_vector(2 downto 0);
signal tile_10_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_10_output_c41 :  std_logic_vector(4 downto 0);
signal tile_10_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w18_3_c41 :  std_logic;
signal bh56_w19_2_c41 :  std_logic;
signal bh56_w20_1_c41 :  std_logic;
signal bh56_w21_0_c41 :  std_logic;
signal bh56_w22_0_c41 :  std_logic;
signal tile_11_X_c41 :  std_logic_vector(0 downto 0);
signal tile_11_Y_c38 :  std_logic_vector(0 downto 0);
signal tile_11_output_c41 :  std_logic_vector(0 downto 0);
signal tile_11_filtered_output_c41 :  unsigned(0-0 downto 0);
signal bh56_w12_6_c41 :  std_logic;
signal tile_12_X_c41 :  std_logic_vector(1 downto 0);
signal tile_12_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_12_output_c41 :  std_logic_vector(3 downto 0);
signal tile_12_filtered_output_c41 :  unsigned(3-0 downto 0);
signal bh56_w12_7_c41 :  std_logic;
signal bh56_w13_4_c41 :  std_logic;
signal bh56_w14_4_c41 :  std_logic;
signal bh56_w15_5_c41 :  std_logic;
signal tile_13_X_c41 :  std_logic_vector(2 downto 0);
signal tile_13_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_13_output_c41 :  std_logic_vector(4 downto 0);
signal tile_13_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w14_5_c41 :  std_logic;
signal bh56_w15_6_c41 :  std_logic;
signal bh56_w16_5_c41 :  std_logic;
signal bh56_w17_4_c41 :  std_logic;
signal bh56_w18_4_c41 :  std_logic;
signal tile_14_X_c41 :  std_logic_vector(2 downto 0);
signal tile_14_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_14_output_c41 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w17_5_c41 :  std_logic;
signal bh56_w18_5_c41 :  std_logic;
signal bh56_w19_3_c41 :  std_logic;
signal bh56_w20_2_c41 :  std_logic;
signal bh56_w21_1_c41 :  std_logic;
signal tile_15_X_c41 :  std_logic_vector(2 downto 0);
signal tile_15_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_15_output_c41 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w20_3_c41 :  std_logic;
signal bh56_w21_2_c41 :  std_logic;
signal bh56_w22_1_c41 :  std_logic;
signal bh56_w23_0_c41 :  std_logic;
signal bh56_w24_0_c41 :  std_logic;
signal tile_16_X_c41 :  std_logic_vector(0 downto 0);
signal tile_16_Y_c38 :  std_logic_vector(0 downto 0);
signal tile_16_output_c41 :  std_logic_vector(0 downto 0);
signal tile_16_filtered_output_c41 :  unsigned(0-0 downto 0);
signal bh56_w12_8_c41 :  std_logic;
signal tile_17_X_c41 :  std_logic_vector(1 downto 0);
signal tile_17_Y_c38 :  std_logic_vector(0 downto 0);
signal tile_17_output_c41 :  std_logic_vector(1 downto 0);
signal tile_17_filtered_output_c41 :  unsigned(1-0 downto 0);
signal bh56_w12_9_c41 :  std_logic;
signal bh56_w13_5_c41 :  std_logic;
signal tile_18_X_c41 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_18_output_c41 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w13_6_c41 :  std_logic;
signal bh56_w14_6_c41 :  std_logic;
signal bh56_w15_7_c41 :  std_logic;
signal bh56_w16_6_c41 :  std_logic;
signal bh56_w17_6_c41 :  std_logic;
signal tile_19_X_c41 :  std_logic_vector(2 downto 0);
signal tile_19_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_19_output_c41 :  std_logic_vector(4 downto 0);
signal tile_19_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w16_7_c41 :  std_logic;
signal bh56_w17_7_c41 :  std_logic;
signal bh56_w18_6_c41 :  std_logic;
signal bh56_w19_4_c41 :  std_logic;
signal bh56_w20_4_c41 :  std_logic;
signal tile_20_X_c41 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_20_output_c41 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w19_5_c41 :  std_logic;
signal bh56_w20_5_c41 :  std_logic;
signal bh56_w21_3_c41 :  std_logic;
signal bh56_w22_2_c41 :  std_logic;
signal bh56_w23_1_c41 :  std_logic;
signal tile_21_X_c41 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_21_output_c41 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w22_3_c41 :  std_logic;
signal bh56_w23_2_c41 :  std_logic;
signal bh56_w24_1_c41 :  std_logic;
signal bh56_w25_0_c41 :  std_logic;
signal bh56_w26_0_c41 :  std_logic;
signal tile_22_X_c41 :  std_logic_vector(0 downto 0);
signal tile_22_Y_c38 :  std_logic_vector(0 downto 0);
signal tile_22_output_c41 :  std_logic_vector(0 downto 0);
signal tile_22_filtered_output_c41 :  unsigned(0-0 downto 0);
signal bh56_w12_10_c41 :  std_logic;
signal tile_23_X_c41 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_23_output_c41 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w12_11_c41 :  std_logic;
signal bh56_w13_7_c41 :  std_logic;
signal bh56_w14_7_c41 :  std_logic;
signal bh56_w15_8_c41 :  std_logic;
signal bh56_w16_8_c41 :  std_logic;
signal tile_24_X_c41 :  std_logic_vector(2 downto 0);
signal tile_24_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_24_output_c41 :  std_logic_vector(4 downto 0);
signal tile_24_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w15_9_c41 :  std_logic;
signal bh56_w16_9_c41 :  std_logic;
signal bh56_w17_8_c41 :  std_logic;
signal bh56_w18_7_c41 :  std_logic;
signal bh56_w19_6_c41, bh56_w19_6_c42 :  std_logic;
signal tile_25_X_c41 :  std_logic_vector(2 downto 0);
signal tile_25_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_25_output_c41 :  std_logic_vector(4 downto 0);
signal tile_25_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w18_8_c41 :  std_logic;
signal bh56_w19_7_c41 :  std_logic;
signal bh56_w20_6_c41 :  std_logic;
signal bh56_w21_4_c41 :  std_logic;
signal bh56_w22_4_c41 :  std_logic;
signal tile_26_X_c41 :  std_logic_vector(2 downto 0);
signal tile_26_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_26_output_c41 :  std_logic_vector(4 downto 0);
signal tile_26_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w21_5_c41 :  std_logic;
signal bh56_w22_5_c41 :  std_logic;
signal bh56_w23_3_c41 :  std_logic;
signal bh56_w24_2_c41 :  std_logic;
signal bh56_w25_1_c41 :  std_logic;
signal tile_27_X_c41 :  std_logic_vector(2 downto 0);
signal tile_27_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_27_output_c41 :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w24_3_c41 :  std_logic;
signal bh56_w25_2_c41 :  std_logic;
signal bh56_w26_1_c41 :  std_logic;
signal bh56_w27_0_c41 :  std_logic;
signal bh56_w28_0_c41 :  std_logic;
signal tile_28_X_c41 :  std_logic_vector(1 downto 0);
signal tile_28_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_28_output_c41 :  std_logic_vector(3 downto 0);
signal tile_28_filtered_output_c41 :  unsigned(3-0 downto 0);
signal bh56_w12_12_c41 :  std_logic;
signal bh56_w13_8_c41 :  std_logic;
signal bh56_w14_8_c41 :  std_logic;
signal bh56_w15_10_c41 :  std_logic;
signal tile_29_X_c41 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_29_output_c41 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w14_9_c41 :  std_logic;
signal bh56_w15_11_c41 :  std_logic;
signal bh56_w16_10_c41 :  std_logic;
signal bh56_w17_9_c41 :  std_logic;
signal bh56_w18_9_c41 :  std_logic;
signal tile_30_X_c41 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_30_output_c41 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w17_10_c41 :  std_logic;
signal bh56_w18_10_c41 :  std_logic;
signal bh56_w19_8_c41 :  std_logic;
signal bh56_w20_7_c41 :  std_logic;
signal bh56_w21_6_c41 :  std_logic;
signal tile_31_X_c41 :  std_logic_vector(2 downto 0);
signal tile_31_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_31_output_c41 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w20_8_c41 :  std_logic;
signal bh56_w21_7_c41 :  std_logic;
signal bh56_w22_6_c41 :  std_logic;
signal bh56_w23_4_c41 :  std_logic;
signal bh56_w24_4_c41 :  std_logic;
signal tile_32_X_c41 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_32_output_c41 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w23_5_c41 :  std_logic;
signal bh56_w24_5_c41 :  std_logic;
signal bh56_w25_3_c41 :  std_logic;
signal bh56_w26_2_c41 :  std_logic;
signal bh56_w27_1_c41 :  std_logic;
signal tile_33_X_c41 :  std_logic_vector(2 downto 0);
signal tile_33_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_33_output_c41 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w26_3_c41 :  std_logic;
signal bh56_w27_2_c41 :  std_logic;
signal bh56_w28_1_c41 :  std_logic;
signal bh56_w29_0_c41 :  std_logic;
signal bh56_w30_0_c41 :  std_logic;
signal tile_34_X_c41 :  std_logic_vector(1 downto 0);
signal tile_34_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_34_output_c41 :  std_logic_vector(3 downto 0);
signal tile_34_filtered_output_c41 :  unsigned(3-0 downto 0);
signal bh56_w14_10_c41 :  std_logic;
signal bh56_w15_12_c41 :  std_logic;
signal bh56_w16_11_c41 :  std_logic;
signal bh56_w17_11_c41 :  std_logic;
signal tile_35_X_c41 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_35_output_c41 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w16_12_c41 :  std_logic;
signal bh56_w17_12_c41 :  std_logic;
signal bh56_w18_11_c41 :  std_logic;
signal bh56_w19_9_c41 :  std_logic;
signal bh56_w20_9_c41 :  std_logic;
signal tile_36_X_c41 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_36_output_c41 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w19_10_c41 :  std_logic;
signal bh56_w20_10_c41 :  std_logic;
signal bh56_w21_8_c41 :  std_logic;
signal bh56_w22_7_c41 :  std_logic;
signal bh56_w23_6_c41 :  std_logic;
signal tile_37_X_c41 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_37_output_c41 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w22_8_c41 :  std_logic;
signal bh56_w23_7_c41 :  std_logic;
signal bh56_w24_6_c41 :  std_logic;
signal bh56_w25_4_c41 :  std_logic;
signal bh56_w26_4_c41 :  std_logic;
signal tile_38_X_c41 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_38_output_c41 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w25_5_c41 :  std_logic;
signal bh56_w26_5_c41 :  std_logic;
signal bh56_w27_3_c41 :  std_logic;
signal bh56_w28_2_c41 :  std_logic;
signal bh56_w29_1_c41 :  std_logic;
signal tile_39_X_c41 :  std_logic_vector(2 downto 0);
signal tile_39_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_39_output_c41 :  std_logic_vector(4 downto 0);
signal tile_39_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w28_3_c41 :  std_logic;
signal bh56_w29_2_c41 :  std_logic;
signal bh56_w30_1_c41 :  std_logic;
signal bh56_w31_0_c41 :  std_logic;
signal bh56_w32_0_c41 :  std_logic;
signal tile_40_X_c41 :  std_logic_vector(1 downto 0);
signal tile_40_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_40_output_c41 :  std_logic_vector(3 downto 0);
signal tile_40_filtered_output_c41 :  unsigned(3-0 downto 0);
signal bh56_w16_13_c41 :  std_logic;
signal bh56_w17_13_c41 :  std_logic;
signal bh56_w18_12_c41 :  std_logic;
signal bh56_w19_11_c41 :  std_logic;
signal tile_41_X_c41 :  std_logic_vector(2 downto 0);
signal tile_41_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_41_output_c41 :  std_logic_vector(4 downto 0);
signal tile_41_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w18_13_c41 :  std_logic;
signal bh56_w19_12_c41 :  std_logic;
signal bh56_w20_11_c41 :  std_logic;
signal bh56_w21_9_c41 :  std_logic;
signal bh56_w22_9_c41 :  std_logic;
signal tile_42_X_c41 :  std_logic_vector(2 downto 0);
signal tile_42_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_42_output_c41 :  std_logic_vector(4 downto 0);
signal tile_42_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w21_10_c41, bh56_w21_10_c42 :  std_logic;
signal bh56_w22_10_c41 :  std_logic;
signal bh56_w23_8_c41 :  std_logic;
signal bh56_w24_7_c41 :  std_logic;
signal bh56_w25_6_c41 :  std_logic;
signal tile_43_X_c41 :  std_logic_vector(2 downto 0);
signal tile_43_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_43_output_c41 :  std_logic_vector(4 downto 0);
signal tile_43_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w24_8_c41 :  std_logic;
signal bh56_w25_7_c41 :  std_logic;
signal bh56_w26_6_c41 :  std_logic;
signal bh56_w27_4_c41 :  std_logic;
signal bh56_w28_4_c41 :  std_logic;
signal tile_44_X_c41 :  std_logic_vector(2 downto 0);
signal tile_44_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_44_output_c41 :  std_logic_vector(4 downto 0);
signal tile_44_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w27_5_c41 :  std_logic;
signal bh56_w28_5_c41 :  std_logic;
signal bh56_w29_3_c41 :  std_logic;
signal bh56_w30_2_c41 :  std_logic;
signal bh56_w31_1_c41 :  std_logic;
signal tile_45_X_c41 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c38 :  std_logic_vector(1 downto 0);
signal tile_45_output_c41 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c41 :  unsigned(4-0 downto 0);
signal bh56_w30_3_c41 :  std_logic;
signal bh56_w31_2_c41, bh56_w31_2_c42 :  std_logic;
signal bh56_w32_1_c41 :  std_logic;
signal bh56_w33_0_c41 :  std_logic;
signal bh56_w34_0_c41, bh56_w34_0_c42 :  std_logic;
signal bh56_w12_13_c0, bh56_w12_13_c1, bh56_w12_13_c2, bh56_w12_13_c3, bh56_w12_13_c4, bh56_w12_13_c5, bh56_w12_13_c6, bh56_w12_13_c7, bh56_w12_13_c8, bh56_w12_13_c9, bh56_w12_13_c10, bh56_w12_13_c11, bh56_w12_13_c12, bh56_w12_13_c13, bh56_w12_13_c14, bh56_w12_13_c15, bh56_w12_13_c16, bh56_w12_13_c17, bh56_w12_13_c18, bh56_w12_13_c19, bh56_w12_13_c20, bh56_w12_13_c21, bh56_w12_13_c22, bh56_w12_13_c23, bh56_w12_13_c24, bh56_w12_13_c25, bh56_w12_13_c26, bh56_w12_13_c27, bh56_w12_13_c28, bh56_w12_13_c29, bh56_w12_13_c30, bh56_w12_13_c31, bh56_w12_13_c32, bh56_w12_13_c33, bh56_w12_13_c34, bh56_w12_13_c35, bh56_w12_13_c36, bh56_w12_13_c37, bh56_w12_13_c38, bh56_w12_13_c39, bh56_w12_13_c40, bh56_w12_13_c41 :  std_logic;
signal bh56_w13_9_c0, bh56_w13_9_c1, bh56_w13_9_c2, bh56_w13_9_c3, bh56_w13_9_c4, bh56_w13_9_c5, bh56_w13_9_c6, bh56_w13_9_c7, bh56_w13_9_c8, bh56_w13_9_c9, bh56_w13_9_c10, bh56_w13_9_c11, bh56_w13_9_c12, bh56_w13_9_c13, bh56_w13_9_c14, bh56_w13_9_c15, bh56_w13_9_c16, bh56_w13_9_c17, bh56_w13_9_c18, bh56_w13_9_c19, bh56_w13_9_c20, bh56_w13_9_c21, bh56_w13_9_c22, bh56_w13_9_c23, bh56_w13_9_c24, bh56_w13_9_c25, bh56_w13_9_c26, bh56_w13_9_c27, bh56_w13_9_c28, bh56_w13_9_c29, bh56_w13_9_c30, bh56_w13_9_c31, bh56_w13_9_c32, bh56_w13_9_c33, bh56_w13_9_c34, bh56_w13_9_c35, bh56_w13_9_c36, bh56_w13_9_c37, bh56_w13_9_c38, bh56_w13_9_c39, bh56_w13_9_c40, bh56_w13_9_c41 :  std_logic;
signal bh56_w14_11_c0, bh56_w14_11_c1, bh56_w14_11_c2, bh56_w14_11_c3, bh56_w14_11_c4, bh56_w14_11_c5, bh56_w14_11_c6, bh56_w14_11_c7, bh56_w14_11_c8, bh56_w14_11_c9, bh56_w14_11_c10, bh56_w14_11_c11, bh56_w14_11_c12, bh56_w14_11_c13, bh56_w14_11_c14, bh56_w14_11_c15, bh56_w14_11_c16, bh56_w14_11_c17, bh56_w14_11_c18, bh56_w14_11_c19, bh56_w14_11_c20, bh56_w14_11_c21, bh56_w14_11_c22, bh56_w14_11_c23, bh56_w14_11_c24, bh56_w14_11_c25, bh56_w14_11_c26, bh56_w14_11_c27, bh56_w14_11_c28, bh56_w14_11_c29, bh56_w14_11_c30, bh56_w14_11_c31, bh56_w14_11_c32, bh56_w14_11_c33, bh56_w14_11_c34, bh56_w14_11_c35, bh56_w14_11_c36, bh56_w14_11_c37, bh56_w14_11_c38, bh56_w14_11_c39, bh56_w14_11_c40, bh56_w14_11_c41 :  std_logic;
signal bh56_w15_13_c0, bh56_w15_13_c1, bh56_w15_13_c2, bh56_w15_13_c3, bh56_w15_13_c4, bh56_w15_13_c5, bh56_w15_13_c6, bh56_w15_13_c7, bh56_w15_13_c8, bh56_w15_13_c9, bh56_w15_13_c10, bh56_w15_13_c11, bh56_w15_13_c12, bh56_w15_13_c13, bh56_w15_13_c14, bh56_w15_13_c15, bh56_w15_13_c16, bh56_w15_13_c17, bh56_w15_13_c18, bh56_w15_13_c19, bh56_w15_13_c20, bh56_w15_13_c21, bh56_w15_13_c22, bh56_w15_13_c23, bh56_w15_13_c24, bh56_w15_13_c25, bh56_w15_13_c26, bh56_w15_13_c27, bh56_w15_13_c28, bh56_w15_13_c29, bh56_w15_13_c30, bh56_w15_13_c31, bh56_w15_13_c32, bh56_w15_13_c33, bh56_w15_13_c34, bh56_w15_13_c35, bh56_w15_13_c36, bh56_w15_13_c37, bh56_w15_13_c38, bh56_w15_13_c39, bh56_w15_13_c40, bh56_w15_13_c41 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid266_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w12_14_c42 :  std_logic;
signal bh56_w13_10_c42 :  std_logic;
signal bh56_w14_12_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_copy267_c41, Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_copy267_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid268_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w12_15_c42 :  std_logic;
signal bh56_w13_11_c42 :  std_logic;
signal bh56_w14_13_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_copy269_c41, Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_copy269_c42 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid272_In0_c41 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid272_In1_c41 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w12_16_c42 :  std_logic;
signal bh56_w13_12_c42 :  std_logic;
signal bh56_w14_14_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_copy273_c41, Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_copy273_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid274_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w13_13_c42 :  std_logic;
signal bh56_w14_15_c42 :  std_logic;
signal bh56_w15_14_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_copy275_c41, Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_copy275_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid278_In0_c41 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_c42 :  std_logic_vector(1 downto 0);
signal bh56_w13_14_c42 :  std_logic;
signal bh56_w14_16_c42 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_copy279_c41, Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_copy279_c42 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid280_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w14_17_c42 :  std_logic;
signal bh56_w15_15_c42 :  std_logic;
signal bh56_w16_14_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_copy281_c41, Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_copy281_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid282_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w14_18_c42 :  std_logic;
signal bh56_w15_16_c42 :  std_logic;
signal bh56_w16_15_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_copy283_c41, Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_copy283_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid284_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w15_17_c42 :  std_logic;
signal bh56_w16_16_c42 :  std_logic;
signal bh56_w17_14_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_copy285_c41, Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_copy285_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid286_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w15_18_c42 :  std_logic;
signal bh56_w16_17_c42 :  std_logic;
signal bh56_w17_15_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_copy287_c41, Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_copy287_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid290_In0_c41 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid290_In1_c41 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w15_19_c42 :  std_logic;
signal bh56_w16_18_c42 :  std_logic;
signal bh56_w17_16_c42 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_copy291_c41, Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_copy291_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid292_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w16_19_c42 :  std_logic;
signal bh56_w17_17_c42 :  std_logic;
signal bh56_w18_14_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_copy293_c41, Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_copy293_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid294_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w16_20_c42 :  std_logic;
signal bh56_w17_18_c42 :  std_logic;
signal bh56_w18_15_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_copy295_c41, Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_copy295_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid296_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w17_19_c42 :  std_logic;
signal bh56_w18_16_c42 :  std_logic;
signal bh56_w19_13_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_copy297_c41, Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_copy297_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid298_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w17_20_c42 :  std_logic;
signal bh56_w18_17_c42 :  std_logic;
signal bh56_w19_14_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_copy299_c41, Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_copy299_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid300_In0_c41 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid300_In1_c41 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w17_21_c42 :  std_logic;
signal bh56_w18_18_c42 :  std_logic;
signal bh56_w19_15_c42 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_copy301_c41, Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_copy301_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid302_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w18_19_c42 :  std_logic;
signal bh56_w19_16_c42 :  std_logic;
signal bh56_w20_12_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_copy303_c41, Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_copy303_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid304_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w18_20_c42 :  std_logic;
signal bh56_w19_17_c42 :  std_logic;
signal bh56_w20_13_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_copy305_c41, Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_copy305_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid306_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w19_18_c42 :  std_logic;
signal bh56_w20_14_c42 :  std_logic;
signal bh56_w21_11_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_copy307_c41, Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_copy307_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid308_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w19_19_c42 :  std_logic;
signal bh56_w20_15_c42 :  std_logic;
signal bh56_w21_12_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_copy309_c41, Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_copy309_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid310_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w20_16_c42 :  std_logic;
signal bh56_w21_13_c42 :  std_logic;
signal bh56_w22_11_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_copy311_c41, Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_copy311_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid312_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w20_17_c42 :  std_logic;
signal bh56_w21_14_c42 :  std_logic;
signal bh56_w22_12_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_copy313_c41, Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_copy313_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid314_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w21_15_c42 :  std_logic;
signal bh56_w22_13_c42 :  std_logic;
signal bh56_w23_9_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_copy315_c41, Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_copy315_c42 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid316_In0_c41 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid316_In1_c41 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w21_16_c42 :  std_logic;
signal bh56_w22_14_c42 :  std_logic;
signal bh56_w23_10_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_copy317_c41, Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_copy317_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid318_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w22_15_c42 :  std_logic;
signal bh56_w23_11_c42 :  std_logic;
signal bh56_w24_9_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_copy319_c41, Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_copy319_c42 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid320_In0_c41 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c0, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c1, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c2, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c3, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c4, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c5, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c6, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c7, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c8, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c9, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c10, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c11, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c12, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c13, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c14, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c15, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c16, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c17, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c18, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c19, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c20, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c21, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c22, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c23, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c24, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c25, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c26, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c27, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c28, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c29, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c30, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c31, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c32, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c33, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c34, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c35, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c36, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c37, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c38, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c39, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c40, Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c41 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w22_16_c42 :  std_logic;
signal bh56_w23_12_c42 :  std_logic;
signal bh56_w24_10_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_copy321_c41, Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_copy321_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid322_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w23_13_c42 :  std_logic;
signal bh56_w24_11_c42 :  std_logic;
signal bh56_w25_8_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_copy323_c41, Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_copy323_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid324_In0_c41 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_c42 :  std_logic_vector(1 downto 0);
signal bh56_w23_14_c42 :  std_logic;
signal bh56_w24_12_c42 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_copy325_c41, Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_copy325_c42 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid326_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w24_13_c42 :  std_logic;
signal bh56_w25_9_c42 :  std_logic;
signal bh56_w26_7_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_copy327_c41, Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_copy327_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid328_In0_c41 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid328_In1_c41 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w24_14_c42 :  std_logic;
signal bh56_w25_10_c42 :  std_logic;
signal bh56_w26_8_c42 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_copy329_c41, Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_copy329_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid330_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w25_11_c42 :  std_logic;
signal bh56_w26_9_c42 :  std_logic;
signal bh56_w27_6_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_copy331_c41, Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_copy331_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid332_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w26_10_c42 :  std_logic;
signal bh56_w27_7_c42 :  std_logic;
signal bh56_w28_6_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_copy333_c41, Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_copy333_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid334_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w27_8_c42 :  std_logic;
signal bh56_w28_7_c42 :  std_logic;
signal bh56_w29_4_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_copy335_c41, Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_copy335_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid336_In0_c41 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w28_8_c42 :  std_logic;
signal bh56_w29_5_c42 :  std_logic;
signal bh56_w30_4_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_copy337_c41, Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_copy337_c42 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid338_In0_c41 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid338_In1_c41 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w29_6_c42 :  std_logic;
signal bh56_w30_5_c42 :  std_logic;
signal bh56_w31_3_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_copy339_c41, Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_copy339_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid340_In0_c41 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid340_In1_c41 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w30_6_c42 :  std_logic;
signal bh56_w31_4_c42 :  std_logic;
signal bh56_w32_2_c42 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_copy341_c41, Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_copy341_c42 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid342_In0_c41 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid342_In1_c41 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w32_3_c42 :  std_logic;
signal bh56_w33_1_c42 :  std_logic;
signal bh56_w34_1_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_copy343_c41, Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_copy343_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid344_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid344_Out0_c42 :  std_logic_vector(1 downto 0);
signal bh56_w12_17_c42, bh56_w12_17_c43 :  std_logic;
signal bh56_w13_15_c42 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid344_Out0_copy345_c42 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid346_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid346_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid346_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w13_16_c42 :  std_logic;
signal bh56_w14_19_c42 :  std_logic;
signal bh56_w15_20_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid346_Out0_copy347_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid348_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid348_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w14_20_c42 :  std_logic;
signal bh56_w15_21_c42 :  std_logic;
signal bh56_w16_21_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid348_Out0_copy349_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid350_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid350_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w15_22_c42 :  std_logic;
signal bh56_w16_22_c42 :  std_logic;
signal bh56_w17_22_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid350_Out0_copy351_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid352_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid352_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w16_23_c42 :  std_logic;
signal bh56_w17_23_c42 :  std_logic;
signal bh56_w18_21_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid352_Out0_copy353_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid354_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid354_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w17_24_c42 :  std_logic;
signal bh56_w18_22_c42 :  std_logic;
signal bh56_w19_20_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid354_Out0_copy355_c42 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid356_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid356_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid356_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w17_25_c42 :  std_logic;
signal bh56_w18_23_c42 :  std_logic;
signal bh56_w19_21_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid356_Out0_copy357_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid358_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid358_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w18_24_c42 :  std_logic;
signal bh56_w19_22_c42 :  std_logic;
signal bh56_w20_18_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid358_Out0_copy359_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid360_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid360_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w19_23_c42 :  std_logic;
signal bh56_w20_19_c42 :  std_logic;
signal bh56_w21_17_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid360_Out0_copy361_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid362_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid362_Out0_c42 :  std_logic_vector(1 downto 0);
signal bh56_w19_24_c42 :  std_logic;
signal bh56_w20_20_c42 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid362_Out0_copy363_c42 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid364_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid364_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w20_21_c42 :  std_logic;
signal bh56_w21_18_c42 :  std_logic;
signal bh56_w22_17_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid364_Out0_copy365_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid366_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid366_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w21_19_c42 :  std_logic;
signal bh56_w22_18_c42 :  std_logic;
signal bh56_w23_15_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid366_Out0_copy367_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid368_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid368_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w22_19_c42 :  std_logic;
signal bh56_w23_16_c42 :  std_logic;
signal bh56_w24_15_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid368_Out0_copy369_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid370_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid370_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w23_17_c42 :  std_logic;
signal bh56_w24_16_c42 :  std_logic;
signal bh56_w25_12_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid370_Out0_copy371_c42 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid372_In0_c42 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid265_bh56_uid372_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w24_17_c42, bh56_w24_17_c43 :  std_logic;
signal bh56_w25_13_c42 :  std_logic;
signal bh56_w26_11_c42 :  std_logic;
signal Compressor_6_3_Freq800_uid265_bh56_uid372_Out0_copy373_c42 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid374_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid374_In1_c41, Compressor_14_3_Freq800_uid271_bh56_uid374_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid374_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w25_14_c42 :  std_logic;
signal bh56_w26_12_c42 :  std_logic;
signal bh56_w27_9_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid374_Out0_copy375_c42 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid376_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c0, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c1, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c2, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c3, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c4, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c5, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c6, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c7, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c8, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c9, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c10, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c11, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c12, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c13, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c14, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c15, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c16, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c17, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c18, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c19, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c20, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c21, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c22, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c23, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c24, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c25, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c26, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c27, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c28, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c29, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c30, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c31, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c32, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c33, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c34, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c35, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c36, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c37, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c38, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c39, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c40, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c41, Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid376_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w26_13_c42, bh56_w26_13_c43 :  std_logic;
signal bh56_w27_10_c42 :  std_logic;
signal bh56_w28_9_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid376_Out0_copy377_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid378_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid378_Out0_c42 :  std_logic_vector(1 downto 0);
signal bh56_w27_11_c42 :  std_logic;
signal bh56_w28_10_c42 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid378_Out0_copy379_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid380_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid380_In1_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid380_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w28_11_c42, bh56_w28_11_c43 :  std_logic;
signal bh56_w29_7_c42 :  std_logic;
signal bh56_w30_7_c42 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid380_Out0_copy381_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid382_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid382_In1_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid382_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w30_8_c42 :  std_logic;
signal bh56_w31_5_c42 :  std_logic;
signal bh56_w32_4_c42 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid382_Out0_copy383_c42 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid384_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid384_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid384_Out0_c42 :  std_logic_vector(2 downto 0);
signal bh56_w32_5_c42 :  std_logic;
signal bh56_w33_2_c42, bh56_w33_2_c43 :  std_logic;
signal bh56_w34_2_c42 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid384_Out0_copy385_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid386_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid386_Out0_c42 :  std_logic_vector(1 downto 0);
signal bh56_w34_3_c42 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid386_Out0_copy387_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid388_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid388_In1_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w13_17_c43 :  std_logic;
signal bh56_w14_21_c43 :  std_logic;
signal bh56_w15_23_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_copy389_c42, Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_copy389_c43 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid390_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_c43 :  std_logic_vector(1 downto 0);
signal bh56_w15_24_c43 :  std_logic;
signal bh56_w16_24_c43 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_copy391_c42, Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_copy391_c43 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid392_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid392_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w16_25_c43 :  std_logic;
signal bh56_w17_26_c43 :  std_logic;
signal bh56_w18_25_c43 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_copy393_c42, Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_copy393_c43 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid394_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_c43 :  std_logic_vector(1 downto 0);
signal bh56_w17_27_c43 :  std_logic;
signal bh56_w18_26_c43 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_copy395_c42, Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_copy395_c43 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid396_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid396_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w18_27_c43 :  std_logic;
signal bh56_w19_25_c43 :  std_logic;
signal bh56_w20_22_c43 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_copy397_c42, Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_copy397_c43 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid398_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid398_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w19_26_c43 :  std_logic;
signal bh56_w20_23_c43 :  std_logic;
signal bh56_w21_20_c43 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_copy399_c42, Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_copy399_c43 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid400_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_c43 :  std_logic_vector(1 downto 0);
signal bh56_w20_24_c43 :  std_logic;
signal bh56_w21_21_c43 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_copy401_c42, Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_copy401_c43 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid402_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c0, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c1, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c2, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c3, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c4, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c5, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c6, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c7, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c8, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c9, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c10, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c11, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c12, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c13, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c14, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c15, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c16, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c17, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c18, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c19, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c20, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c21, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c22, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c23, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c24, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c25, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c26, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c27, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c28, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c29, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c30, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c31, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c32, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c33, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c34, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c35, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c36, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c37, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c38, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c39, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c40, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c41, Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w21_22_c43 :  std_logic;
signal bh56_w22_20_c43 :  std_logic;
signal bh56_w23_18_c43 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_copy403_c42, Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_copy403_c43 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid404_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_c43 :  std_logic_vector(1 downto 0);
signal bh56_w22_21_c43 :  std_logic;
signal bh56_w23_19_c43 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_copy405_c42, Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_copy405_c43 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid406_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid406_In1_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w23_20_c43 :  std_logic;
signal bh56_w24_18_c43 :  std_logic;
signal bh56_w25_15_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_copy407_c42, Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_copy407_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid408_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid408_In1_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w25_16_c43 :  std_logic;
signal bh56_w26_14_c43 :  std_logic;
signal bh56_w27_12_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_copy409_c42, Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_copy409_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid410_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid410_In1_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w27_13_c43 :  std_logic;
signal bh56_w28_12_c43 :  std_logic;
signal bh56_w29_8_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_copy411_c42, Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_copy411_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid412_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid412_In1_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w29_9_c43 :  std_logic;
signal bh56_w30_9_c43 :  std_logic;
signal bh56_w31_6_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_copy413_c42, Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_copy413_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid414_In0_c42 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid414_In1_c42 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w31_7_c43 :  std_logic;
signal bh56_w32_6_c43 :  std_logic;
signal bh56_w33_3_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_copy415_c42, Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_copy415_c43 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid416_In0_c42 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c0, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c1, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c2, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c3, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c4, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c5, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c6, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c7, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c8, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c9, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c10, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c11, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c12, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c13, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c14, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c15, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c16, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c17, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c18, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c19, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c20, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c21, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c22, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c23, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c24, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c25, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c26, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c27, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c28, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c29, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c30, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c31, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c32, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c33, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c34, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c35, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c36, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c37, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c38, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c39, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c40, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c41, Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c42 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid416_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w34_4_c43 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid416_Out0_copy417_c42, Compressor_14_3_Freq800_uid271_bh56_uid416_Out0_copy417_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid418_In0_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid418_In1_c43 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid418_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w15_25_c43 :  std_logic;
signal bh56_w16_26_c43 :  std_logic;
signal bh56_w17_28_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid418_Out0_copy419_c43 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid420_In0_c43 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid277_bh56_uid420_Out0_c43 :  std_logic_vector(1 downto 0);
signal bh56_w17_29_c43 :  std_logic;
signal bh56_w18_28_c43 :  std_logic;
signal Compressor_3_2_Freq800_uid277_bh56_uid420_Out0_copy421_c43 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid422_In0_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid422_In1_c43 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid422_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w18_29_c43 :  std_logic;
signal bh56_w19_27_c43 :  std_logic;
signal bh56_w20_25_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid422_Out0_copy423_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid424_In0_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c0, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c1, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c2, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c3, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c4, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c5, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c6, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c7, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c8, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c9, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c10, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c11, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c12, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c13, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c14, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c15, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c16, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c17, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c18, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c19, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c20, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c21, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c22, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c23, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c24, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c25, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c26, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c27, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c28, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c29, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c30, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c31, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c32, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c33, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c34, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c35, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c36, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c37, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c38, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c39, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c40, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c41, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c42, Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c43 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid424_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w20_26_c43 :  std_logic;
signal bh56_w21_23_c43 :  std_logic;
signal bh56_w22_22_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid424_Out0_copy425_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid426_In0_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid426_In1_c43 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid426_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w21_24_c43 :  std_logic;
signal bh56_w22_23_c43 :  std_logic;
signal bh56_w23_21_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid426_Out0_copy427_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid428_In0_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid428_In1_c43 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid428_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w23_22_c43 :  std_logic;
signal bh56_w24_19_c43 :  std_logic;
signal bh56_w25_17_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid428_Out0_copy429_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid430_In0_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid430_In1_c43 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid430_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w25_18_c43 :  std_logic;
signal bh56_w26_15_c43 :  std_logic;
signal bh56_w27_14_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid430_Out0_copy431_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid432_In0_c43 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid432_In1_c43 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid289_bh56_uid432_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w27_15_c43 :  std_logic;
signal bh56_w28_13_c43 :  std_logic;
signal bh56_w29_10_c43 :  std_logic;
signal Compressor_23_3_Freq800_uid289_bh56_uid432_Out0_copy433_c43 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid434_In0_c43 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid434_In1_c43 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid434_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w29_11_c43 :  std_logic;
signal bh56_w30_10_c43 :  std_logic;
signal bh56_w31_8_c43 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid434_Out0_copy435_c43 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid436_In0_c43 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid436_In1_c43 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid436_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w31_9_c43 :  std_logic;
signal bh56_w32_7_c43 :  std_logic;
signal bh56_w33_4_c43 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid436_Out0_copy437_c43 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid438_In0_c43 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid438_In1_c43 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid271_bh56_uid438_Out0_c43 :  std_logic_vector(2 downto 0);
signal bh56_w33_5_c43 :  std_logic;
signal bh56_w34_5_c43 :  std_logic;
signal Compressor_14_3_Freq800_uid271_bh56_uid438_Out0_copy439_c43 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh56_16_c43, tmp_bitheapResult_bh56_16_c44, tmp_bitheapResult_bh56_16_c45, tmp_bitheapResult_bh56_16_c46, tmp_bitheapResult_bh56_16_c47, tmp_bitheapResult_bh56_16_c48, tmp_bitheapResult_bh56_16_c49, tmp_bitheapResult_bh56_16_c50 :  std_logic_vector(16 downto 0);
signal bitheapFinalAdd_bh56_In0_c43 :  std_logic_vector(18 downto 0);
signal bitheapFinalAdd_bh56_In1_c43 :  std_logic_vector(18 downto 0);
signal bitheapFinalAdd_bh56_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh56_Out_c50 :  std_logic_vector(18 downto 0);
signal bitheapResult_bh56_c50 :  std_logic_vector(34 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_39 = '1' then
               bh56_w12_13_c39 <= bh56_w12_13_c38;
               bh56_w13_9_c39 <= bh56_w13_9_c38;
               bh56_w14_11_c39 <= bh56_w14_11_c38;
               bh56_w15_13_c39 <= bh56_w15_13_c38;
               Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c39 <= Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c38;
               Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c39 <= Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c38;
               Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c39 <= Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c38;
               Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c39 <= Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c38;
               Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c39 <= Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c38;
            end if;
            if ce_40 = '1' then
               bh56_w12_13_c40 <= bh56_w12_13_c39;
               bh56_w13_9_c40 <= bh56_w13_9_c39;
               bh56_w14_11_c40 <= bh56_w14_11_c39;
               bh56_w15_13_c40 <= bh56_w15_13_c39;
               Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c40 <= Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c39;
               Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c40 <= Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c39;
               Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c40 <= Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c39;
               Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c40 <= Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c39;
               Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c40 <= Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c39;
            end if;
            if ce_41 = '1' then
               bh56_w12_13_c41 <= bh56_w12_13_c40;
               bh56_w13_9_c41 <= bh56_w13_9_c40;
               bh56_w14_11_c41 <= bh56_w14_11_c40;
               bh56_w15_13_c41 <= bh56_w15_13_c40;
               Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c41 <= Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c40;
               Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c41 <= Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c40;
               Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c41 <= Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c40;
               Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c41 <= Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c40;
               Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c41 <= Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c40;
            end if;
            if ce_42 = '1' then
               bh56_w19_6_c42 <= bh56_w19_6_c41;
               bh56_w21_10_c42 <= bh56_w21_10_c41;
               bh56_w31_2_c42 <= bh56_w31_2_c41;
               bh56_w34_0_c42 <= bh56_w34_0_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_copy267_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_copy267_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_copy269_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_copy269_c41;
               Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_copy273_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_copy273_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_copy275_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_copy275_c41;
               Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_copy279_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_copy279_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_copy281_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_copy281_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_copy283_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_copy283_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_copy285_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_copy285_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_copy287_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_copy287_c41;
               Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_copy291_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_copy291_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_copy293_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_copy293_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_copy295_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_copy295_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_copy297_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_copy297_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_copy299_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_copy299_c41;
               Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_copy301_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_copy301_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_copy303_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_copy303_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_copy305_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_copy305_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_copy307_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_copy307_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_copy309_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_copy309_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_copy311_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_copy311_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_copy313_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_copy313_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_copy315_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_copy315_c41;
               Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_copy317_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_copy317_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_copy319_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_copy319_c41;
               Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_copy321_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_copy321_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_copy323_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_copy323_c41;
               Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_copy325_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_copy325_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_copy327_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_copy327_c41;
               Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_copy329_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_copy329_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_copy331_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_copy331_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_copy333_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_copy333_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_copy335_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_copy335_c41;
               Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_copy337_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_copy337_c41;
               Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_copy339_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_copy339_c41;
               Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_copy341_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_copy341_c41;
               Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_copy343_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_copy343_c41;
               Compressor_14_3_Freq800_uid271_bh56_uid374_In1_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid374_In1_c41;
               Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c41;
               Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c41;
               Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c41;
               Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c41;
            end if;
            if ce_43 = '1' then
               bh56_w12_17_c43 <= bh56_w12_17_c42;
               bh56_w24_17_c43 <= bh56_w24_17_c42;
               bh56_w26_13_c43 <= bh56_w26_13_c42;
               bh56_w28_11_c43 <= bh56_w28_11_c42;
               bh56_w33_2_c43 <= bh56_w33_2_c42;
               Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_copy389_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_copy389_c42;
               Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_copy391_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_copy391_c42;
               Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_copy393_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_copy393_c42;
               Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_copy395_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_copy395_c42;
               Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_copy397_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_copy397_c42;
               Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_copy399_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_copy399_c42;
               Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_copy401_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_copy401_c42;
               Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_copy403_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_copy403_c42;
               Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_copy405_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_copy405_c42;
               Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_copy407_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_copy407_c42;
               Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_copy409_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_copy409_c42;
               Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_copy411_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_copy411_c42;
               Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_copy413_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_copy413_c42;
               Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_copy415_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_copy415_c42;
               Compressor_14_3_Freq800_uid271_bh56_uid416_Out0_copy417_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid416_Out0_copy417_c42;
               Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c42;
            end if;
            if ce_44 = '1' then
               tmp_bitheapResult_bh56_16_c44 <= tmp_bitheapResult_bh56_16_c43;
            end if;
            if ce_45 = '1' then
               tmp_bitheapResult_bh56_16_c45 <= tmp_bitheapResult_bh56_16_c44;
            end if;
            if ce_46 = '1' then
               tmp_bitheapResult_bh56_16_c46 <= tmp_bitheapResult_bh56_16_c45;
            end if;
            if ce_47 = '1' then
               tmp_bitheapResult_bh56_16_c47 <= tmp_bitheapResult_bh56_16_c46;
            end if;
            if ce_48 = '1' then
               tmp_bitheapResult_bh56_16_c48 <= tmp_bitheapResult_bh56_16_c47;
            end if;
            if ce_49 = '1' then
               tmp_bitheapResult_bh56_16_c49 <= tmp_bitheapResult_bh56_16_c48;
            end if;
            if ce_50 = '1' then
               tmp_bitheapResult_bh56_16_c50 <= tmp_bitheapResult_bh56_16_c49;
            end if;
         end if;
      end process;
   XX_m55_c41 <= X ;
   YY_m55_c38 <= Y ;
   tile_0_X_c41 <= X(11 downto 11);
   tile_0_Y_c38 <= Y(1 downto 1);
   tile_0_mult: IntMultiplierLUT_1x1_Freq800_uid58
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_0_X_c41,
                 Y => tile_0_Y_c38,
                 R => tile_0_output_c41);

   tile_0_filtered_output_c41 <= unsigned(tile_0_output_c41(0 downto 0));
   bh56_w12_0_c41 <= tile_0_filtered_output_c41(0);
   tile_1_X_c41 <= X(13 downto 12);
   tile_1_Y_c38 <= Y(1 downto 0);
   tile_1_mult: IntMultiplierLUT_2x2_Freq800_uid60
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_1_X_c41,
                 Y => tile_1_Y_c38,
                 R => tile_1_output_c41);

   tile_1_filtered_output_c41 <= unsigned(tile_1_output_c41(3 downto 0));
   bh56_w12_1_c41 <= tile_1_filtered_output_c41(0);
   bh56_w13_0_c41 <= tile_1_filtered_output_c41(1);
   bh56_w14_0_c41 <= tile_1_filtered_output_c41(2);
   bh56_w15_0_c41 <= tile_1_filtered_output_c41(3);
   tile_2_X_c41 <= X(16 downto 14);
   tile_2_Y_c38 <= Y(1 downto 0);
   tile_2_mult: IntMultiplierLUT_3x2_Freq800_uid65
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_2_X_c41,
                 Y => tile_2_Y_c38,
                 R => tile_2_output_c41);

   tile_2_filtered_output_c41 <= unsigned(tile_2_output_c41(4 downto 0));
   bh56_w14_1_c41 <= tile_2_filtered_output_c41(0);
   bh56_w15_1_c41 <= tile_2_filtered_output_c41(1);
   bh56_w16_0_c41 <= tile_2_filtered_output_c41(2);
   bh56_w17_0_c41 <= tile_2_filtered_output_c41(3);
   bh56_w18_0_c41 <= tile_2_filtered_output_c41(4);
   tile_3_X_c41 <= X(10 downto 10);
   tile_3_Y_c38 <= Y(2 downto 2);
   tile_3_mult: IntMultiplierLUT_1x1_Freq800_uid70
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_3_X_c41,
                 Y => tile_3_Y_c38,
                 R => tile_3_output_c41);

   tile_3_filtered_output_c41 <= unsigned(tile_3_output_c41(0 downto 0));
   bh56_w12_2_c41 <= tile_3_filtered_output_c41(0);
   tile_4_X_c41 <= X(10 downto 9);
   tile_4_Y_c38 <= Y(3 downto 3);
   tile_4_mult: IntMultiplierLUT_2x1_Freq800_uid72
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_4_X_c41,
                 Y => tile_4_Y_c38,
                 R => tile_4_output_c41);

   tile_4_filtered_output_c41 <= unsigned(tile_4_output_c41(1 downto 0));
   bh56_w12_3_c41 <= tile_4_filtered_output_c41(0);
   bh56_w13_1_c41 <= tile_4_filtered_output_c41(1);
   tile_5_X_c41 <= X(13 downto 11);
   tile_5_Y_c38 <= Y(3 downto 2);
   tile_5_mult: IntMultiplierLUT_3x2_Freq800_uid74
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_5_X_c41,
                 Y => tile_5_Y_c38,
                 R => tile_5_output_c41);

   tile_5_filtered_output_c41 <= unsigned(tile_5_output_c41(4 downto 0));
   bh56_w13_2_c41 <= tile_5_filtered_output_c41(0);
   bh56_w14_2_c41 <= tile_5_filtered_output_c41(1);
   bh56_w15_2_c41 <= tile_5_filtered_output_c41(2);
   bh56_w16_1_c41 <= tile_5_filtered_output_c41(3);
   bh56_w17_1_c41 <= tile_5_filtered_output_c41(4);
   tile_6_X_c41 <= X(16 downto 14);
   tile_6_Y_c38 <= Y(3 downto 2);
   tile_6_mult: IntMultiplierLUT_3x2_Freq800_uid79
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_6_X_c41,
                 Y => tile_6_Y_c38,
                 R => tile_6_output_c41);

   tile_6_filtered_output_c41 <= unsigned(tile_6_output_c41(4 downto 0));
   bh56_w16_2_c41 <= tile_6_filtered_output_c41(0);
   bh56_w17_2_c41 <= tile_6_filtered_output_c41(1);
   bh56_w18_1_c41 <= tile_6_filtered_output_c41(2);
   bh56_w19_0_c41 <= tile_6_filtered_output_c41(3);
   bh56_w20_0_c41 <= tile_6_filtered_output_c41(4);
   tile_7_X_c41 <= X(7 downto 7);
   tile_7_Y_c38 <= Y(5 downto 5);
   tile_7_mult: IntMultiplierLUT_1x1_Freq800_uid84
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_7_X_c41,
                 Y => tile_7_Y_c38,
                 R => tile_7_output_c41);

   tile_7_filtered_output_c41 <= unsigned(tile_7_output_c41(0 downto 0));
   bh56_w12_4_c41 <= tile_7_filtered_output_c41(0);
   tile_8_X_c41 <= X(10 downto 8);
   tile_8_Y_c38 <= Y(5 downto 4);
   tile_8_mult: IntMultiplierLUT_3x2_Freq800_uid86
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_8_X_c41,
                 Y => tile_8_Y_c38,
                 R => tile_8_output_c41);

   tile_8_filtered_output_c41 <= unsigned(tile_8_output_c41(4 downto 0));
   bh56_w12_5_c41 <= tile_8_filtered_output_c41(0);
   bh56_w13_3_c41 <= tile_8_filtered_output_c41(1);
   bh56_w14_3_c41 <= tile_8_filtered_output_c41(2);
   bh56_w15_3_c41 <= tile_8_filtered_output_c41(3);
   bh56_w16_3_c41 <= tile_8_filtered_output_c41(4);
   tile_9_X_c41 <= X(13 downto 11);
   tile_9_Y_c38 <= Y(5 downto 4);
   tile_9_mult: IntMultiplierLUT_3x2_Freq800_uid91
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_9_X_c41,
                 Y => tile_9_Y_c38,
                 R => tile_9_output_c41);

   tile_9_filtered_output_c41 <= unsigned(tile_9_output_c41(4 downto 0));
   bh56_w15_4_c41 <= tile_9_filtered_output_c41(0);
   bh56_w16_4_c41 <= tile_9_filtered_output_c41(1);
   bh56_w17_3_c41 <= tile_9_filtered_output_c41(2);
   bh56_w18_2_c41 <= tile_9_filtered_output_c41(3);
   bh56_w19_1_c41 <= tile_9_filtered_output_c41(4);
   tile_10_X_c41 <= X(16 downto 14);
   tile_10_Y_c38 <= Y(5 downto 4);
   tile_10_mult: IntMultiplierLUT_3x2_Freq800_uid96
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_10_X_c41,
                 Y => tile_10_Y_c38,
                 R => tile_10_output_c41);

   tile_10_filtered_output_c41 <= unsigned(tile_10_output_c41(4 downto 0));
   bh56_w18_3_c41 <= tile_10_filtered_output_c41(0);
   bh56_w19_2_c41 <= tile_10_filtered_output_c41(1);
   bh56_w20_1_c41 <= tile_10_filtered_output_c41(2);
   bh56_w21_0_c41 <= tile_10_filtered_output_c41(3);
   bh56_w22_0_c41 <= tile_10_filtered_output_c41(4);
   tile_11_X_c41 <= X(5 downto 5);
   tile_11_Y_c38 <= Y(7 downto 7);
   tile_11_mult: IntMultiplierLUT_1x1_Freq800_uid101
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_11_X_c41,
                 Y => tile_11_Y_c38,
                 R => tile_11_output_c41);

   tile_11_filtered_output_c41 <= unsigned(tile_11_output_c41(0 downto 0));
   bh56_w12_6_c41 <= tile_11_filtered_output_c41(0);
   tile_12_X_c41 <= X(7 downto 6);
   tile_12_Y_c38 <= Y(7 downto 6);
   tile_12_mult: IntMultiplierLUT_2x2_Freq800_uid103
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_12_X_c41,
                 Y => tile_12_Y_c38,
                 R => tile_12_output_c41);

   tile_12_filtered_output_c41 <= unsigned(tile_12_output_c41(3 downto 0));
   bh56_w12_7_c41 <= tile_12_filtered_output_c41(0);
   bh56_w13_4_c41 <= tile_12_filtered_output_c41(1);
   bh56_w14_4_c41 <= tile_12_filtered_output_c41(2);
   bh56_w15_5_c41 <= tile_12_filtered_output_c41(3);
   tile_13_X_c41 <= X(10 downto 8);
   tile_13_Y_c38 <= Y(7 downto 6);
   tile_13_mult: IntMultiplierLUT_3x2_Freq800_uid108
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_13_X_c41,
                 Y => tile_13_Y_c38,
                 R => tile_13_output_c41);

   tile_13_filtered_output_c41 <= unsigned(tile_13_output_c41(4 downto 0));
   bh56_w14_5_c41 <= tile_13_filtered_output_c41(0);
   bh56_w15_6_c41 <= tile_13_filtered_output_c41(1);
   bh56_w16_5_c41 <= tile_13_filtered_output_c41(2);
   bh56_w17_4_c41 <= tile_13_filtered_output_c41(3);
   bh56_w18_4_c41 <= tile_13_filtered_output_c41(4);
   tile_14_X_c41 <= X(13 downto 11);
   tile_14_Y_c38 <= Y(7 downto 6);
   tile_14_mult: IntMultiplierLUT_3x2_Freq800_uid113
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_14_X_c41,
                 Y => tile_14_Y_c38,
                 R => tile_14_output_c41);

   tile_14_filtered_output_c41 <= unsigned(tile_14_output_c41(4 downto 0));
   bh56_w17_5_c41 <= tile_14_filtered_output_c41(0);
   bh56_w18_5_c41 <= tile_14_filtered_output_c41(1);
   bh56_w19_3_c41 <= tile_14_filtered_output_c41(2);
   bh56_w20_2_c41 <= tile_14_filtered_output_c41(3);
   bh56_w21_1_c41 <= tile_14_filtered_output_c41(4);
   tile_15_X_c41 <= X(16 downto 14);
   tile_15_Y_c38 <= Y(7 downto 6);
   tile_15_mult: IntMultiplierLUT_3x2_Freq800_uid118
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_15_X_c41,
                 Y => tile_15_Y_c38,
                 R => tile_15_output_c41);

   tile_15_filtered_output_c41 <= unsigned(tile_15_output_c41(4 downto 0));
   bh56_w20_3_c41 <= tile_15_filtered_output_c41(0);
   bh56_w21_2_c41 <= tile_15_filtered_output_c41(1);
   bh56_w22_1_c41 <= tile_15_filtered_output_c41(2);
   bh56_w23_0_c41 <= tile_15_filtered_output_c41(3);
   bh56_w24_0_c41 <= tile_15_filtered_output_c41(4);
   tile_16_X_c41 <= X(4 downto 4);
   tile_16_Y_c38 <= Y(8 downto 8);
   tile_16_mult: IntMultiplierLUT_1x1_Freq800_uid123
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_16_X_c41,
                 Y => tile_16_Y_c38,
                 R => tile_16_output_c41);

   tile_16_filtered_output_c41 <= unsigned(tile_16_output_c41(0 downto 0));
   bh56_w12_8_c41 <= tile_16_filtered_output_c41(0);
   tile_17_X_c41 <= X(4 downto 3);
   tile_17_Y_c38 <= Y(9 downto 9);
   tile_17_mult: IntMultiplierLUT_2x1_Freq800_uid125
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_17_X_c41,
                 Y => tile_17_Y_c38,
                 R => tile_17_output_c41);

   tile_17_filtered_output_c41 <= unsigned(tile_17_output_c41(1 downto 0));
   bh56_w12_9_c41 <= tile_17_filtered_output_c41(0);
   bh56_w13_5_c41 <= tile_17_filtered_output_c41(1);
   tile_18_X_c41 <= X(7 downto 5);
   tile_18_Y_c38 <= Y(9 downto 8);
   tile_18_mult: IntMultiplierLUT_3x2_Freq800_uid127
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_18_X_c41,
                 Y => tile_18_Y_c38,
                 R => tile_18_output_c41);

   tile_18_filtered_output_c41 <= unsigned(tile_18_output_c41(4 downto 0));
   bh56_w13_6_c41 <= tile_18_filtered_output_c41(0);
   bh56_w14_6_c41 <= tile_18_filtered_output_c41(1);
   bh56_w15_7_c41 <= tile_18_filtered_output_c41(2);
   bh56_w16_6_c41 <= tile_18_filtered_output_c41(3);
   bh56_w17_6_c41 <= tile_18_filtered_output_c41(4);
   tile_19_X_c41 <= X(10 downto 8);
   tile_19_Y_c38 <= Y(9 downto 8);
   tile_19_mult: IntMultiplierLUT_3x2_Freq800_uid132
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_19_X_c41,
                 Y => tile_19_Y_c38,
                 R => tile_19_output_c41);

   tile_19_filtered_output_c41 <= unsigned(tile_19_output_c41(4 downto 0));
   bh56_w16_7_c41 <= tile_19_filtered_output_c41(0);
   bh56_w17_7_c41 <= tile_19_filtered_output_c41(1);
   bh56_w18_6_c41 <= tile_19_filtered_output_c41(2);
   bh56_w19_4_c41 <= tile_19_filtered_output_c41(3);
   bh56_w20_4_c41 <= tile_19_filtered_output_c41(4);
   tile_20_X_c41 <= X(13 downto 11);
   tile_20_Y_c38 <= Y(9 downto 8);
   tile_20_mult: IntMultiplierLUT_3x2_Freq800_uid137
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_20_X_c41,
                 Y => tile_20_Y_c38,
                 R => tile_20_output_c41);

   tile_20_filtered_output_c41 <= unsigned(tile_20_output_c41(4 downto 0));
   bh56_w19_5_c41 <= tile_20_filtered_output_c41(0);
   bh56_w20_5_c41 <= tile_20_filtered_output_c41(1);
   bh56_w21_3_c41 <= tile_20_filtered_output_c41(2);
   bh56_w22_2_c41 <= tile_20_filtered_output_c41(3);
   bh56_w23_1_c41 <= tile_20_filtered_output_c41(4);
   tile_21_X_c41 <= X(16 downto 14);
   tile_21_Y_c38 <= Y(9 downto 8);
   tile_21_mult: IntMultiplierLUT_3x2_Freq800_uid142
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_21_X_c41,
                 Y => tile_21_Y_c38,
                 R => tile_21_output_c41);

   tile_21_filtered_output_c41 <= unsigned(tile_21_output_c41(4 downto 0));
   bh56_w22_3_c41 <= tile_21_filtered_output_c41(0);
   bh56_w23_2_c41 <= tile_21_filtered_output_c41(1);
   bh56_w24_1_c41 <= tile_21_filtered_output_c41(2);
   bh56_w25_0_c41 <= tile_21_filtered_output_c41(3);
   bh56_w26_0_c41 <= tile_21_filtered_output_c41(4);
   tile_22_X_c41 <= X(1 downto 1);
   tile_22_Y_c38 <= Y(11 downto 11);
   tile_22_mult: IntMultiplierLUT_1x1_Freq800_uid147
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_22_X_c41,
                 Y => tile_22_Y_c38,
                 R => tile_22_output_c41);

   tile_22_filtered_output_c41 <= unsigned(tile_22_output_c41(0 downto 0));
   bh56_w12_10_c41 <= tile_22_filtered_output_c41(0);
   tile_23_X_c41 <= X(4 downto 2);
   tile_23_Y_c38 <= Y(11 downto 10);
   tile_23_mult: IntMultiplierLUT_3x2_Freq800_uid149
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_23_X_c41,
                 Y => tile_23_Y_c38,
                 R => tile_23_output_c41);

   tile_23_filtered_output_c41 <= unsigned(tile_23_output_c41(4 downto 0));
   bh56_w12_11_c41 <= tile_23_filtered_output_c41(0);
   bh56_w13_7_c41 <= tile_23_filtered_output_c41(1);
   bh56_w14_7_c41 <= tile_23_filtered_output_c41(2);
   bh56_w15_8_c41 <= tile_23_filtered_output_c41(3);
   bh56_w16_8_c41 <= tile_23_filtered_output_c41(4);
   tile_24_X_c41 <= X(7 downto 5);
   tile_24_Y_c38 <= Y(11 downto 10);
   tile_24_mult: IntMultiplierLUT_3x2_Freq800_uid154
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_24_X_c41,
                 Y => tile_24_Y_c38,
                 R => tile_24_output_c41);

   tile_24_filtered_output_c41 <= unsigned(tile_24_output_c41(4 downto 0));
   bh56_w15_9_c41 <= tile_24_filtered_output_c41(0);
   bh56_w16_9_c41 <= tile_24_filtered_output_c41(1);
   bh56_w17_8_c41 <= tile_24_filtered_output_c41(2);
   bh56_w18_7_c41 <= tile_24_filtered_output_c41(3);
   bh56_w19_6_c41 <= tile_24_filtered_output_c41(4);
   tile_25_X_c41 <= X(10 downto 8);
   tile_25_Y_c38 <= Y(11 downto 10);
   tile_25_mult: IntMultiplierLUT_3x2_Freq800_uid159
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_25_X_c41,
                 Y => tile_25_Y_c38,
                 R => tile_25_output_c41);

   tile_25_filtered_output_c41 <= unsigned(tile_25_output_c41(4 downto 0));
   bh56_w18_8_c41 <= tile_25_filtered_output_c41(0);
   bh56_w19_7_c41 <= tile_25_filtered_output_c41(1);
   bh56_w20_6_c41 <= tile_25_filtered_output_c41(2);
   bh56_w21_4_c41 <= tile_25_filtered_output_c41(3);
   bh56_w22_4_c41 <= tile_25_filtered_output_c41(4);
   tile_26_X_c41 <= X(13 downto 11);
   tile_26_Y_c38 <= Y(11 downto 10);
   tile_26_mult: IntMultiplierLUT_3x2_Freq800_uid164
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_26_X_c41,
                 Y => tile_26_Y_c38,
                 R => tile_26_output_c41);

   tile_26_filtered_output_c41 <= unsigned(tile_26_output_c41(4 downto 0));
   bh56_w21_5_c41 <= tile_26_filtered_output_c41(0);
   bh56_w22_5_c41 <= tile_26_filtered_output_c41(1);
   bh56_w23_3_c41 <= tile_26_filtered_output_c41(2);
   bh56_w24_2_c41 <= tile_26_filtered_output_c41(3);
   bh56_w25_1_c41 <= tile_26_filtered_output_c41(4);
   tile_27_X_c41 <= X(16 downto 14);
   tile_27_Y_c38 <= Y(11 downto 10);
   tile_27_mult: IntMultiplierLUT_3x2_Freq800_uid169
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_27_X_c41,
                 Y => tile_27_Y_c38,
                 R => tile_27_output_c41);

   tile_27_filtered_output_c41 <= unsigned(tile_27_output_c41(4 downto 0));
   bh56_w24_3_c41 <= tile_27_filtered_output_c41(0);
   bh56_w25_2_c41 <= tile_27_filtered_output_c41(1);
   bh56_w26_1_c41 <= tile_27_filtered_output_c41(2);
   bh56_w27_0_c41 <= tile_27_filtered_output_c41(3);
   bh56_w28_0_c41 <= tile_27_filtered_output_c41(4);
   tile_28_X_c41 <= X(1 downto 0);
   tile_28_Y_c38 <= Y(13 downto 12);
   tile_28_mult: IntMultiplierLUT_2x2_Freq800_uid174
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_28_X_c41,
                 Y => tile_28_Y_c38,
                 R => tile_28_output_c41);

   tile_28_filtered_output_c41 <= unsigned(tile_28_output_c41(3 downto 0));
   bh56_w12_12_c41 <= tile_28_filtered_output_c41(0);
   bh56_w13_8_c41 <= tile_28_filtered_output_c41(1);
   bh56_w14_8_c41 <= tile_28_filtered_output_c41(2);
   bh56_w15_10_c41 <= tile_28_filtered_output_c41(3);
   tile_29_X_c41 <= X(4 downto 2);
   tile_29_Y_c38 <= Y(13 downto 12);
   tile_29_mult: IntMultiplierLUT_3x2_Freq800_uid179
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_29_X_c41,
                 Y => tile_29_Y_c38,
                 R => tile_29_output_c41);

   tile_29_filtered_output_c41 <= unsigned(tile_29_output_c41(4 downto 0));
   bh56_w14_9_c41 <= tile_29_filtered_output_c41(0);
   bh56_w15_11_c41 <= tile_29_filtered_output_c41(1);
   bh56_w16_10_c41 <= tile_29_filtered_output_c41(2);
   bh56_w17_9_c41 <= tile_29_filtered_output_c41(3);
   bh56_w18_9_c41 <= tile_29_filtered_output_c41(4);
   tile_30_X_c41 <= X(7 downto 5);
   tile_30_Y_c38 <= Y(13 downto 12);
   tile_30_mult: IntMultiplierLUT_3x2_Freq800_uid184
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_30_X_c41,
                 Y => tile_30_Y_c38,
                 R => tile_30_output_c41);

   tile_30_filtered_output_c41 <= unsigned(tile_30_output_c41(4 downto 0));
   bh56_w17_10_c41 <= tile_30_filtered_output_c41(0);
   bh56_w18_10_c41 <= tile_30_filtered_output_c41(1);
   bh56_w19_8_c41 <= tile_30_filtered_output_c41(2);
   bh56_w20_7_c41 <= tile_30_filtered_output_c41(3);
   bh56_w21_6_c41 <= tile_30_filtered_output_c41(4);
   tile_31_X_c41 <= X(10 downto 8);
   tile_31_Y_c38 <= Y(13 downto 12);
   tile_31_mult: IntMultiplierLUT_3x2_Freq800_uid189
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_31_X_c41,
                 Y => tile_31_Y_c38,
                 R => tile_31_output_c41);

   tile_31_filtered_output_c41 <= unsigned(tile_31_output_c41(4 downto 0));
   bh56_w20_8_c41 <= tile_31_filtered_output_c41(0);
   bh56_w21_7_c41 <= tile_31_filtered_output_c41(1);
   bh56_w22_6_c41 <= tile_31_filtered_output_c41(2);
   bh56_w23_4_c41 <= tile_31_filtered_output_c41(3);
   bh56_w24_4_c41 <= tile_31_filtered_output_c41(4);
   tile_32_X_c41 <= X(13 downto 11);
   tile_32_Y_c38 <= Y(13 downto 12);
   tile_32_mult: IntMultiplierLUT_3x2_Freq800_uid194
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_32_X_c41,
                 Y => tile_32_Y_c38,
                 R => tile_32_output_c41);

   tile_32_filtered_output_c41 <= unsigned(tile_32_output_c41(4 downto 0));
   bh56_w23_5_c41 <= tile_32_filtered_output_c41(0);
   bh56_w24_5_c41 <= tile_32_filtered_output_c41(1);
   bh56_w25_3_c41 <= tile_32_filtered_output_c41(2);
   bh56_w26_2_c41 <= tile_32_filtered_output_c41(3);
   bh56_w27_1_c41 <= tile_32_filtered_output_c41(4);
   tile_33_X_c41 <= X(16 downto 14);
   tile_33_Y_c38 <= Y(13 downto 12);
   tile_33_mult: IntMultiplierLUT_3x2_Freq800_uid199
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_33_X_c41,
                 Y => tile_33_Y_c38,
                 R => tile_33_output_c41);

   tile_33_filtered_output_c41 <= unsigned(tile_33_output_c41(4 downto 0));
   bh56_w26_3_c41 <= tile_33_filtered_output_c41(0);
   bh56_w27_2_c41 <= tile_33_filtered_output_c41(1);
   bh56_w28_1_c41 <= tile_33_filtered_output_c41(2);
   bh56_w29_0_c41 <= tile_33_filtered_output_c41(3);
   bh56_w30_0_c41 <= tile_33_filtered_output_c41(4);
   tile_34_X_c41 <= X(1 downto 0);
   tile_34_Y_c38 <= Y(15 downto 14);
   tile_34_mult: IntMultiplierLUT_2x2_Freq800_uid204
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_34_X_c41,
                 Y => tile_34_Y_c38,
                 R => tile_34_output_c41);

   tile_34_filtered_output_c41 <= unsigned(tile_34_output_c41(3 downto 0));
   bh56_w14_10_c41 <= tile_34_filtered_output_c41(0);
   bh56_w15_12_c41 <= tile_34_filtered_output_c41(1);
   bh56_w16_11_c41 <= tile_34_filtered_output_c41(2);
   bh56_w17_11_c41 <= tile_34_filtered_output_c41(3);
   tile_35_X_c41 <= X(4 downto 2);
   tile_35_Y_c38 <= Y(15 downto 14);
   tile_35_mult: IntMultiplierLUT_3x2_Freq800_uid209
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_35_X_c41,
                 Y => tile_35_Y_c38,
                 R => tile_35_output_c41);

   tile_35_filtered_output_c41 <= unsigned(tile_35_output_c41(4 downto 0));
   bh56_w16_12_c41 <= tile_35_filtered_output_c41(0);
   bh56_w17_12_c41 <= tile_35_filtered_output_c41(1);
   bh56_w18_11_c41 <= tile_35_filtered_output_c41(2);
   bh56_w19_9_c41 <= tile_35_filtered_output_c41(3);
   bh56_w20_9_c41 <= tile_35_filtered_output_c41(4);
   tile_36_X_c41 <= X(7 downto 5);
   tile_36_Y_c38 <= Y(15 downto 14);
   tile_36_mult: IntMultiplierLUT_3x2_Freq800_uid214
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_36_X_c41,
                 Y => tile_36_Y_c38,
                 R => tile_36_output_c41);

   tile_36_filtered_output_c41 <= unsigned(tile_36_output_c41(4 downto 0));
   bh56_w19_10_c41 <= tile_36_filtered_output_c41(0);
   bh56_w20_10_c41 <= tile_36_filtered_output_c41(1);
   bh56_w21_8_c41 <= tile_36_filtered_output_c41(2);
   bh56_w22_7_c41 <= tile_36_filtered_output_c41(3);
   bh56_w23_6_c41 <= tile_36_filtered_output_c41(4);
   tile_37_X_c41 <= X(10 downto 8);
   tile_37_Y_c38 <= Y(15 downto 14);
   tile_37_mult: IntMultiplierLUT_3x2_Freq800_uid219
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_37_X_c41,
                 Y => tile_37_Y_c38,
                 R => tile_37_output_c41);

   tile_37_filtered_output_c41 <= unsigned(tile_37_output_c41(4 downto 0));
   bh56_w22_8_c41 <= tile_37_filtered_output_c41(0);
   bh56_w23_7_c41 <= tile_37_filtered_output_c41(1);
   bh56_w24_6_c41 <= tile_37_filtered_output_c41(2);
   bh56_w25_4_c41 <= tile_37_filtered_output_c41(3);
   bh56_w26_4_c41 <= tile_37_filtered_output_c41(4);
   tile_38_X_c41 <= X(13 downto 11);
   tile_38_Y_c38 <= Y(15 downto 14);
   tile_38_mult: IntMultiplierLUT_3x2_Freq800_uid224
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_38_X_c41,
                 Y => tile_38_Y_c38,
                 R => tile_38_output_c41);

   tile_38_filtered_output_c41 <= unsigned(tile_38_output_c41(4 downto 0));
   bh56_w25_5_c41 <= tile_38_filtered_output_c41(0);
   bh56_w26_5_c41 <= tile_38_filtered_output_c41(1);
   bh56_w27_3_c41 <= tile_38_filtered_output_c41(2);
   bh56_w28_2_c41 <= tile_38_filtered_output_c41(3);
   bh56_w29_1_c41 <= tile_38_filtered_output_c41(4);
   tile_39_X_c41 <= X(16 downto 14);
   tile_39_Y_c38 <= Y(15 downto 14);
   tile_39_mult: IntMultiplierLUT_3x2_Freq800_uid229
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_39_X_c41,
                 Y => tile_39_Y_c38,
                 R => tile_39_output_c41);

   tile_39_filtered_output_c41 <= unsigned(tile_39_output_c41(4 downto 0));
   bh56_w28_3_c41 <= tile_39_filtered_output_c41(0);
   bh56_w29_2_c41 <= tile_39_filtered_output_c41(1);
   bh56_w30_1_c41 <= tile_39_filtered_output_c41(2);
   bh56_w31_0_c41 <= tile_39_filtered_output_c41(3);
   bh56_w32_0_c41 <= tile_39_filtered_output_c41(4);
   tile_40_X_c41 <= X(1 downto 0);
   tile_40_Y_c38 <= Y(17 downto 16);
   tile_40_mult: IntMultiplierLUT_2x2_Freq800_uid234
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_40_X_c41,
                 Y => tile_40_Y_c38,
                 R => tile_40_output_c41);

   tile_40_filtered_output_c41 <= unsigned(tile_40_output_c41(3 downto 0));
   bh56_w16_13_c41 <= tile_40_filtered_output_c41(0);
   bh56_w17_13_c41 <= tile_40_filtered_output_c41(1);
   bh56_w18_12_c41 <= tile_40_filtered_output_c41(2);
   bh56_w19_11_c41 <= tile_40_filtered_output_c41(3);
   tile_41_X_c41 <= X(4 downto 2);
   tile_41_Y_c38 <= Y(17 downto 16);
   tile_41_mult: IntMultiplierLUT_3x2_Freq800_uid239
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_41_X_c41,
                 Y => tile_41_Y_c38,
                 R => tile_41_output_c41);

   tile_41_filtered_output_c41 <= unsigned(tile_41_output_c41(4 downto 0));
   bh56_w18_13_c41 <= tile_41_filtered_output_c41(0);
   bh56_w19_12_c41 <= tile_41_filtered_output_c41(1);
   bh56_w20_11_c41 <= tile_41_filtered_output_c41(2);
   bh56_w21_9_c41 <= tile_41_filtered_output_c41(3);
   bh56_w22_9_c41 <= tile_41_filtered_output_c41(4);
   tile_42_X_c41 <= X(7 downto 5);
   tile_42_Y_c38 <= Y(17 downto 16);
   tile_42_mult: IntMultiplierLUT_3x2_Freq800_uid244
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_42_X_c41,
                 Y => tile_42_Y_c38,
                 R => tile_42_output_c41);

   tile_42_filtered_output_c41 <= unsigned(tile_42_output_c41(4 downto 0));
   bh56_w21_10_c41 <= tile_42_filtered_output_c41(0);
   bh56_w22_10_c41 <= tile_42_filtered_output_c41(1);
   bh56_w23_8_c41 <= tile_42_filtered_output_c41(2);
   bh56_w24_7_c41 <= tile_42_filtered_output_c41(3);
   bh56_w25_6_c41 <= tile_42_filtered_output_c41(4);
   tile_43_X_c41 <= X(10 downto 8);
   tile_43_Y_c38 <= Y(17 downto 16);
   tile_43_mult: IntMultiplierLUT_3x2_Freq800_uid249
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_43_X_c41,
                 Y => tile_43_Y_c38,
                 R => tile_43_output_c41);

   tile_43_filtered_output_c41 <= unsigned(tile_43_output_c41(4 downto 0));
   bh56_w24_8_c41 <= tile_43_filtered_output_c41(0);
   bh56_w25_7_c41 <= tile_43_filtered_output_c41(1);
   bh56_w26_6_c41 <= tile_43_filtered_output_c41(2);
   bh56_w27_4_c41 <= tile_43_filtered_output_c41(3);
   bh56_w28_4_c41 <= tile_43_filtered_output_c41(4);
   tile_44_X_c41 <= X(13 downto 11);
   tile_44_Y_c38 <= Y(17 downto 16);
   tile_44_mult: IntMultiplierLUT_3x2_Freq800_uid254
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_44_X_c41,
                 Y => tile_44_Y_c38,
                 R => tile_44_output_c41);

   tile_44_filtered_output_c41 <= unsigned(tile_44_output_c41(4 downto 0));
   bh56_w27_5_c41 <= tile_44_filtered_output_c41(0);
   bh56_w28_5_c41 <= tile_44_filtered_output_c41(1);
   bh56_w29_3_c41 <= tile_44_filtered_output_c41(2);
   bh56_w30_2_c41 <= tile_44_filtered_output_c41(3);
   bh56_w31_1_c41 <= tile_44_filtered_output_c41(4);
   tile_45_X_c41 <= X(16 downto 14);
   tile_45_Y_c38 <= Y(17 downto 16);
   tile_45_mult: IntMultiplierLUT_3x2_Freq800_uid259
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 X => tile_45_X_c41,
                 Y => tile_45_Y_c38,
                 R => tile_45_output_c41);

   tile_45_filtered_output_c41 <= unsigned(tile_45_output_c41(4 downto 0));
   bh56_w30_3_c41 <= tile_45_filtered_output_c41(0);
   bh56_w31_2_c41 <= tile_45_filtered_output_c41(1);
   bh56_w32_1_c41 <= tile_45_filtered_output_c41(2);
   bh56_w33_0_c41 <= tile_45_filtered_output_c41(3);
   bh56_w34_0_c41 <= tile_45_filtered_output_c41(4);

   -- Adding the constant bits 
   bh56_w12_13_c0 <= '1';
   bh56_w13_9_c0 <= '1';
   bh56_w14_11_c0 <= '1';
   bh56_w15_13_c0 <= '1';


   Compressor_6_3_Freq800_uid265_bh56_uid266_In0_c41 <= "" & bh56_w12_0_c41 & bh56_w12_1_c41 & bh56_w12_2_c41 & bh56_w12_3_c41 & "0" & "0";
   bh56_w12_14_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_c42(0);
   bh56_w13_10_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_c42(1);
   bh56_w14_12_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid266: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid266_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_copy267_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid266_Out0_copy267_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid268_In0_c41 <= "" & bh56_w12_4_c41 & bh56_w12_5_c41 & bh56_w12_6_c41 & bh56_w12_7_c41 & bh56_w12_8_c41 & bh56_w12_9_c41;
   bh56_w12_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_c42(0);
   bh56_w13_11_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_c42(1);
   bh56_w14_13_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid268: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid268_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_copy269_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid268_Out0_copy269_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid272_In0_c41 <= "" & bh56_w12_10_c41 & bh56_w12_11_c41 & bh56_w12_12_c41 & bh56_w12_13_c41;
   Compressor_14_3_Freq800_uid271_bh56_uid272_In1_c41 <= "" & bh56_w13_0_c41;
   bh56_w12_16_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_c42(0);
   bh56_w13_12_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_c42(1);
   bh56_w14_14_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid272: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid272_In0_c41,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid272_In1_c41,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_copy273_c41);
   Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid272_Out0_copy273_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid274_In0_c41 <= "" & bh56_w13_1_c41 & bh56_w13_2_c41 & bh56_w13_3_c41 & bh56_w13_4_c41 & bh56_w13_5_c41 & bh56_w13_6_c41;
   bh56_w13_13_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_c42(0);
   bh56_w14_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_c42(1);
   bh56_w15_14_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid274: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid274_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_copy275_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid274_Out0_copy275_c42; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid278_In0_c41 <= "" & bh56_w13_7_c41 & bh56_w13_8_c41 & bh56_w13_9_c41;
   bh56_w13_14_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_c42(0);
   bh56_w14_16_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_c42(1);
   Compressor_3_2_Freq800_uid277_uid278: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid278_In0_c41,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_copy279_c41);
   Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid278_Out0_copy279_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid280_In0_c41 <= "" & bh56_w14_8_c41 & bh56_w14_11_c41 & bh56_w14_10_c41 & bh56_w14_9_c41 & bh56_w14_0_c41 & bh56_w14_7_c41;
   bh56_w14_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_c42(0);
   bh56_w15_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_c42(1);
   bh56_w16_14_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid280: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid280_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_copy281_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid280_Out0_copy281_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid282_In0_c41 <= "" & bh56_w14_1_c41 & bh56_w14_2_c41 & bh56_w14_3_c41 & bh56_w14_4_c41 & bh56_w14_5_c41 & bh56_w14_6_c41;
   bh56_w14_18_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_c42(0);
   bh56_w15_16_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_c42(1);
   bh56_w16_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid282: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid282_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_copy283_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid282_Out0_copy283_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid284_In0_c41 <= "" & bh56_w15_8_c41 & bh56_w15_13_c41 & bh56_w15_12_c41 & bh56_w15_11_c41 & bh56_w15_10_c41 & "0";
   bh56_w15_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_c42(0);
   bh56_w16_16_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_c42(1);
   bh56_w17_14_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid284: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid284_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_copy285_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid284_Out0_copy285_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid286_In0_c41 <= "" & bh56_w15_0_c41 & bh56_w15_1_c41 & bh56_w15_2_c41 & bh56_w15_3_c41 & bh56_w15_4_c41 & bh56_w15_5_c41;
   bh56_w15_18_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_c42(0);
   bh56_w16_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_c42(1);
   bh56_w17_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid286: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid286_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_copy287_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid286_Out0_copy287_c42; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid290_In0_c41 <= "" & bh56_w15_9_c41 & bh56_w15_7_c41 & bh56_w15_6_c41;
   Compressor_23_3_Freq800_uid289_bh56_uid290_In1_c41 <= "" & bh56_w16_0_c41 & bh56_w16_1_c41;
   bh56_w15_19_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_c42(0);
   bh56_w16_18_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_c42(1);
   bh56_w17_16_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_c42(2);
   Compressor_23_3_Freq800_uid289_uid290: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid290_In0_c41,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid290_In1_c41,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_copy291_c41);
   Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid290_Out0_copy291_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid292_In0_c41 <= "" & bh56_w16_8_c41 & bh56_w16_13_c41 & bh56_w16_12_c41 & bh56_w16_11_c41 & bh56_w16_10_c41 & bh56_w16_9_c41;
   bh56_w16_19_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_c42(0);
   bh56_w17_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_c42(1);
   bh56_w18_14_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid292: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid292_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_copy293_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid292_Out0_copy293_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid294_In0_c41 <= "" & bh56_w16_2_c41 & bh56_w16_3_c41 & bh56_w16_4_c41 & bh56_w16_5_c41 & bh56_w16_6_c41 & bh56_w16_7_c41;
   bh56_w16_20_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_c42(0);
   bh56_w17_18_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_c42(1);
   bh56_w18_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid294: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid294_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_copy295_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid294_Out0_copy295_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid296_In0_c41 <= "" & bh56_w17_8_c41 & bh56_w17_13_c41 & bh56_w17_12_c41 & bh56_w17_11_c41 & bh56_w17_10_c41 & "0";
   bh56_w17_19_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_c42(0);
   bh56_w18_16_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_c42(1);
   bh56_w19_13_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid296: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid296_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_copy297_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid296_Out0_copy297_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid298_In0_c41 <= "" & bh56_w17_0_c41 & bh56_w17_1_c41 & bh56_w17_2_c41 & bh56_w17_3_c41 & bh56_w17_4_c41 & bh56_w17_5_c41;
   bh56_w17_20_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_c42(0);
   bh56_w18_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_c42(1);
   bh56_w19_14_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid298: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid298_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_copy299_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid298_Out0_copy299_c42; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid300_In0_c41 <= "" & bh56_w17_9_c41 & bh56_w17_7_c41 & bh56_w17_6_c41;
   Compressor_23_3_Freq800_uid289_bh56_uid300_In1_c41 <= "" & bh56_w18_0_c41 & bh56_w18_1_c41;
   bh56_w17_21_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_c42(0);
   bh56_w18_18_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_c42(1);
   bh56_w19_15_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_c42(2);
   Compressor_23_3_Freq800_uid289_uid300: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid300_In0_c41,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid300_In1_c41,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_copy301_c41);
   Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid300_Out0_copy301_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid302_In0_c41 <= "" & bh56_w18_8_c41 & bh56_w18_13_c41 & bh56_w18_12_c41 & bh56_w18_11_c41 & bh56_w18_10_c41 & bh56_w18_9_c41;
   bh56_w18_19_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_c42(0);
   bh56_w19_16_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_c42(1);
   bh56_w20_12_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid302: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid302_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_copy303_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid302_Out0_copy303_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid304_In0_c41 <= "" & bh56_w18_2_c41 & bh56_w18_3_c41 & bh56_w18_4_c41 & bh56_w18_5_c41 & bh56_w18_6_c41 & bh56_w18_7_c41;
   bh56_w18_20_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_c42(0);
   bh56_w19_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_c42(1);
   bh56_w20_13_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid304: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid304_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_copy305_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid304_Out0_copy305_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid306_In0_c41 <= "" & bh56_w19_0_c41 & bh56_w19_1_c41 & bh56_w19_2_c41 & bh56_w19_3_c41 & bh56_w19_4_c41 & bh56_w19_5_c41;
   bh56_w19_18_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_c42(0);
   bh56_w20_14_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_c42(1);
   bh56_w21_11_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid306: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid306_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_copy307_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid306_Out0_copy307_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid308_In0_c41 <= "" & bh56_w19_8_c41 & bh56_w19_12_c41 & bh56_w19_11_c41 & bh56_w19_10_c41 & bh56_w19_9_c41 & bh56_w19_7_c41;
   bh56_w19_19_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_c42(0);
   bh56_w20_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_c42(1);
   bh56_w21_12_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid308: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid308_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_copy309_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid308_Out0_copy309_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid310_In0_c41 <= "" & bh56_w20_0_c41 & bh56_w20_1_c41 & bh56_w20_2_c41 & bh56_w20_3_c41 & bh56_w20_4_c41 & bh56_w20_5_c41;
   bh56_w20_16_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_c42(0);
   bh56_w21_13_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_c42(1);
   bh56_w22_11_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid310: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid310_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_copy311_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid310_Out0_copy311_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid312_In0_c41 <= "" & bh56_w20_8_c41 & bh56_w20_11_c41 & bh56_w20_10_c41 & bh56_w20_9_c41 & bh56_w20_7_c41 & bh56_w20_6_c41;
   bh56_w20_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_c42(0);
   bh56_w21_14_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_c42(1);
   bh56_w22_12_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid312: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid312_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_copy313_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid312_Out0_copy313_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid314_In0_c41 <= "" & bh56_w21_0_c41 & bh56_w21_1_c41 & bh56_w21_2_c41 & bh56_w21_3_c41 & bh56_w21_4_c41 & bh56_w21_5_c41;
   bh56_w21_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_c42(0);
   bh56_w22_13_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_c42(1);
   bh56_w23_9_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid314: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid314_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_copy315_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid314_Out0_copy315_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid316_In0_c41 <= "" & bh56_w21_6_c41 & bh56_w21_7_c41 & bh56_w21_8_c41 & bh56_w21_9_c41;
   Compressor_14_3_Freq800_uid271_bh56_uid316_In1_c41 <= "" & bh56_w22_0_c41;
   bh56_w21_16_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_c42(0);
   bh56_w22_14_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_c42(1);
   bh56_w23_10_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid316: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid316_In0_c41,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid316_In1_c41,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_copy317_c41);
   Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid316_Out0_copy317_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid318_In0_c41 <= "" & bh56_w22_1_c41 & bh56_w22_2_c41 & bh56_w22_3_c41 & bh56_w22_4_c41 & bh56_w22_5_c41 & bh56_w22_6_c41;
   bh56_w22_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_c42(0);
   bh56_w23_11_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_c42(1);
   bh56_w24_9_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid318: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid318_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_copy319_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid318_Out0_copy319_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid320_In0_c41 <= "" & bh56_w22_7_c41 & bh56_w22_8_c41 & bh56_w22_9_c41 & bh56_w22_10_c41;
   Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c0 <= "" & "0";
   bh56_w22_16_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_c42(0);
   bh56_w23_12_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_c42(1);
   bh56_w24_10_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid320: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid320_In0_c41,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid320_In1_c41,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_copy321_c41);
   Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid320_Out0_copy321_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid322_In0_c41 <= "" & bh56_w23_0_c41 & bh56_w23_1_c41 & bh56_w23_2_c41 & bh56_w23_3_c41 & bh56_w23_4_c41 & bh56_w23_5_c41;
   bh56_w23_13_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_c42(0);
   bh56_w24_11_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_c42(1);
   bh56_w25_8_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid322: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid322_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_copy323_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid322_Out0_copy323_c42; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid324_In0_c41 <= "" & bh56_w23_6_c41 & bh56_w23_7_c41 & bh56_w23_8_c41;
   bh56_w23_14_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_c42(0);
   bh56_w24_12_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_c42(1);
   Compressor_3_2_Freq800_uid277_uid324: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid324_In0_c41,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_copy325_c41);
   Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid324_Out0_copy325_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid326_In0_c41 <= "" & bh56_w24_0_c41 & bh56_w24_1_c41 & bh56_w24_2_c41 & bh56_w24_3_c41 & bh56_w24_4_c41 & bh56_w24_5_c41;
   bh56_w24_13_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_c42(0);
   bh56_w25_9_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_c42(1);
   bh56_w26_7_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid326: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid326_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_copy327_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid326_Out0_copy327_c42; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid328_In0_c41 <= "" & bh56_w24_6_c41 & bh56_w24_7_c41 & bh56_w24_8_c41;
   Compressor_23_3_Freq800_uid289_bh56_uid328_In1_c41 <= "" & bh56_w25_0_c41 & bh56_w25_1_c41;
   bh56_w24_14_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_c42(0);
   bh56_w25_10_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_c42(1);
   bh56_w26_8_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_c42(2);
   Compressor_23_3_Freq800_uid289_uid328: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid328_In0_c41,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid328_In1_c41,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_copy329_c41);
   Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid328_Out0_copy329_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid330_In0_c41 <= "" & bh56_w25_2_c41 & bh56_w25_3_c41 & bh56_w25_4_c41 & bh56_w25_5_c41 & bh56_w25_6_c41 & bh56_w25_7_c41;
   bh56_w25_11_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_c42(0);
   bh56_w26_9_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_c42(1);
   bh56_w27_6_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid330: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid330_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_copy331_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid330_Out0_copy331_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid332_In0_c41 <= "" & bh56_w26_0_c41 & bh56_w26_1_c41 & bh56_w26_2_c41 & bh56_w26_3_c41 & bh56_w26_4_c41 & bh56_w26_5_c41;
   bh56_w26_10_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_c42(0);
   bh56_w27_7_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_c42(1);
   bh56_w28_6_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid332: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid332_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_copy333_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid332_Out0_copy333_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid334_In0_c41 <= "" & bh56_w27_0_c41 & bh56_w27_1_c41 & bh56_w27_2_c41 & bh56_w27_3_c41 & bh56_w27_4_c41 & bh56_w27_5_c41;
   bh56_w27_8_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_c42(0);
   bh56_w28_7_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_c42(1);
   bh56_w29_4_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid334: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid334_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_copy335_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid334_Out0_copy335_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid336_In0_c41 <= "" & bh56_w28_0_c41 & bh56_w28_1_c41 & bh56_w28_2_c41 & bh56_w28_3_c41 & bh56_w28_4_c41 & bh56_w28_5_c41;
   bh56_w28_8_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_c42(0);
   bh56_w29_5_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_c42(1);
   bh56_w30_4_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid336: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid336_In0_c41,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_copy337_c41);
   Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid336_Out0_copy337_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid338_In0_c41 <= "" & bh56_w29_0_c41 & bh56_w29_1_c41 & bh56_w29_2_c41 & bh56_w29_3_c41;
   Compressor_14_3_Freq800_uid271_bh56_uid338_In1_c41 <= "" & bh56_w30_0_c41;
   bh56_w29_6_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_c42(0);
   bh56_w30_5_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_c42(1);
   bh56_w31_3_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid338: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid338_In0_c41,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid338_In1_c41,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_copy339_c41);
   Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid338_Out0_copy339_c42; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid340_In0_c41 <= "" & bh56_w30_1_c41 & bh56_w30_2_c41 & bh56_w30_3_c41;
   Compressor_23_3_Freq800_uid289_bh56_uid340_In1_c41 <= "" & bh56_w31_0_c41 & bh56_w31_1_c41;
   bh56_w30_6_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_c42(0);
   bh56_w31_4_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_c42(1);
   bh56_w32_2_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_c42(2);
   Compressor_23_3_Freq800_uid289_uid340: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid340_In0_c41,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid340_In1_c41,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_copy341_c41);
   Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid340_Out0_copy341_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid342_In0_c41 <= "" & bh56_w32_0_c41 & bh56_w32_1_c41 & "0" & "0";
   Compressor_14_3_Freq800_uid271_bh56_uid342_In1_c41 <= "" & bh56_w33_0_c41;
   bh56_w32_3_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_c42(0);
   bh56_w33_1_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_c42(1);
   bh56_w34_1_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid342: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid342_In0_c41,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid342_In1_c41,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_copy343_c41);
   Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid342_Out0_copy343_c42; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid344_In0_c42 <= "" & bh56_w12_14_c42 & bh56_w12_15_c42 & bh56_w12_16_c42;
   bh56_w12_17_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid344_Out0_c42(0);
   bh56_w13_15_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid344_Out0_c42(1);
   Compressor_3_2_Freq800_uid277_uid344: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid344_In0_c42,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid344_Out0_copy345_c42);
   Compressor_3_2_Freq800_uid277_bh56_uid344_Out0_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid344_Out0_copy345_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid346_In0_c42 <= "" & bh56_w13_10_c42 & bh56_w13_11_c42 & bh56_w13_12_c42 & bh56_w13_13_c42;
   Compressor_14_3_Freq800_uid271_bh56_uid346_In1_c42 <= "" & bh56_w14_17_c42;
   bh56_w13_16_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid346_Out0_c42(0);
   bh56_w14_19_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid346_Out0_c42(1);
   bh56_w15_20_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid346_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid346: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid346_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid346_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid346_Out0_copy347_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid346_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid346_Out0_copy347_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid348_In0_c42 <= "" & bh56_w14_12_c42 & bh56_w14_13_c42 & bh56_w14_14_c42 & bh56_w14_15_c42 & bh56_w14_16_c42 & bh56_w14_18_c42;
   bh56_w14_20_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid348_Out0_c42(0);
   bh56_w15_21_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid348_Out0_c42(1);
   bh56_w16_21_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid348_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid348: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid348_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid348_Out0_copy349_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid348_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid348_Out0_copy349_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid350_In0_c42 <= "" & bh56_w15_19_c42 & bh56_w15_17_c42 & bh56_w15_14_c42 & bh56_w15_15_c42 & bh56_w15_16_c42 & bh56_w15_18_c42;
   bh56_w15_22_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid350_Out0_c42(0);
   bh56_w16_22_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid350_Out0_c42(1);
   bh56_w17_22_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid350_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid350: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid350_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid350_Out0_copy351_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid350_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid350_Out0_copy351_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid352_In0_c42 <= "" & bh56_w16_20_c42 & bh56_w16_18_c42 & bh56_w16_16_c42 & bh56_w16_15_c42 & bh56_w16_14_c42 & bh56_w16_17_c42;
   bh56_w16_23_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid352_Out0_c42(0);
   bh56_w17_23_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid352_Out0_c42(1);
   bh56_w18_21_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid352_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid352: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid352_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid352_Out0_copy353_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid352_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid352_Out0_copy353_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid354_In0_c42 <= "" & bh56_w17_20_c42 & bh56_w17_18_c42 & bh56_w17_16_c42 & bh56_w17_15_c42 & "0" & "0";
   bh56_w17_24_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid354_Out0_c42(0);
   bh56_w18_22_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid354_Out0_c42(1);
   bh56_w19_20_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid354_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid354: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid354_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid354_Out0_copy355_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid354_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid354_Out0_copy355_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid356_In0_c42 <= "" & bh56_w17_14_c42 & bh56_w17_17_c42 & bh56_w17_19_c42 & bh56_w17_21_c42;
   Compressor_14_3_Freq800_uid271_bh56_uid356_In1_c42 <= "" & bh56_w18_19_c42;
   bh56_w17_25_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid356_Out0_c42(0);
   bh56_w18_23_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid356_Out0_c42(1);
   bh56_w19_21_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid356_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid356: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid356_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid356_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid356_Out0_copy357_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid356_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid356_Out0_copy357_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid358_In0_c42 <= "" & bh56_w18_17_c42 & bh56_w18_14_c42 & bh56_w18_15_c42 & bh56_w18_16_c42 & bh56_w18_18_c42 & bh56_w18_20_c42;
   bh56_w18_24_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid358_Out0_c42(0);
   bh56_w19_22_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid358_Out0_c42(1);
   bh56_w20_18_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid358_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid358: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid358_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid358_Out0_copy359_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid358_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid358_Out0_copy359_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid360_In0_c42 <= "" & bh56_w19_18_c42 & bh56_w19_16_c42 & bh56_w19_15_c42 & bh56_w19_14_c42 & bh56_w19_13_c42 & "0";
   bh56_w19_23_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid360_Out0_c42(0);
   bh56_w20_19_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid360_Out0_c42(1);
   bh56_w21_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid360_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid360: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid360_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid360_Out0_copy361_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid360_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid360_Out0_copy361_c42; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid362_In0_c42 <= "" & bh56_w19_6_c42 & bh56_w19_17_c42 & bh56_w19_19_c42;
   bh56_w19_24_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid362_Out0_c42(0);
   bh56_w20_20_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid362_Out0_c42(1);
   Compressor_3_2_Freq800_uid277_uid362: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid362_In0_c42,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid362_Out0_copy363_c42);
   Compressor_3_2_Freq800_uid277_bh56_uid362_Out0_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid362_Out0_copy363_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid364_In0_c42 <= "" & bh56_w20_16_c42 & bh56_w20_15_c42 & bh56_w20_14_c42 & bh56_w20_13_c42 & bh56_w20_12_c42 & bh56_w20_17_c42;
   bh56_w20_21_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid364_Out0_c42(0);
   bh56_w21_18_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid364_Out0_c42(1);
   bh56_w22_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid364_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid364: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid364_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid364_Out0_copy365_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid364_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid364_Out0_copy365_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid366_In0_c42 <= "" & bh56_w21_10_c42 & bh56_w21_11_c42 & bh56_w21_12_c42 & bh56_w21_13_c42 & bh56_w21_14_c42 & bh56_w21_15_c42;
   bh56_w21_19_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid366_Out0_c42(0);
   bh56_w22_18_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid366_Out0_c42(1);
   bh56_w23_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid366_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid366: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid366_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid366_Out0_copy367_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid366_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid366_Out0_copy367_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid368_In0_c42 <= "" & bh56_w22_11_c42 & bh56_w22_12_c42 & bh56_w22_13_c42 & bh56_w22_14_c42 & bh56_w22_15_c42 & bh56_w22_16_c42;
   bh56_w22_19_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid368_Out0_c42(0);
   bh56_w23_16_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid368_Out0_c42(1);
   bh56_w24_15_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid368_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid368: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid368_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid368_Out0_copy369_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid368_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid368_Out0_copy369_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid370_In0_c42 <= "" & bh56_w23_9_c42 & bh56_w23_10_c42 & bh56_w23_11_c42 & bh56_w23_12_c42 & bh56_w23_13_c42 & bh56_w23_14_c42;
   bh56_w23_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid370_Out0_c42(0);
   bh56_w24_16_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid370_Out0_c42(1);
   bh56_w25_12_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid370_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid370: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid370_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid370_Out0_copy371_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid370_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid370_Out0_copy371_c42; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid265_bh56_uid372_In0_c42 <= "" & bh56_w24_9_c42 & bh56_w24_10_c42 & bh56_w24_11_c42 & bh56_w24_12_c42 & bh56_w24_13_c42 & bh56_w24_14_c42;
   bh56_w24_17_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid372_Out0_c42(0);
   bh56_w25_13_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid372_Out0_c42(1);
   bh56_w26_11_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid372_Out0_c42(2);
   Compressor_6_3_Freq800_uid265_uid372: Compressor_6_3_Freq800_uid265
      port map ( X0 => Compressor_6_3_Freq800_uid265_bh56_uid372_In0_c42,
                 R => Compressor_6_3_Freq800_uid265_bh56_uid372_Out0_copy373_c42);
   Compressor_6_3_Freq800_uid265_bh56_uid372_Out0_c42 <= Compressor_6_3_Freq800_uid265_bh56_uid372_Out0_copy373_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid374_In0_c42 <= "" & bh56_w25_8_c42 & bh56_w25_9_c42 & bh56_w25_10_c42 & bh56_w25_11_c42;
   Compressor_14_3_Freq800_uid271_bh56_uid374_In1_c41 <= "" & bh56_w26_6_c41;
   bh56_w25_14_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid374_Out0_c42(0);
   bh56_w26_12_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid374_Out0_c42(1);
   bh56_w27_9_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid374_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid374: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid374_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid374_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid374_Out0_copy375_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid374_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid374_Out0_copy375_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid376_In0_c42 <= "" & bh56_w26_7_c42 & bh56_w26_8_c42 & bh56_w26_9_c42 & bh56_w26_10_c42;
   Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c0 <= "" & "0";
   bh56_w26_13_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid376_Out0_c42(0);
   bh56_w27_10_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid376_Out0_c42(1);
   bh56_w28_9_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid376_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid376: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid376_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid376_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid376_Out0_copy377_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid376_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid376_Out0_copy377_c42; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid378_In0_c42 <= "" & bh56_w27_6_c42 & bh56_w27_7_c42 & bh56_w27_8_c42;
   bh56_w27_11_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid378_Out0_c42(0);
   bh56_w28_10_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid378_Out0_c42(1);
   Compressor_3_2_Freq800_uid277_uid378: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid378_In0_c42,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid378_Out0_copy379_c42);
   Compressor_3_2_Freq800_uid277_bh56_uid378_Out0_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid378_Out0_copy379_c42; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid380_In0_c42 <= "" & bh56_w28_6_c42 & bh56_w28_7_c42 & bh56_w28_8_c42;
   Compressor_23_3_Freq800_uid289_bh56_uid380_In1_c42 <= "" & bh56_w29_4_c42 & bh56_w29_5_c42;
   bh56_w28_11_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid380_Out0_c42(0);
   bh56_w29_7_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid380_Out0_c42(1);
   bh56_w30_7_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid380_Out0_c42(2);
   Compressor_23_3_Freq800_uid289_uid380: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid380_In0_c42,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid380_In1_c42,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid380_Out0_copy381_c42);
   Compressor_23_3_Freq800_uid289_bh56_uid380_Out0_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid380_Out0_copy381_c42; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid382_In0_c42 <= "" & bh56_w30_4_c42 & bh56_w30_5_c42 & bh56_w30_6_c42;
   Compressor_23_3_Freq800_uid289_bh56_uid382_In1_c42 <= "" & bh56_w31_2_c42 & bh56_w31_3_c42;
   bh56_w30_8_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid382_Out0_c42(0);
   bh56_w31_5_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid382_Out0_c42(1);
   bh56_w32_4_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid382_Out0_c42(2);
   Compressor_23_3_Freq800_uid289_uid382: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid382_In0_c42,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid382_In1_c42,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid382_Out0_copy383_c42);
   Compressor_23_3_Freq800_uid289_bh56_uid382_Out0_c42 <= Compressor_23_3_Freq800_uid289_bh56_uid382_Out0_copy383_c42; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid384_In0_c42 <= "" & bh56_w32_2_c42 & bh56_w32_3_c42 & "0" & "0";
   Compressor_14_3_Freq800_uid271_bh56_uid384_In1_c42 <= "" & bh56_w33_1_c42;
   bh56_w32_5_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid384_Out0_c42(0);
   bh56_w33_2_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid384_Out0_c42(1);
   bh56_w34_2_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid384_Out0_c42(2);
   Compressor_14_3_Freq800_uid271_uid384: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid384_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid384_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid384_Out0_copy385_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid384_Out0_c42 <= Compressor_14_3_Freq800_uid271_bh56_uid384_Out0_copy385_c42; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid386_In0_c42 <= "" & bh56_w34_0_c42 & bh56_w34_1_c42 & "0";
   bh56_w34_3_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid386_Out0_c42(0);
   Compressor_3_2_Freq800_uid277_uid386: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid386_In0_c42,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid386_Out0_copy387_c42);
   Compressor_3_2_Freq800_uid277_bh56_uid386_Out0_c42 <= Compressor_3_2_Freq800_uid277_bh56_uid386_Out0_copy387_c42; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid388_In0_c42 <= "" & bh56_w13_14_c42 & bh56_w13_15_c42 & bh56_w13_16_c42;
   Compressor_23_3_Freq800_uid289_bh56_uid388_In1_c42 <= "" & bh56_w14_19_c42 & bh56_w14_20_c42;
   bh56_w13_17_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_c43(0);
   bh56_w14_21_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_c43(1);
   bh56_w15_23_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid388: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid388_In0_c42,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid388_In1_c42,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_copy389_c42);
   Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid388_Out0_copy389_c43; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid390_In0_c42 <= "" & bh56_w15_20_c42 & bh56_w15_21_c42 & bh56_w15_22_c42;
   bh56_w15_24_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_c43(0);
   bh56_w16_24_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_c43(1);
   Compressor_3_2_Freq800_uid277_uid390: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid390_In0_c42,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_copy391_c42);
   Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid390_Out0_copy391_c43; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid392_In0_c42 <= "" & bh56_w16_19_c42 & bh56_w16_21_c42 & bh56_w16_22_c42 & bh56_w16_23_c42;
   Compressor_14_3_Freq800_uid271_bh56_uid392_In1_c42 <= "" & bh56_w17_22_c42;
   bh56_w16_25_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_c43(0);
   bh56_w17_26_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_c43(1);
   bh56_w18_25_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_c43(2);
   Compressor_14_3_Freq800_uid271_uid392: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid392_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid392_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_copy393_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid392_Out0_copy393_c43; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid394_In0_c42 <= "" & bh56_w17_23_c42 & bh56_w17_24_c42 & bh56_w17_25_c42;
   bh56_w17_27_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_c43(0);
   bh56_w18_26_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_c43(1);
   Compressor_3_2_Freq800_uid277_uid394: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid394_In0_c42,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_copy395_c42);
   Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid394_Out0_copy395_c43; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid396_In0_c42 <= "" & bh56_w18_21_c42 & bh56_w18_22_c42 & bh56_w18_23_c42 & bh56_w18_24_c42;
   Compressor_14_3_Freq800_uid271_bh56_uid396_In1_c42 <= "" & bh56_w19_20_c42;
   bh56_w18_27_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_c43(0);
   bh56_w19_25_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_c43(1);
   bh56_w20_22_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_c43(2);
   Compressor_14_3_Freq800_uid271_uid396: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid396_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid396_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_copy397_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid396_Out0_copy397_c43; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid398_In0_c42 <= "" & bh56_w19_21_c42 & bh56_w19_22_c42 & bh56_w19_23_c42 & bh56_w19_24_c42;
   Compressor_14_3_Freq800_uid271_bh56_uid398_In1_c42 <= "" & bh56_w20_18_c42;
   bh56_w19_26_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_c43(0);
   bh56_w20_23_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_c43(1);
   bh56_w21_20_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_c43(2);
   Compressor_14_3_Freq800_uid271_uid398: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid398_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid398_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_copy399_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid398_Out0_copy399_c43; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid400_In0_c42 <= "" & bh56_w20_19_c42 & bh56_w20_20_c42 & bh56_w20_21_c42;
   bh56_w20_24_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_c43(0);
   bh56_w21_21_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_c43(1);
   Compressor_3_2_Freq800_uid277_uid400: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid400_In0_c42,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_copy401_c42);
   Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid400_Out0_copy401_c43; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid402_In0_c42 <= "" & bh56_w21_16_c42 & bh56_w21_17_c42 & bh56_w21_18_c42 & bh56_w21_19_c42;
   Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c0 <= "" & "0";
   bh56_w21_22_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_c43(0);
   bh56_w22_20_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_c43(1);
   bh56_w23_18_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_c43(2);
   Compressor_14_3_Freq800_uid271_uid402: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid402_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid402_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_copy403_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid402_Out0_copy403_c43; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid404_In0_c42 <= "" & bh56_w22_17_c42 & bh56_w22_18_c42 & bh56_w22_19_c42;
   bh56_w22_21_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_c43(0);
   bh56_w23_19_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_c43(1);
   Compressor_3_2_Freq800_uid277_uid404: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid404_In0_c42,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_copy405_c42);
   Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid404_Out0_copy405_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid406_In0_c42 <= "" & bh56_w23_15_c42 & bh56_w23_16_c42 & bh56_w23_17_c42;
   Compressor_23_3_Freq800_uid289_bh56_uid406_In1_c42 <= "" & bh56_w24_15_c42 & bh56_w24_16_c42;
   bh56_w23_20_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_c43(0);
   bh56_w24_18_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_c43(1);
   bh56_w25_15_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid406: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid406_In0_c42,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid406_In1_c42,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_copy407_c42);
   Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid406_Out0_copy407_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid408_In0_c42 <= "" & bh56_w25_12_c42 & bh56_w25_13_c42 & bh56_w25_14_c42;
   Compressor_23_3_Freq800_uid289_bh56_uid408_In1_c42 <= "" & bh56_w26_11_c42 & bh56_w26_12_c42;
   bh56_w25_16_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_c43(0);
   bh56_w26_14_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_c43(1);
   bh56_w27_12_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid408: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid408_In0_c42,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid408_In1_c42,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_copy409_c42);
   Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid408_Out0_copy409_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid410_In0_c42 <= "" & bh56_w27_9_c42 & bh56_w27_10_c42 & bh56_w27_11_c42;
   Compressor_23_3_Freq800_uid289_bh56_uid410_In1_c42 <= "" & bh56_w28_9_c42 & bh56_w28_10_c42;
   bh56_w27_13_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_c43(0);
   bh56_w28_12_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_c43(1);
   bh56_w29_8_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid410: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid410_In0_c42,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid410_In1_c42,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_copy411_c42);
   Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid410_Out0_copy411_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid412_In0_c42 <= "" & bh56_w29_6_c42 & bh56_w29_7_c42 & "0";
   Compressor_23_3_Freq800_uid289_bh56_uid412_In1_c42 <= "" & bh56_w30_7_c42 & bh56_w30_8_c42;
   bh56_w29_9_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_c43(0);
   bh56_w30_9_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_c43(1);
   bh56_w31_6_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid412: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid412_In0_c42,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid412_In1_c42,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_copy413_c42);
   Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid412_Out0_copy413_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid414_In0_c42 <= "" & bh56_w31_4_c42 & bh56_w31_5_c42 & "0";
   Compressor_23_3_Freq800_uid289_bh56_uid414_In1_c42 <= "" & bh56_w32_4_c42 & bh56_w32_5_c42;
   bh56_w31_7_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_c43(0);
   bh56_w32_6_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_c43(1);
   bh56_w33_3_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid414: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid414_In0_c42,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid414_In1_c42,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_copy415_c42);
   Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid414_Out0_copy415_c43; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid416_In0_c42 <= "" & bh56_w34_2_c42 & bh56_w34_3_c42 & "0" & "0";
   Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c0 <= "" & "0";
   bh56_w34_4_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid416_Out0_c43(0);
   Compressor_14_3_Freq800_uid271_uid416: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid416_In0_c42,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid416_In1_c42,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid416_Out0_copy417_c42);
   Compressor_14_3_Freq800_uid271_bh56_uid416_Out0_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid416_Out0_copy417_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid418_In0_c43 <= "" & bh56_w15_23_c43 & bh56_w15_24_c43 & "0";
   Compressor_23_3_Freq800_uid289_bh56_uid418_In1_c43 <= "" & bh56_w16_24_c43 & bh56_w16_25_c43;
   bh56_w15_25_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid418_Out0_c43(0);
   bh56_w16_26_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid418_Out0_c43(1);
   bh56_w17_28_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid418_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid418: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid418_In0_c43,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid418_In1_c43,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid418_Out0_copy419_c43);
   Compressor_23_3_Freq800_uid289_bh56_uid418_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid418_Out0_copy419_c43; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid277_bh56_uid420_In0_c43 <= "" & bh56_w17_26_c43 & bh56_w17_27_c43 & "0";
   bh56_w17_29_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid420_Out0_c43(0);
   bh56_w18_28_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid420_Out0_c43(1);
   Compressor_3_2_Freq800_uid277_uid420: Compressor_3_2_Freq800_uid277
      port map ( X0 => Compressor_3_2_Freq800_uid277_bh56_uid420_In0_c43,
                 R => Compressor_3_2_Freq800_uid277_bh56_uid420_Out0_copy421_c43);
   Compressor_3_2_Freq800_uid277_bh56_uid420_Out0_c43 <= Compressor_3_2_Freq800_uid277_bh56_uid420_Out0_copy421_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid422_In0_c43 <= "" & bh56_w18_25_c43 & bh56_w18_26_c43 & bh56_w18_27_c43;
   Compressor_23_3_Freq800_uid289_bh56_uid422_In1_c43 <= "" & bh56_w19_25_c43 & bh56_w19_26_c43;
   bh56_w18_29_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid422_Out0_c43(0);
   bh56_w19_27_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid422_Out0_c43(1);
   bh56_w20_25_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid422_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid422: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid422_In0_c43,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid422_In1_c43,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid422_Out0_copy423_c43);
   Compressor_23_3_Freq800_uid289_bh56_uid422_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid422_Out0_copy423_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid424_In0_c43 <= "" & bh56_w20_22_c43 & bh56_w20_23_c43 & bh56_w20_24_c43;
   Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c0 <= "" & "0" & "0";
   bh56_w20_26_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid424_Out0_c43(0);
   bh56_w21_23_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid424_Out0_c43(1);
   bh56_w22_22_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid424_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid424: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid424_In0_c43,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid424_In1_c43,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid424_Out0_copy425_c43);
   Compressor_23_3_Freq800_uid289_bh56_uid424_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid424_Out0_copy425_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid426_In0_c43 <= "" & bh56_w21_20_c43 & bh56_w21_21_c43 & bh56_w21_22_c43;
   Compressor_23_3_Freq800_uid289_bh56_uid426_In1_c43 <= "" & bh56_w22_20_c43 & bh56_w22_21_c43;
   bh56_w21_24_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid426_Out0_c43(0);
   bh56_w22_23_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid426_Out0_c43(1);
   bh56_w23_21_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid426_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid426: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid426_In0_c43,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid426_In1_c43,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid426_Out0_copy427_c43);
   Compressor_23_3_Freq800_uid289_bh56_uid426_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid426_Out0_copy427_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid428_In0_c43 <= "" & bh56_w23_18_c43 & bh56_w23_19_c43 & bh56_w23_20_c43;
   Compressor_23_3_Freq800_uid289_bh56_uid428_In1_c43 <= "" & bh56_w24_17_c43 & bh56_w24_18_c43;
   bh56_w23_22_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid428_Out0_c43(0);
   bh56_w24_19_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid428_Out0_c43(1);
   bh56_w25_17_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid428_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid428: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid428_In0_c43,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid428_In1_c43,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid428_Out0_copy429_c43);
   Compressor_23_3_Freq800_uid289_bh56_uid428_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid428_Out0_copy429_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid430_In0_c43 <= "" & bh56_w25_15_c43 & bh56_w25_16_c43 & "0";
   Compressor_23_3_Freq800_uid289_bh56_uid430_In1_c43 <= "" & bh56_w26_13_c43 & bh56_w26_14_c43;
   bh56_w25_18_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid430_Out0_c43(0);
   bh56_w26_15_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid430_Out0_c43(1);
   bh56_w27_14_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid430_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid430: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid430_In0_c43,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid430_In1_c43,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid430_Out0_copy431_c43);
   Compressor_23_3_Freq800_uid289_bh56_uid430_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid430_Out0_copy431_c43; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid289_bh56_uid432_In0_c43 <= "" & bh56_w27_12_c43 & bh56_w27_13_c43 & "0";
   Compressor_23_3_Freq800_uid289_bh56_uid432_In1_c43 <= "" & bh56_w28_11_c43 & bh56_w28_12_c43;
   bh56_w27_15_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid432_Out0_c43(0);
   bh56_w28_13_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid432_Out0_c43(1);
   bh56_w29_10_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid432_Out0_c43(2);
   Compressor_23_3_Freq800_uid289_uid432: Compressor_23_3_Freq800_uid289
      port map ( X0 => Compressor_23_3_Freq800_uid289_bh56_uid432_In0_c43,
                 X1 => Compressor_23_3_Freq800_uid289_bh56_uid432_In1_c43,
                 R => Compressor_23_3_Freq800_uid289_bh56_uid432_Out0_copy433_c43);
   Compressor_23_3_Freq800_uid289_bh56_uid432_Out0_c43 <= Compressor_23_3_Freq800_uid289_bh56_uid432_Out0_copy433_c43; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid434_In0_c43 <= "" & bh56_w29_8_c43 & bh56_w29_9_c43 & "0" & "0";
   Compressor_14_3_Freq800_uid271_bh56_uid434_In1_c43 <= "" & bh56_w30_9_c43;
   bh56_w29_11_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid434_Out0_c43(0);
   bh56_w30_10_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid434_Out0_c43(1);
   bh56_w31_8_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid434_Out0_c43(2);
   Compressor_14_3_Freq800_uid271_uid434: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid434_In0_c43,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid434_In1_c43,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid434_Out0_copy435_c43);
   Compressor_14_3_Freq800_uid271_bh56_uid434_Out0_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid434_Out0_copy435_c43; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid436_In0_c43 <= "" & bh56_w31_6_c43 & bh56_w31_7_c43 & "0" & "0";
   Compressor_14_3_Freq800_uid271_bh56_uid436_In1_c43 <= "" & bh56_w32_6_c43;
   bh56_w31_9_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid436_Out0_c43(0);
   bh56_w32_7_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid436_Out0_c43(1);
   bh56_w33_4_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid436_Out0_c43(2);
   Compressor_14_3_Freq800_uid271_uid436: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid436_In0_c43,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid436_In1_c43,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid436_Out0_copy437_c43);
   Compressor_14_3_Freq800_uid271_bh56_uid436_Out0_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid436_Out0_copy437_c43; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid271_bh56_uid438_In0_c43 <= "" & bh56_w33_2_c43 & bh56_w33_3_c43 & "0" & "0";
   Compressor_14_3_Freq800_uid271_bh56_uid438_In1_c43 <= "" & bh56_w34_4_c43;
   bh56_w33_5_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid438_Out0_c43(0);
   bh56_w34_5_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid438_Out0_c43(1);
   Compressor_14_3_Freq800_uid271_uid438: Compressor_14_3_Freq800_uid271
      port map ( X0 => Compressor_14_3_Freq800_uid271_bh56_uid438_In0_c43,
                 X1 => Compressor_14_3_Freq800_uid271_bh56_uid438_In1_c43,
                 R => Compressor_14_3_Freq800_uid271_bh56_uid438_Out0_copy439_c43);
   Compressor_14_3_Freq800_uid271_bh56_uid438_Out0_c43 <= Compressor_14_3_Freq800_uid271_bh56_uid438_Out0_copy439_c43; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh56_16_c43 <= bh56_w16_26_c43 & bh56_w15_25_c43 & bh56_w14_21_c43 & bh56_w13_17_c43 & bh56_w12_17_c43 & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0" & "0";

   bitheapFinalAdd_bh56_In0_c43 <= "0" & bh56_w34_5_c43 & bh56_w33_4_c43 & bh56_w32_7_c43 & bh56_w31_8_c43 & bh56_w30_10_c43 & bh56_w29_10_c43 & bh56_w28_13_c43 & bh56_w27_14_c43 & bh56_w26_15_c43 & bh56_w25_17_c43 & bh56_w24_19_c43 & bh56_w23_21_c43 & bh56_w22_22_c43 & bh56_w21_23_c43 & bh56_w20_25_c43 & bh56_w19_27_c43 & bh56_w18_28_c43 & bh56_w17_28_c43;
   bitheapFinalAdd_bh56_In1_c43 <= "0" & "0" & bh56_w33_5_c43 & "0" & bh56_w31_9_c43 & "0" & bh56_w29_11_c43 & "0" & bh56_w27_15_c43 & "0" & bh56_w25_18_c43 & "0" & bh56_w23_22_c43 & bh56_w22_23_c43 & bh56_w21_24_c43 & bh56_w20_26_c43 & "0" & bh56_w18_29_c43 & bh56_w17_29_c43;
   bitheapFinalAdd_bh56_Cin_c0 <= '0';

   bitheapFinalAdd_bh56: IntAdder_19_Freq800_uid441
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 ce_36=> ce_36,
                 ce_37=> ce_37,
                 ce_38=> ce_38,
                 ce_39=> ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 ce_42=> ce_42,
                 ce_43=> ce_43,
                 ce_44=> ce_44,
                 ce_45=> ce_45,
                 ce_46=> ce_46,
                 ce_47=> ce_47,
                 ce_48=> ce_48,
                 ce_49=> ce_49,
                 ce_50=> ce_50,
                 Cin => bitheapFinalAdd_bh56_Cin_c0,
                 X => bitheapFinalAdd_bh56_In0_c43,
                 Y => bitheapFinalAdd_bh56_In1_c43,
                 R => bitheapFinalAdd_bh56_Out_c50);
   bitheapResult_bh56_c50 <= bitheapFinalAdd_bh56_Out_c50(17 downto 0) & tmp_bitheapResult_bh56_16_c50;
   R <= bitheapResult_bh56_c50(34 downto 16);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_28_Freq800_uid444
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 61 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_28_Freq800_uid444 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56, ce_57, ce_58, ce_59, ce_60, ce_61 : in std_logic;
          X : in  std_logic_vector(27 downto 0);
          Y : in  std_logic_vector(27 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of IntAdder_28_Freq800_uid444 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3, Cin_0_c4, Cin_0_c5, Cin_0_c6, Cin_0_c7, Cin_0_c8, Cin_0_c9, Cin_0_c10, Cin_0_c11, Cin_0_c12, Cin_0_c13, Cin_0_c14, Cin_0_c15, Cin_0_c16, Cin_0_c17, Cin_0_c18, Cin_0_c19, Cin_0_c20, Cin_0_c21, Cin_0_c22, Cin_0_c23, Cin_0_c24, Cin_0_c25, Cin_0_c26, Cin_0_c27, Cin_0_c28, Cin_0_c29, Cin_0_c30, Cin_0_c31, Cin_0_c32, Cin_0_c33, Cin_0_c34, Cin_0_c35, Cin_0_c36, Cin_0_c37, Cin_0_c38, Cin_0_c39, Cin_0_c40, Cin_0_c41, Cin_0_c42, Cin_0_c43, Cin_0_c44, Cin_0_c45, Cin_0_c46, Cin_0_c47, Cin_0_c48, Cin_0_c49, Cin_0_c50, Cin_0_c51 :  std_logic;
signal X_0_c35, X_0_c36, X_0_c37, X_0_c38, X_0_c39, X_0_c40, X_0_c41, X_0_c42, X_0_c43, X_0_c44, X_0_c45, X_0_c46, X_0_c47, X_0_c48, X_0_c49, X_0_c50, X_0_c51 :  std_logic_vector(3 downto 0);
signal Y_0_c50, Y_0_c51 :  std_logic_vector(3 downto 0);
signal S_0_c51 :  std_logic_vector(3 downto 0);
signal R_0_c51, R_0_c52, R_0_c53, R_0_c54, R_0_c55, R_0_c56, R_0_c57, R_0_c58, R_0_c59, R_0_c60, R_0_c61 :  std_logic_vector(2 downto 0);
signal Cin_1_c51, Cin_1_c52 :  std_logic;
signal X_1_c35, X_1_c36, X_1_c37, X_1_c38, X_1_c39, X_1_c40, X_1_c41, X_1_c42, X_1_c43, X_1_c44, X_1_c45, X_1_c46, X_1_c47, X_1_c48, X_1_c49, X_1_c50, X_1_c51, X_1_c52 :  std_logic_vector(3 downto 0);
signal Y_1_c50, Y_1_c51, Y_1_c52 :  std_logic_vector(3 downto 0);
signal S_1_c52 :  std_logic_vector(3 downto 0);
signal R_1_c52, R_1_c53, R_1_c54, R_1_c55, R_1_c56, R_1_c57, R_1_c58, R_1_c59, R_1_c60, R_1_c61 :  std_logic_vector(2 downto 0);
signal Cin_2_c52, Cin_2_c53 :  std_logic;
signal X_2_c35, X_2_c36, X_2_c37, X_2_c38, X_2_c39, X_2_c40, X_2_c41, X_2_c42, X_2_c43, X_2_c44, X_2_c45, X_2_c46, X_2_c47, X_2_c48, X_2_c49, X_2_c50, X_2_c51, X_2_c52, X_2_c53 :  std_logic_vector(3 downto 0);
signal Y_2_c50, Y_2_c51, Y_2_c52, Y_2_c53 :  std_logic_vector(3 downto 0);
signal S_2_c53 :  std_logic_vector(3 downto 0);
signal R_2_c53, R_2_c54, R_2_c55, R_2_c56, R_2_c57, R_2_c58, R_2_c59, R_2_c60, R_2_c61 :  std_logic_vector(2 downto 0);
signal Cin_3_c53, Cin_3_c54, Cin_3_c55 :  std_logic;
signal X_3_c35, X_3_c36, X_3_c37, X_3_c38, X_3_c39, X_3_c40, X_3_c41, X_3_c42, X_3_c43, X_3_c44, X_3_c45, X_3_c46, X_3_c47, X_3_c48, X_3_c49, X_3_c50, X_3_c51, X_3_c52, X_3_c53, X_3_c54, X_3_c55 :  std_logic_vector(3 downto 0);
signal Y_3_c50, Y_3_c51, Y_3_c52, Y_3_c53, Y_3_c54, Y_3_c55 :  std_logic_vector(3 downto 0);
signal S_3_c55 :  std_logic_vector(3 downto 0);
signal R_3_c55, R_3_c56, R_3_c57, R_3_c58, R_3_c59, R_3_c60, R_3_c61 :  std_logic_vector(2 downto 0);
signal Cin_4_c55, Cin_4_c56 :  std_logic;
signal X_4_c35, X_4_c36, X_4_c37, X_4_c38, X_4_c39, X_4_c40, X_4_c41, X_4_c42, X_4_c43, X_4_c44, X_4_c45, X_4_c46, X_4_c47, X_4_c48, X_4_c49, X_4_c50, X_4_c51, X_4_c52, X_4_c53, X_4_c54, X_4_c55, X_4_c56 :  std_logic_vector(3 downto 0);
signal Y_4_c50, Y_4_c51, Y_4_c52, Y_4_c53, Y_4_c54, Y_4_c55, Y_4_c56 :  std_logic_vector(3 downto 0);
signal S_4_c56 :  std_logic_vector(3 downto 0);
signal R_4_c56, R_4_c57, R_4_c58, R_4_c59, R_4_c60, R_4_c61 :  std_logic_vector(2 downto 0);
signal Cin_5_c56, Cin_5_c57 :  std_logic;
signal X_5_c35, X_5_c36, X_5_c37, X_5_c38, X_5_c39, X_5_c40, X_5_c41, X_5_c42, X_5_c43, X_5_c44, X_5_c45, X_5_c46, X_5_c47, X_5_c48, X_5_c49, X_5_c50, X_5_c51, X_5_c52, X_5_c53, X_5_c54, X_5_c55, X_5_c56, X_5_c57 :  std_logic_vector(3 downto 0);
signal Y_5_c50, Y_5_c51, Y_5_c52, Y_5_c53, Y_5_c54, Y_5_c55, Y_5_c56, Y_5_c57 :  std_logic_vector(3 downto 0);
signal S_5_c57 :  std_logic_vector(3 downto 0);
signal R_5_c57, R_5_c58, R_5_c59, R_5_c60, R_5_c61 :  std_logic_vector(2 downto 0);
signal Cin_6_c57, Cin_6_c58 :  std_logic;
signal X_6_c35, X_6_c36, X_6_c37, X_6_c38, X_6_c39, X_6_c40, X_6_c41, X_6_c42, X_6_c43, X_6_c44, X_6_c45, X_6_c46, X_6_c47, X_6_c48, X_6_c49, X_6_c50, X_6_c51, X_6_c52, X_6_c53, X_6_c54, X_6_c55, X_6_c56, X_6_c57, X_6_c58 :  std_logic_vector(3 downto 0);
signal Y_6_c50, Y_6_c51, Y_6_c52, Y_6_c53, Y_6_c54, Y_6_c55, Y_6_c56, Y_6_c57, Y_6_c58 :  std_logic_vector(3 downto 0);
signal S_6_c58 :  std_logic_vector(3 downto 0);
signal R_6_c58, R_6_c59, R_6_c60, R_6_c61 :  std_logic_vector(2 downto 0);
signal Cin_7_c58, Cin_7_c59 :  std_logic;
signal X_7_c35, X_7_c36, X_7_c37, X_7_c38, X_7_c39, X_7_c40, X_7_c41, X_7_c42, X_7_c43, X_7_c44, X_7_c45, X_7_c46, X_7_c47, X_7_c48, X_7_c49, X_7_c50, X_7_c51, X_7_c52, X_7_c53, X_7_c54, X_7_c55, X_7_c56, X_7_c57, X_7_c58, X_7_c59 :  std_logic_vector(3 downto 0);
signal Y_7_c50, Y_7_c51, Y_7_c52, Y_7_c53, Y_7_c54, Y_7_c55, Y_7_c56, Y_7_c57, Y_7_c58, Y_7_c59 :  std_logic_vector(3 downto 0);
signal S_7_c59 :  std_logic_vector(3 downto 0);
signal R_7_c59, R_7_c60, R_7_c61 :  std_logic_vector(2 downto 0);
signal Cin_8_c59, Cin_8_c60 :  std_logic;
signal X_8_c35, X_8_c36, X_8_c37, X_8_c38, X_8_c39, X_8_c40, X_8_c41, X_8_c42, X_8_c43, X_8_c44, X_8_c45, X_8_c46, X_8_c47, X_8_c48, X_8_c49, X_8_c50, X_8_c51, X_8_c52, X_8_c53, X_8_c54, X_8_c55, X_8_c56, X_8_c57, X_8_c58, X_8_c59, X_8_c60 :  std_logic_vector(3 downto 0);
signal Y_8_c50, Y_8_c51, Y_8_c52, Y_8_c53, Y_8_c54, Y_8_c55, Y_8_c56, Y_8_c57, Y_8_c58, Y_8_c59, Y_8_c60 :  std_logic_vector(3 downto 0);
signal S_8_c60 :  std_logic_vector(3 downto 0);
signal R_8_c60, R_8_c61 :  std_logic_vector(2 downto 0);
signal Cin_9_c60, Cin_9_c61 :  std_logic;
signal X_9_c35, X_9_c36, X_9_c37, X_9_c38, X_9_c39, X_9_c40, X_9_c41, X_9_c42, X_9_c43, X_9_c44, X_9_c45, X_9_c46, X_9_c47, X_9_c48, X_9_c49, X_9_c50, X_9_c51, X_9_c52, X_9_c53, X_9_c54, X_9_c55, X_9_c56, X_9_c57, X_9_c58, X_9_c59, X_9_c60, X_9_c61 :  std_logic_vector(1 downto 0);
signal Y_9_c50, Y_9_c51, Y_9_c52, Y_9_c53, Y_9_c54, Y_9_c55, Y_9_c56, Y_9_c57, Y_9_c58, Y_9_c59, Y_9_c60, Y_9_c61 :  std_logic_vector(1 downto 0);
signal S_9_c61 :  std_logic_vector(1 downto 0);
signal R_9_c61 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
            end if;
            if ce_4 = '1' then
               Cin_0_c4 <= Cin_0_c3;
            end if;
            if ce_5 = '1' then
               Cin_0_c5 <= Cin_0_c4;
            end if;
            if ce_6 = '1' then
               Cin_0_c6 <= Cin_0_c5;
            end if;
            if ce_7 = '1' then
               Cin_0_c7 <= Cin_0_c6;
            end if;
            if ce_8 = '1' then
               Cin_0_c8 <= Cin_0_c7;
            end if;
            if ce_9 = '1' then
               Cin_0_c9 <= Cin_0_c8;
            end if;
            if ce_10 = '1' then
               Cin_0_c10 <= Cin_0_c9;
            end if;
            if ce_11 = '1' then
               Cin_0_c11 <= Cin_0_c10;
            end if;
            if ce_12 = '1' then
               Cin_0_c12 <= Cin_0_c11;
            end if;
            if ce_13 = '1' then
               Cin_0_c13 <= Cin_0_c12;
            end if;
            if ce_14 = '1' then
               Cin_0_c14 <= Cin_0_c13;
            end if;
            if ce_15 = '1' then
               Cin_0_c15 <= Cin_0_c14;
            end if;
            if ce_16 = '1' then
               Cin_0_c16 <= Cin_0_c15;
            end if;
            if ce_17 = '1' then
               Cin_0_c17 <= Cin_0_c16;
            end if;
            if ce_18 = '1' then
               Cin_0_c18 <= Cin_0_c17;
            end if;
            if ce_19 = '1' then
               Cin_0_c19 <= Cin_0_c18;
            end if;
            if ce_20 = '1' then
               Cin_0_c20 <= Cin_0_c19;
            end if;
            if ce_21 = '1' then
               Cin_0_c21 <= Cin_0_c20;
            end if;
            if ce_22 = '1' then
               Cin_0_c22 <= Cin_0_c21;
            end if;
            if ce_23 = '1' then
               Cin_0_c23 <= Cin_0_c22;
            end if;
            if ce_24 = '1' then
               Cin_0_c24 <= Cin_0_c23;
            end if;
            if ce_25 = '1' then
               Cin_0_c25 <= Cin_0_c24;
            end if;
            if ce_26 = '1' then
               Cin_0_c26 <= Cin_0_c25;
            end if;
            if ce_27 = '1' then
               Cin_0_c27 <= Cin_0_c26;
            end if;
            if ce_28 = '1' then
               Cin_0_c28 <= Cin_0_c27;
            end if;
            if ce_29 = '1' then
               Cin_0_c29 <= Cin_0_c28;
            end if;
            if ce_30 = '1' then
               Cin_0_c30 <= Cin_0_c29;
            end if;
            if ce_31 = '1' then
               Cin_0_c31 <= Cin_0_c30;
            end if;
            if ce_32 = '1' then
               Cin_0_c32 <= Cin_0_c31;
            end if;
            if ce_33 = '1' then
               Cin_0_c33 <= Cin_0_c32;
            end if;
            if ce_34 = '1' then
               Cin_0_c34 <= Cin_0_c33;
            end if;
            if ce_35 = '1' then
               Cin_0_c35 <= Cin_0_c34;
            end if;
            if ce_36 = '1' then
               Cin_0_c36 <= Cin_0_c35;
               X_0_c36 <= X_0_c35;
               X_1_c36 <= X_1_c35;
               X_2_c36 <= X_2_c35;
               X_3_c36 <= X_3_c35;
               X_4_c36 <= X_4_c35;
               X_5_c36 <= X_5_c35;
               X_6_c36 <= X_6_c35;
               X_7_c36 <= X_7_c35;
               X_8_c36 <= X_8_c35;
               X_9_c36 <= X_9_c35;
            end if;
            if ce_37 = '1' then
               Cin_0_c37 <= Cin_0_c36;
               X_0_c37 <= X_0_c36;
               X_1_c37 <= X_1_c36;
               X_2_c37 <= X_2_c36;
               X_3_c37 <= X_3_c36;
               X_4_c37 <= X_4_c36;
               X_5_c37 <= X_5_c36;
               X_6_c37 <= X_6_c36;
               X_7_c37 <= X_7_c36;
               X_8_c37 <= X_8_c36;
               X_9_c37 <= X_9_c36;
            end if;
            if ce_38 = '1' then
               Cin_0_c38 <= Cin_0_c37;
               X_0_c38 <= X_0_c37;
               X_1_c38 <= X_1_c37;
               X_2_c38 <= X_2_c37;
               X_3_c38 <= X_3_c37;
               X_4_c38 <= X_4_c37;
               X_5_c38 <= X_5_c37;
               X_6_c38 <= X_6_c37;
               X_7_c38 <= X_7_c37;
               X_8_c38 <= X_8_c37;
               X_9_c38 <= X_9_c37;
            end if;
            if ce_39 = '1' then
               Cin_0_c39 <= Cin_0_c38;
               X_0_c39 <= X_0_c38;
               X_1_c39 <= X_1_c38;
               X_2_c39 <= X_2_c38;
               X_3_c39 <= X_3_c38;
               X_4_c39 <= X_4_c38;
               X_5_c39 <= X_5_c38;
               X_6_c39 <= X_6_c38;
               X_7_c39 <= X_7_c38;
               X_8_c39 <= X_8_c38;
               X_9_c39 <= X_9_c38;
            end if;
            if ce_40 = '1' then
               Cin_0_c40 <= Cin_0_c39;
               X_0_c40 <= X_0_c39;
               X_1_c40 <= X_1_c39;
               X_2_c40 <= X_2_c39;
               X_3_c40 <= X_3_c39;
               X_4_c40 <= X_4_c39;
               X_5_c40 <= X_5_c39;
               X_6_c40 <= X_6_c39;
               X_7_c40 <= X_7_c39;
               X_8_c40 <= X_8_c39;
               X_9_c40 <= X_9_c39;
            end if;
            if ce_41 = '1' then
               Cin_0_c41 <= Cin_0_c40;
               X_0_c41 <= X_0_c40;
               X_1_c41 <= X_1_c40;
               X_2_c41 <= X_2_c40;
               X_3_c41 <= X_3_c40;
               X_4_c41 <= X_4_c40;
               X_5_c41 <= X_5_c40;
               X_6_c41 <= X_6_c40;
               X_7_c41 <= X_7_c40;
               X_8_c41 <= X_8_c40;
               X_9_c41 <= X_9_c40;
            end if;
            if ce_42 = '1' then
               Cin_0_c42 <= Cin_0_c41;
               X_0_c42 <= X_0_c41;
               X_1_c42 <= X_1_c41;
               X_2_c42 <= X_2_c41;
               X_3_c42 <= X_3_c41;
               X_4_c42 <= X_4_c41;
               X_5_c42 <= X_5_c41;
               X_6_c42 <= X_6_c41;
               X_7_c42 <= X_7_c41;
               X_8_c42 <= X_8_c41;
               X_9_c42 <= X_9_c41;
            end if;
            if ce_43 = '1' then
               Cin_0_c43 <= Cin_0_c42;
               X_0_c43 <= X_0_c42;
               X_1_c43 <= X_1_c42;
               X_2_c43 <= X_2_c42;
               X_3_c43 <= X_3_c42;
               X_4_c43 <= X_4_c42;
               X_5_c43 <= X_5_c42;
               X_6_c43 <= X_6_c42;
               X_7_c43 <= X_7_c42;
               X_8_c43 <= X_8_c42;
               X_9_c43 <= X_9_c42;
            end if;
            if ce_44 = '1' then
               Cin_0_c44 <= Cin_0_c43;
               X_0_c44 <= X_0_c43;
               X_1_c44 <= X_1_c43;
               X_2_c44 <= X_2_c43;
               X_3_c44 <= X_3_c43;
               X_4_c44 <= X_4_c43;
               X_5_c44 <= X_5_c43;
               X_6_c44 <= X_6_c43;
               X_7_c44 <= X_7_c43;
               X_8_c44 <= X_8_c43;
               X_9_c44 <= X_9_c43;
            end if;
            if ce_45 = '1' then
               Cin_0_c45 <= Cin_0_c44;
               X_0_c45 <= X_0_c44;
               X_1_c45 <= X_1_c44;
               X_2_c45 <= X_2_c44;
               X_3_c45 <= X_3_c44;
               X_4_c45 <= X_4_c44;
               X_5_c45 <= X_5_c44;
               X_6_c45 <= X_6_c44;
               X_7_c45 <= X_7_c44;
               X_8_c45 <= X_8_c44;
               X_9_c45 <= X_9_c44;
            end if;
            if ce_46 = '1' then
               Cin_0_c46 <= Cin_0_c45;
               X_0_c46 <= X_0_c45;
               X_1_c46 <= X_1_c45;
               X_2_c46 <= X_2_c45;
               X_3_c46 <= X_3_c45;
               X_4_c46 <= X_4_c45;
               X_5_c46 <= X_5_c45;
               X_6_c46 <= X_6_c45;
               X_7_c46 <= X_7_c45;
               X_8_c46 <= X_8_c45;
               X_9_c46 <= X_9_c45;
            end if;
            if ce_47 = '1' then
               Cin_0_c47 <= Cin_0_c46;
               X_0_c47 <= X_0_c46;
               X_1_c47 <= X_1_c46;
               X_2_c47 <= X_2_c46;
               X_3_c47 <= X_3_c46;
               X_4_c47 <= X_4_c46;
               X_5_c47 <= X_5_c46;
               X_6_c47 <= X_6_c46;
               X_7_c47 <= X_7_c46;
               X_8_c47 <= X_8_c46;
               X_9_c47 <= X_9_c46;
            end if;
            if ce_48 = '1' then
               Cin_0_c48 <= Cin_0_c47;
               X_0_c48 <= X_0_c47;
               X_1_c48 <= X_1_c47;
               X_2_c48 <= X_2_c47;
               X_3_c48 <= X_3_c47;
               X_4_c48 <= X_4_c47;
               X_5_c48 <= X_5_c47;
               X_6_c48 <= X_6_c47;
               X_7_c48 <= X_7_c47;
               X_8_c48 <= X_8_c47;
               X_9_c48 <= X_9_c47;
            end if;
            if ce_49 = '1' then
               Cin_0_c49 <= Cin_0_c48;
               X_0_c49 <= X_0_c48;
               X_1_c49 <= X_1_c48;
               X_2_c49 <= X_2_c48;
               X_3_c49 <= X_3_c48;
               X_4_c49 <= X_4_c48;
               X_5_c49 <= X_5_c48;
               X_6_c49 <= X_6_c48;
               X_7_c49 <= X_7_c48;
               X_8_c49 <= X_8_c48;
               X_9_c49 <= X_9_c48;
            end if;
            if ce_50 = '1' then
               Cin_0_c50 <= Cin_0_c49;
               X_0_c50 <= X_0_c49;
               X_1_c50 <= X_1_c49;
               X_2_c50 <= X_2_c49;
               X_3_c50 <= X_3_c49;
               X_4_c50 <= X_4_c49;
               X_5_c50 <= X_5_c49;
               X_6_c50 <= X_6_c49;
               X_7_c50 <= X_7_c49;
               X_8_c50 <= X_8_c49;
               X_9_c50 <= X_9_c49;
            end if;
            if ce_51 = '1' then
               Cin_0_c51 <= Cin_0_c50;
               X_0_c51 <= X_0_c50;
               Y_0_c51 <= Y_0_c50;
               X_1_c51 <= X_1_c50;
               Y_1_c51 <= Y_1_c50;
               X_2_c51 <= X_2_c50;
               Y_2_c51 <= Y_2_c50;
               X_3_c51 <= X_3_c50;
               Y_3_c51 <= Y_3_c50;
               X_4_c51 <= X_4_c50;
               Y_4_c51 <= Y_4_c50;
               X_5_c51 <= X_5_c50;
               Y_5_c51 <= Y_5_c50;
               X_6_c51 <= X_6_c50;
               Y_6_c51 <= Y_6_c50;
               X_7_c51 <= X_7_c50;
               Y_7_c51 <= Y_7_c50;
               X_8_c51 <= X_8_c50;
               Y_8_c51 <= Y_8_c50;
               X_9_c51 <= X_9_c50;
               Y_9_c51 <= Y_9_c50;
            end if;
            if ce_52 = '1' then
               R_0_c52 <= R_0_c51;
               Cin_1_c52 <= Cin_1_c51;
               X_1_c52 <= X_1_c51;
               Y_1_c52 <= Y_1_c51;
               X_2_c52 <= X_2_c51;
               Y_2_c52 <= Y_2_c51;
               X_3_c52 <= X_3_c51;
               Y_3_c52 <= Y_3_c51;
               X_4_c52 <= X_4_c51;
               Y_4_c52 <= Y_4_c51;
               X_5_c52 <= X_5_c51;
               Y_5_c52 <= Y_5_c51;
               X_6_c52 <= X_6_c51;
               Y_6_c52 <= Y_6_c51;
               X_7_c52 <= X_7_c51;
               Y_7_c52 <= Y_7_c51;
               X_8_c52 <= X_8_c51;
               Y_8_c52 <= Y_8_c51;
               X_9_c52 <= X_9_c51;
               Y_9_c52 <= Y_9_c51;
            end if;
            if ce_53 = '1' then
               R_0_c53 <= R_0_c52;
               R_1_c53 <= R_1_c52;
               Cin_2_c53 <= Cin_2_c52;
               X_2_c53 <= X_2_c52;
               Y_2_c53 <= Y_2_c52;
               X_3_c53 <= X_3_c52;
               Y_3_c53 <= Y_3_c52;
               X_4_c53 <= X_4_c52;
               Y_4_c53 <= Y_4_c52;
               X_5_c53 <= X_5_c52;
               Y_5_c53 <= Y_5_c52;
               X_6_c53 <= X_6_c52;
               Y_6_c53 <= Y_6_c52;
               X_7_c53 <= X_7_c52;
               Y_7_c53 <= Y_7_c52;
               X_8_c53 <= X_8_c52;
               Y_8_c53 <= Y_8_c52;
               X_9_c53 <= X_9_c52;
               Y_9_c53 <= Y_9_c52;
            end if;
            if ce_54 = '1' then
               R_0_c54 <= R_0_c53;
               R_1_c54 <= R_1_c53;
               R_2_c54 <= R_2_c53;
               Cin_3_c54 <= Cin_3_c53;
               X_3_c54 <= X_3_c53;
               Y_3_c54 <= Y_3_c53;
               X_4_c54 <= X_4_c53;
               Y_4_c54 <= Y_4_c53;
               X_5_c54 <= X_5_c53;
               Y_5_c54 <= Y_5_c53;
               X_6_c54 <= X_6_c53;
               Y_6_c54 <= Y_6_c53;
               X_7_c54 <= X_7_c53;
               Y_7_c54 <= Y_7_c53;
               X_8_c54 <= X_8_c53;
               Y_8_c54 <= Y_8_c53;
               X_9_c54 <= X_9_c53;
               Y_9_c54 <= Y_9_c53;
            end if;
            if ce_55 = '1' then
               R_0_c55 <= R_0_c54;
               R_1_c55 <= R_1_c54;
               R_2_c55 <= R_2_c54;
               Cin_3_c55 <= Cin_3_c54;
               X_3_c55 <= X_3_c54;
               Y_3_c55 <= Y_3_c54;
               X_4_c55 <= X_4_c54;
               Y_4_c55 <= Y_4_c54;
               X_5_c55 <= X_5_c54;
               Y_5_c55 <= Y_5_c54;
               X_6_c55 <= X_6_c54;
               Y_6_c55 <= Y_6_c54;
               X_7_c55 <= X_7_c54;
               Y_7_c55 <= Y_7_c54;
               X_8_c55 <= X_8_c54;
               Y_8_c55 <= Y_8_c54;
               X_9_c55 <= X_9_c54;
               Y_9_c55 <= Y_9_c54;
            end if;
            if ce_56 = '1' then
               R_0_c56 <= R_0_c55;
               R_1_c56 <= R_1_c55;
               R_2_c56 <= R_2_c55;
               R_3_c56 <= R_3_c55;
               Cin_4_c56 <= Cin_4_c55;
               X_4_c56 <= X_4_c55;
               Y_4_c56 <= Y_4_c55;
               X_5_c56 <= X_5_c55;
               Y_5_c56 <= Y_5_c55;
               X_6_c56 <= X_6_c55;
               Y_6_c56 <= Y_6_c55;
               X_7_c56 <= X_7_c55;
               Y_7_c56 <= Y_7_c55;
               X_8_c56 <= X_8_c55;
               Y_8_c56 <= Y_8_c55;
               X_9_c56 <= X_9_c55;
               Y_9_c56 <= Y_9_c55;
            end if;
            if ce_57 = '1' then
               R_0_c57 <= R_0_c56;
               R_1_c57 <= R_1_c56;
               R_2_c57 <= R_2_c56;
               R_3_c57 <= R_3_c56;
               R_4_c57 <= R_4_c56;
               Cin_5_c57 <= Cin_5_c56;
               X_5_c57 <= X_5_c56;
               Y_5_c57 <= Y_5_c56;
               X_6_c57 <= X_6_c56;
               Y_6_c57 <= Y_6_c56;
               X_7_c57 <= X_7_c56;
               Y_7_c57 <= Y_7_c56;
               X_8_c57 <= X_8_c56;
               Y_8_c57 <= Y_8_c56;
               X_9_c57 <= X_9_c56;
               Y_9_c57 <= Y_9_c56;
            end if;
            if ce_58 = '1' then
               R_0_c58 <= R_0_c57;
               R_1_c58 <= R_1_c57;
               R_2_c58 <= R_2_c57;
               R_3_c58 <= R_3_c57;
               R_4_c58 <= R_4_c57;
               R_5_c58 <= R_5_c57;
               Cin_6_c58 <= Cin_6_c57;
               X_6_c58 <= X_6_c57;
               Y_6_c58 <= Y_6_c57;
               X_7_c58 <= X_7_c57;
               Y_7_c58 <= Y_7_c57;
               X_8_c58 <= X_8_c57;
               Y_8_c58 <= Y_8_c57;
               X_9_c58 <= X_9_c57;
               Y_9_c58 <= Y_9_c57;
            end if;
            if ce_59 = '1' then
               R_0_c59 <= R_0_c58;
               R_1_c59 <= R_1_c58;
               R_2_c59 <= R_2_c58;
               R_3_c59 <= R_3_c58;
               R_4_c59 <= R_4_c58;
               R_5_c59 <= R_5_c58;
               R_6_c59 <= R_6_c58;
               Cin_7_c59 <= Cin_7_c58;
               X_7_c59 <= X_7_c58;
               Y_7_c59 <= Y_7_c58;
               X_8_c59 <= X_8_c58;
               Y_8_c59 <= Y_8_c58;
               X_9_c59 <= X_9_c58;
               Y_9_c59 <= Y_9_c58;
            end if;
            if ce_60 = '1' then
               R_0_c60 <= R_0_c59;
               R_1_c60 <= R_1_c59;
               R_2_c60 <= R_2_c59;
               R_3_c60 <= R_3_c59;
               R_4_c60 <= R_4_c59;
               R_5_c60 <= R_5_c59;
               R_6_c60 <= R_6_c59;
               R_7_c60 <= R_7_c59;
               Cin_8_c60 <= Cin_8_c59;
               X_8_c60 <= X_8_c59;
               Y_8_c60 <= Y_8_c59;
               X_9_c60 <= X_9_c59;
               Y_9_c60 <= Y_9_c59;
            end if;
            if ce_61 = '1' then
               R_0_c61 <= R_0_c60;
               R_1_c61 <= R_1_c60;
               R_2_c61 <= R_2_c60;
               R_3_c61 <= R_3_c60;
               R_4_c61 <= R_4_c60;
               R_5_c61 <= R_5_c60;
               R_6_c61 <= R_6_c60;
               R_7_c61 <= R_7_c60;
               R_8_c61 <= R_8_c60;
               Cin_9_c61 <= Cin_9_c60;
               X_9_c61 <= X_9_c60;
               Y_9_c61 <= Y_9_c60;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c35 <= '0' & X(2 downto 0);
   Y_0_c50 <= '0' & Y(2 downto 0);
   S_0_c51 <= X_0_c51 + Y_0_c51 + Cin_0_c51;
   R_0_c51 <= S_0_c51(2 downto 0);
   Cin_1_c51 <= S_0_c51(3);
   X_1_c35 <= '0' & X(5 downto 3);
   Y_1_c50 <= '0' & Y(5 downto 3);
   S_1_c52 <= X_1_c52 + Y_1_c52 + Cin_1_c52;
   R_1_c52 <= S_1_c52(2 downto 0);
   Cin_2_c52 <= S_1_c52(3);
   X_2_c35 <= '0' & X(8 downto 6);
   Y_2_c50 <= '0' & Y(8 downto 6);
   S_2_c53 <= X_2_c53 + Y_2_c53 + Cin_2_c53;
   R_2_c53 <= S_2_c53(2 downto 0);
   Cin_3_c53 <= S_2_c53(3);
   X_3_c35 <= '0' & X(11 downto 9);
   Y_3_c50 <= '0' & Y(11 downto 9);
   S_3_c55 <= X_3_c55 + Y_3_c55 + Cin_3_c55;
   R_3_c55 <= S_3_c55(2 downto 0);
   Cin_4_c55 <= S_3_c55(3);
   X_4_c35 <= '0' & X(14 downto 12);
   Y_4_c50 <= '0' & Y(14 downto 12);
   S_4_c56 <= X_4_c56 + Y_4_c56 + Cin_4_c56;
   R_4_c56 <= S_4_c56(2 downto 0);
   Cin_5_c56 <= S_4_c56(3);
   X_5_c35 <= '0' & X(17 downto 15);
   Y_5_c50 <= '0' & Y(17 downto 15);
   S_5_c57 <= X_5_c57 + Y_5_c57 + Cin_5_c57;
   R_5_c57 <= S_5_c57(2 downto 0);
   Cin_6_c57 <= S_5_c57(3);
   X_6_c35 <= '0' & X(20 downto 18);
   Y_6_c50 <= '0' & Y(20 downto 18);
   S_6_c58 <= X_6_c58 + Y_6_c58 + Cin_6_c58;
   R_6_c58 <= S_6_c58(2 downto 0);
   Cin_7_c58 <= S_6_c58(3);
   X_7_c35 <= '0' & X(23 downto 21);
   Y_7_c50 <= '0' & Y(23 downto 21);
   S_7_c59 <= X_7_c59 + Y_7_c59 + Cin_7_c59;
   R_7_c59 <= S_7_c59(2 downto 0);
   Cin_8_c59 <= S_7_c59(3);
   X_8_c35 <= '0' & X(26 downto 24);
   Y_8_c50 <= '0' & Y(26 downto 24);
   S_8_c60 <= X_8_c60 + Y_8_c60 + Cin_8_c60;
   R_8_c60 <= S_8_c60(2 downto 0);
   Cin_9_c60 <= S_8_c60(3);
   X_9_c35 <= '0' & X(27 downto 27);
   Y_9_c50 <= '0' & Y(27 downto 27);
   S_9_c61 <= X_9_c61 + Y_9_c61 + Cin_9_c61;
   R_9_c61 <= S_9_c61(0 downto 0);
   R <= R_9_c61 & R_8_c61 & R_7_c61 & R_6_c61 & R_5_c61 & R_4_c61 & R_3_c61 & R_2_c61 & R_1_c61 & R_0_c61 ;
end architecture;

--------------------------------------------------------------------------------
--                           Exp_8_23_Freq800_uid6
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca (2008-2021)
--------------------------------------------------------------------------------
-- Pipeline depth: 61 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: ufixX_i XSign
-- Output signals: expY K

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Exp_8_23_Freq800_uid6 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56, ce_57, ce_58, ce_59, ce_60, ce_61 : in std_logic;
          ufixX_i : in  std_logic_vector(33 downto 0);
          XSign : in  std_logic;
          expY : out  std_logic_vector(27 downto 0);
          K : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of Exp_8_23_Freq800_uid6 is
   component FixRealKCM_Freq800_uid8 is
      port ( clk, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10 : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             R : out  std_logic_vector(7 downto 0)   );
   end component;

   component FixRealKCM_Freq800_uid20 is
      port ( clk, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23 : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             R : out  std_logic_vector(34 downto 0)   );
   end component;

   component IntAdder_27_Freq800_uid33 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32 : in std_logic;
             X : in  std_logic_vector(26 downto 0);
             Y : in  std_logic_vector(26 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(26 downto 0)   );
   end component;

   component FixFunctionByTable_Freq800_uid35 is
      port ( clk, ce_33, ce_34, ce_35 : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(27 downto 0)   );
   end component;

   component FixFunctionByTable_Freq800_uid44 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

   component IntAdder_18_Freq800_uid48 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38 : in std_logic;
             X : in  std_logic_vector(17 downto 0);
             Y : in  std_logic_vector(17 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(17 downto 0)   );
   end component;

   component IntAdder_18_Freq800_uid52 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41 : in std_logic;
             X : in  std_logic_vector(17 downto 0);
             Y : in  std_logic_vector(17 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(17 downto 0)   );
   end component;

   component IntMultiplier_17x18_19_Freq800_uid54 is
      port ( clk, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(17 downto 0);
             R : out  std_logic_vector(18 downto 0)   );
   end component;

   component IntAdder_28_Freq800_uid444 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56, ce_57, ce_58, ce_59, ce_60, ce_61 : in std_logic;
             X : in  std_logic_vector(27 downto 0);
             Y : in  std_logic_vector(27 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(27 downto 0)   );
   end component;

signal ufixX_c4, ufixX_c5 :  unsigned(6+27 downto 0);
signal xMulIn_c4 :  unsigned(6+3 downto 0);
signal absK_c10, absK_c11 :  std_logic_vector(7 downto 0);
signal minusAbsK_c11 :  std_logic_vector(8 downto 0);
signal absKLog2_c23 :  std_logic_vector(34 downto 0);
signal subOp1_c5 :  std_logic_vector(26 downto 0);
signal subOp2_c23 :  std_logic_vector(26 downto 0);
signal Y_c32 :  std_logic_vector(26 downto 0);
signal A_c32 :  std_logic_vector(9 downto 0);
signal Z_c32 :  std_logic_vector(16 downto 0);
signal expA_c35 :  std_logic_vector(27 downto 0);
signal Ztrunc_c32 :  std_logic_vector(6 downto 0);
signal expZmZm1_c32 :  std_logic_vector(5 downto 0);
signal expZmZm1_copy45_c32 :  std_logic_vector(5 downto 0);
signal expZm1adderX_c32 :  std_logic_vector(17 downto 0);
signal expZm1adderY_c32 :  std_logic_vector(17 downto 0);
signal expZm1_c38 :  std_logic_vector(17 downto 0);
signal expA_T_c35 :  std_logic_vector(17 downto 0);
signal expArounded0_c41 :  std_logic_vector(17 downto 0);
signal expArounded_c41 :  std_logic_vector(16 downto 0);
signal lowerProduct_c50 :  std_logic_vector(18 downto 0);
signal extendedLowerProduct_c50 :  std_logic_vector(27 downto 0);
signal XSign_c1, XSign_c2, XSign_c3, XSign_c4, XSign_c5, XSign_c6, XSign_c7, XSign_c8, XSign_c9, XSign_c10, XSign_c11, XSign_c12, XSign_c13, XSign_c14, XSign_c15, XSign_c16, XSign_c17, XSign_c18, XSign_c19, XSign_c20, XSign_c21, XSign_c22, XSign_c23 :  std_logic;
constant g: positive := 4;
constant wE: positive := 8;
constant wF: positive := 23;
constant wFIn: positive := 23;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               XSign_c1 <= XSign;
            end if;
            if ce_2 = '1' then
               XSign_c2 <= XSign_c1;
            end if;
            if ce_3 = '1' then
               XSign_c3 <= XSign_c2;
            end if;
            if ce_4 = '1' then
               XSign_c4 <= XSign_c3;
            end if;
            if ce_5 = '1' then
               ufixX_c5 <= ufixX_c4;
               XSign_c5 <= XSign_c4;
            end if;
            if ce_6 = '1' then
               XSign_c6 <= XSign_c5;
            end if;
            if ce_7 = '1' then
               XSign_c7 <= XSign_c6;
            end if;
            if ce_8 = '1' then
               XSign_c8 <= XSign_c7;
            end if;
            if ce_9 = '1' then
               XSign_c9 <= XSign_c8;
            end if;
            if ce_10 = '1' then
               XSign_c10 <= XSign_c9;
            end if;
            if ce_11 = '1' then
               absK_c11 <= absK_c10;
               XSign_c11 <= XSign_c10;
            end if;
            if ce_12 = '1' then
               XSign_c12 <= XSign_c11;
            end if;
            if ce_13 = '1' then
               XSign_c13 <= XSign_c12;
            end if;
            if ce_14 = '1' then
               XSign_c14 <= XSign_c13;
            end if;
            if ce_15 = '1' then
               XSign_c15 <= XSign_c14;
            end if;
            if ce_16 = '1' then
               XSign_c16 <= XSign_c15;
            end if;
            if ce_17 = '1' then
               XSign_c17 <= XSign_c16;
            end if;
            if ce_18 = '1' then
               XSign_c18 <= XSign_c17;
            end if;
            if ce_19 = '1' then
               XSign_c19 <= XSign_c18;
            end if;
            if ce_20 = '1' then
               XSign_c20 <= XSign_c19;
            end if;
            if ce_21 = '1' then
               XSign_c21 <= XSign_c20;
            end if;
            if ce_22 = '1' then
               XSign_c22 <= XSign_c21;
            end if;
            if ce_23 = '1' then
               XSign_c23 <= XSign_c22;
            end if;
            if ce_24 = '1' then
            end if;
            if ce_25 = '1' then
            end if;
            if ce_26 = '1' then
            end if;
            if ce_27 = '1' then
            end if;
            if ce_28 = '1' then
            end if;
            if ce_29 = '1' then
            end if;
            if ce_30 = '1' then
            end if;
            if ce_31 = '1' then
            end if;
            if ce_32 = '1' then
            end if;
            if ce_33 = '1' then
            end if;
            if ce_34 = '1' then
            end if;
            if ce_35 = '1' then
            end if;
            if ce_36 = '1' then
            end if;
            if ce_37 = '1' then
            end if;
            if ce_38 = '1' then
            end if;
            if ce_39 = '1' then
            end if;
            if ce_40 = '1' then
            end if;
            if ce_41 = '1' then
            end if;
            if ce_42 = '1' then
            end if;
            if ce_43 = '1' then
            end if;
            if ce_44 = '1' then
            end if;
            if ce_45 = '1' then
            end if;
            if ce_46 = '1' then
            end if;
            if ce_47 = '1' then
            end if;
            if ce_48 = '1' then
            end if;
            if ce_49 = '1' then
            end if;
            if ce_50 = '1' then
            end if;
            if ce_51 = '1' then
            end if;
            if ce_52 = '1' then
            end if;
            if ce_53 = '1' then
            end if;
            if ce_54 = '1' then
            end if;
            if ce_55 = '1' then
            end if;
            if ce_56 = '1' then
            end if;
            if ce_57 = '1' then
            end if;
            if ce_58 = '1' then
            end if;
            if ce_59 = '1' then
            end if;
            if ce_60 = '1' then
            end if;
            if ce_61 = '1' then
            end if;
         end if;
      end process;
ufixX_c4 <= unsigned(ufixX_i);
   xMulIn_c4 <= ufixX_c4(33 downto 24); -- fix resize from (6, -27) to (6, -3)
   MulInvLog2: FixRealKCM_Freq800_uid8
      port map ( clk  => clk,
                 ce_5 => ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 X => std_logic_vector(xMulIn_c4),
                 R => absK_c10);
   minusAbsK_c11 <= (8 downto 0 => '0') - ('0' & absK_c11);
   K <= minusAbsK_c11 when  XSign_c11='1'   else ('0' & absK_c11);
   MulLog2: FixRealKCM_Freq800_uid20
      port map ( clk  => clk,
                 ce_11 => ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 X => absK_c10,
                 R => absKLog2_c23);
   subOp1_c5 <= std_logic_vector(ufixX_c5(26 downto 0)) when XSign_c5='0' else not (std_logic_vector(ufixX_c5(26 downto 0)));
   subOp2_c23 <= absKLog2_c23(26 downto 0) when XSign_c23='1' else not (absKLog2_c23(26 downto 0));
   theYAdder: IntAdder_27_Freq800_uid33
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 Cin => '1',
                 X => subOp1_c5,
                 Y => subOp2_c23,
                 R => Y_c32);
   -- Now compute the exp of this fixed-point value
   A_c32 <= Y_c32(26 downto 17);
   Z_c32 <= Y_c32(16 downto 0);
   ExpATable: FixFunctionByTable_Freq800_uid35
      port map ( clk  => clk,
                 ce_33 => ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 X => A_c32,
                 Y => expA_c35);
   Ztrunc_c32 <= Z_c32(16 downto 10);
   ExpZmZm1Table: FixFunctionByTable_Freq800_uid44
      port map ( X => Ztrunc_c32,
                 Y => expZmZm1_copy45_c32);
   expZmZm1_c32 <= expZmZm1_copy45_c32; -- output copy to hold a pipeline register if needed
   -- Computing Z + (exp(Z)-1-Z)
   expZm1adderX_c32 <= '0' & Z_c32;
   expZm1adderY_c32 <= (11 downto 0 => '0') & expZmZm1_c32 ;
   Adder_expZm1: IntAdder_18_Freq800_uid48
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 ce_36=> ce_36,
                 ce_37=> ce_37,
                 ce_38=> ce_38,
                 Cin => '0',
                 X => expZm1adderX_c32,
                 Y => expZm1adderY_c32,
                 R => expZm1_c38);
   -- Rounding expA to the same accuracy as expZm1
   --   (truncation would not be accurate enough and require one more guard bit)
   expA_T_c35 <= expA_c35(27 downto 10);
   Adder_expArounded0: IntAdder_18_Freq800_uid52
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 ce_36=> ce_36,
                 ce_37=> ce_37,
                 ce_38=> ce_38,
                 ce_39=> ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 Cin => '1',
                 X => expA_T_c35,
                 Y => "000000000000000000",
                 R => expArounded0_c41);
   expArounded_c41 <= expArounded0_c41(17 downto 1);
   TheLowerProduct: IntMultiplier_17x18_19_Freq800_uid54
      port map ( clk  => clk,
                 ce_39 => ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 ce_42=> ce_42,
                 ce_43=> ce_43,
                 ce_44=> ce_44,
                 ce_45=> ce_45,
                 ce_46=> ce_46,
                 ce_47=> ce_47,
                 ce_48=> ce_48,
                 ce_49=> ce_49,
                 ce_50=> ce_50,
                 X => expArounded_c41,
                 Y => expZm1_c38,
                 R => lowerProduct_c50);
   extendedLowerProduct_c50 <= ((27 downto 19 => '0') & lowerProduct_c50(18 downto 0));
   -- Final addition -- the product MSB bit weight is -k+2 = -8
   TheFinalAdder: IntAdder_28_Freq800_uid444
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 ce_36=> ce_36,
                 ce_37=> ce_37,
                 ce_38=> ce_38,
                 ce_39=> ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 ce_42=> ce_42,
                 ce_43=> ce_43,
                 ce_44=> ce_44,
                 ce_45=> ce_45,
                 ce_46=> ce_46,
                 ce_47=> ce_47,
                 ce_48=> ce_48,
                 ce_49=> ce_49,
                 ce_50=> ce_50,
                 ce_51=> ce_51,
                 ce_52=> ce_52,
                 ce_53=> ce_53,
                 ce_54=> ce_54,
                 ce_55=> ce_55,
                 ce_56=> ce_56,
                 ce_57=> ce_57,
                 ce_58=> ce_58,
                 ce_59=> ce_59,
                 ce_60=> ce_60,
                 ce_61=> ce_61,
                 Cin => '0',
                 X => expA_c35,
                 Y => extendedLowerProduct_c50,
                 R => expY);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_Freq800_uid447
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 72 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_Freq800_uid447 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56, ce_57, ce_58, ce_59, ce_60, ce_61, ce_62, ce_63, ce_64, ce_65, ce_66, ce_67, ce_68, ce_69, ce_70, ce_71, ce_72 : in std_logic;
          X : in  std_logic_vector(32 downto 0);
          Y : in  std_logic_vector(32 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_Freq800_uid447 is
signal Cin_1_c0, Cin_1_c1, Cin_1_c2, Cin_1_c3, Cin_1_c4, Cin_1_c5, Cin_1_c6, Cin_1_c7, Cin_1_c8, Cin_1_c9, Cin_1_c10, Cin_1_c11, Cin_1_c12, Cin_1_c13, Cin_1_c14, Cin_1_c15, Cin_1_c16, Cin_1_c17, Cin_1_c18, Cin_1_c19, Cin_1_c20, Cin_1_c21, Cin_1_c22, Cin_1_c23, Cin_1_c24, Cin_1_c25, Cin_1_c26, Cin_1_c27, Cin_1_c28, Cin_1_c29, Cin_1_c30, Cin_1_c31, Cin_1_c32, Cin_1_c33, Cin_1_c34, Cin_1_c35, Cin_1_c36, Cin_1_c37, Cin_1_c38, Cin_1_c39, Cin_1_c40, Cin_1_c41, Cin_1_c42, Cin_1_c43, Cin_1_c44, Cin_1_c45, Cin_1_c46, Cin_1_c47, Cin_1_c48, Cin_1_c49, Cin_1_c50, Cin_1_c51, Cin_1_c52, Cin_1_c53, Cin_1_c54, Cin_1_c55, Cin_1_c56, Cin_1_c57, Cin_1_c58, Cin_1_c59, Cin_1_c60, Cin_1_c61, Cin_1_c62 :  std_logic;
signal X_1_c61, X_1_c62 :  std_logic_vector(3 downto 0);
signal Y_1_c61, Y_1_c62 :  std_logic_vector(3 downto 0);
signal S_1_c62 :  std_logic_vector(3 downto 0);
signal R_1_c62, R_1_c63, R_1_c64, R_1_c65, R_1_c66, R_1_c67, R_1_c68, R_1_c69, R_1_c70, R_1_c71, R_1_c72 :  std_logic_vector(2 downto 0);
signal Cin_2_c62, Cin_2_c63 :  std_logic;
signal X_2_c61, X_2_c62, X_2_c63 :  std_logic_vector(3 downto 0);
signal Y_2_c61, Y_2_c62, Y_2_c63 :  std_logic_vector(3 downto 0);
signal S_2_c63 :  std_logic_vector(3 downto 0);
signal R_2_c63, R_2_c64, R_2_c65, R_2_c66, R_2_c67, R_2_c68, R_2_c69, R_2_c70, R_2_c71, R_2_c72 :  std_logic_vector(2 downto 0);
signal Cin_3_c63, Cin_3_c64 :  std_logic;
signal X_3_c61, X_3_c62, X_3_c63, X_3_c64 :  std_logic_vector(3 downto 0);
signal Y_3_c61, Y_3_c62, Y_3_c63, Y_3_c64 :  std_logic_vector(3 downto 0);
signal S_3_c64 :  std_logic_vector(3 downto 0);
signal R_3_c64, R_3_c65, R_3_c66, R_3_c67, R_3_c68, R_3_c69, R_3_c70, R_3_c71, R_3_c72 :  std_logic_vector(2 downto 0);
signal Cin_4_c64, Cin_4_c65 :  std_logic;
signal X_4_c61, X_4_c62, X_4_c63, X_4_c64, X_4_c65 :  std_logic_vector(3 downto 0);
signal Y_4_c61, Y_4_c62, Y_4_c63, Y_4_c64, Y_4_c65 :  std_logic_vector(3 downto 0);
signal S_4_c65 :  std_logic_vector(3 downto 0);
signal R_4_c65, R_4_c66, R_4_c67, R_4_c68, R_4_c69, R_4_c70, R_4_c71, R_4_c72 :  std_logic_vector(2 downto 0);
signal Cin_5_c65, Cin_5_c66 :  std_logic;
signal X_5_c61, X_5_c62, X_5_c63, X_5_c64, X_5_c65, X_5_c66 :  std_logic_vector(3 downto 0);
signal Y_5_c61, Y_5_c62, Y_5_c63, Y_5_c64, Y_5_c65, Y_5_c66 :  std_logic_vector(3 downto 0);
signal S_5_c66 :  std_logic_vector(3 downto 0);
signal R_5_c66, R_5_c67, R_5_c68, R_5_c69, R_5_c70, R_5_c71, R_5_c72 :  std_logic_vector(2 downto 0);
signal Cin_6_c66, Cin_6_c67 :  std_logic;
signal X_6_c61, X_6_c62, X_6_c63, X_6_c64, X_6_c65, X_6_c66, X_6_c67 :  std_logic_vector(3 downto 0);
signal Y_6_c61, Y_6_c62, Y_6_c63, Y_6_c64, Y_6_c65, Y_6_c66, Y_6_c67 :  std_logic_vector(3 downto 0);
signal S_6_c67 :  std_logic_vector(3 downto 0);
signal R_6_c67, R_6_c68, R_6_c69, R_6_c70, R_6_c71, R_6_c72 :  std_logic_vector(2 downto 0);
signal Cin_7_c67, Cin_7_c68 :  std_logic;
signal X_7_c61, X_7_c62, X_7_c63, X_7_c64, X_7_c65, X_7_c66, X_7_c67, X_7_c68 :  std_logic_vector(3 downto 0);
signal Y_7_c61, Y_7_c62, Y_7_c63, Y_7_c64, Y_7_c65, Y_7_c66, Y_7_c67, Y_7_c68 :  std_logic_vector(3 downto 0);
signal S_7_c68 :  std_logic_vector(3 downto 0);
signal R_7_c68, R_7_c69, R_7_c70, R_7_c71, R_7_c72 :  std_logic_vector(2 downto 0);
signal Cin_8_c68, Cin_8_c69 :  std_logic;
signal X_8_c61, X_8_c62, X_8_c63, X_8_c64, X_8_c65, X_8_c66, X_8_c67, X_8_c68, X_8_c69 :  std_logic_vector(3 downto 0);
signal Y_8_c61, Y_8_c62, Y_8_c63, Y_8_c64, Y_8_c65, Y_8_c66, Y_8_c67, Y_8_c68, Y_8_c69 :  std_logic_vector(3 downto 0);
signal S_8_c69 :  std_logic_vector(3 downto 0);
signal R_8_c69, R_8_c70, R_8_c71, R_8_c72 :  std_logic_vector(2 downto 0);
signal Cin_9_c69, Cin_9_c70 :  std_logic;
signal X_9_c61, X_9_c62, X_9_c63, X_9_c64, X_9_c65, X_9_c66, X_9_c67, X_9_c68, X_9_c69, X_9_c70 :  std_logic_vector(3 downto 0);
signal Y_9_c61, Y_9_c62, Y_9_c63, Y_9_c64, Y_9_c65, Y_9_c66, Y_9_c67, Y_9_c68, Y_9_c69, Y_9_c70 :  std_logic_vector(3 downto 0);
signal S_9_c70 :  std_logic_vector(3 downto 0);
signal R_9_c70, R_9_c71, R_9_c72 :  std_logic_vector(2 downto 0);
signal Cin_10_c70, Cin_10_c71 :  std_logic;
signal X_10_c61, X_10_c62, X_10_c63, X_10_c64, X_10_c65, X_10_c66, X_10_c67, X_10_c68, X_10_c69, X_10_c70, X_10_c71 :  std_logic_vector(3 downto 0);
signal Y_10_c61, Y_10_c62, Y_10_c63, Y_10_c64, Y_10_c65, Y_10_c66, Y_10_c67, Y_10_c68, Y_10_c69, Y_10_c70, Y_10_c71 :  std_logic_vector(3 downto 0);
signal S_10_c71 :  std_logic_vector(3 downto 0);
signal R_10_c71, R_10_c72 :  std_logic_vector(2 downto 0);
signal Cin_11_c71, Cin_11_c72 :  std_logic;
signal X_11_c61, X_11_c62, X_11_c63, X_11_c64, X_11_c65, X_11_c66, X_11_c67, X_11_c68, X_11_c69, X_11_c70, X_11_c71, X_11_c72 :  std_logic_vector(3 downto 0);
signal Y_11_c61, Y_11_c62, Y_11_c63, Y_11_c64, Y_11_c65, Y_11_c66, Y_11_c67, Y_11_c68, Y_11_c69, Y_11_c70, Y_11_c71, Y_11_c72 :  std_logic_vector(3 downto 0);
signal S_11_c72 :  std_logic_vector(3 downto 0);
signal R_11_c72 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_1_c1 <= Cin_1_c0;
            end if;
            if ce_2 = '1' then
               Cin_1_c2 <= Cin_1_c1;
            end if;
            if ce_3 = '1' then
               Cin_1_c3 <= Cin_1_c2;
            end if;
            if ce_4 = '1' then
               Cin_1_c4 <= Cin_1_c3;
            end if;
            if ce_5 = '1' then
               Cin_1_c5 <= Cin_1_c4;
            end if;
            if ce_6 = '1' then
               Cin_1_c6 <= Cin_1_c5;
            end if;
            if ce_7 = '1' then
               Cin_1_c7 <= Cin_1_c6;
            end if;
            if ce_8 = '1' then
               Cin_1_c8 <= Cin_1_c7;
            end if;
            if ce_9 = '1' then
               Cin_1_c9 <= Cin_1_c8;
            end if;
            if ce_10 = '1' then
               Cin_1_c10 <= Cin_1_c9;
            end if;
            if ce_11 = '1' then
               Cin_1_c11 <= Cin_1_c10;
            end if;
            if ce_12 = '1' then
               Cin_1_c12 <= Cin_1_c11;
            end if;
            if ce_13 = '1' then
               Cin_1_c13 <= Cin_1_c12;
            end if;
            if ce_14 = '1' then
               Cin_1_c14 <= Cin_1_c13;
            end if;
            if ce_15 = '1' then
               Cin_1_c15 <= Cin_1_c14;
            end if;
            if ce_16 = '1' then
               Cin_1_c16 <= Cin_1_c15;
            end if;
            if ce_17 = '1' then
               Cin_1_c17 <= Cin_1_c16;
            end if;
            if ce_18 = '1' then
               Cin_1_c18 <= Cin_1_c17;
            end if;
            if ce_19 = '1' then
               Cin_1_c19 <= Cin_1_c18;
            end if;
            if ce_20 = '1' then
               Cin_1_c20 <= Cin_1_c19;
            end if;
            if ce_21 = '1' then
               Cin_1_c21 <= Cin_1_c20;
            end if;
            if ce_22 = '1' then
               Cin_1_c22 <= Cin_1_c21;
            end if;
            if ce_23 = '1' then
               Cin_1_c23 <= Cin_1_c22;
            end if;
            if ce_24 = '1' then
               Cin_1_c24 <= Cin_1_c23;
            end if;
            if ce_25 = '1' then
               Cin_1_c25 <= Cin_1_c24;
            end if;
            if ce_26 = '1' then
               Cin_1_c26 <= Cin_1_c25;
            end if;
            if ce_27 = '1' then
               Cin_1_c27 <= Cin_1_c26;
            end if;
            if ce_28 = '1' then
               Cin_1_c28 <= Cin_1_c27;
            end if;
            if ce_29 = '1' then
               Cin_1_c29 <= Cin_1_c28;
            end if;
            if ce_30 = '1' then
               Cin_1_c30 <= Cin_1_c29;
            end if;
            if ce_31 = '1' then
               Cin_1_c31 <= Cin_1_c30;
            end if;
            if ce_32 = '1' then
               Cin_1_c32 <= Cin_1_c31;
            end if;
            if ce_33 = '1' then
               Cin_1_c33 <= Cin_1_c32;
            end if;
            if ce_34 = '1' then
               Cin_1_c34 <= Cin_1_c33;
            end if;
            if ce_35 = '1' then
               Cin_1_c35 <= Cin_1_c34;
            end if;
            if ce_36 = '1' then
               Cin_1_c36 <= Cin_1_c35;
            end if;
            if ce_37 = '1' then
               Cin_1_c37 <= Cin_1_c36;
            end if;
            if ce_38 = '1' then
               Cin_1_c38 <= Cin_1_c37;
            end if;
            if ce_39 = '1' then
               Cin_1_c39 <= Cin_1_c38;
            end if;
            if ce_40 = '1' then
               Cin_1_c40 <= Cin_1_c39;
            end if;
            if ce_41 = '1' then
               Cin_1_c41 <= Cin_1_c40;
            end if;
            if ce_42 = '1' then
               Cin_1_c42 <= Cin_1_c41;
            end if;
            if ce_43 = '1' then
               Cin_1_c43 <= Cin_1_c42;
            end if;
            if ce_44 = '1' then
               Cin_1_c44 <= Cin_1_c43;
            end if;
            if ce_45 = '1' then
               Cin_1_c45 <= Cin_1_c44;
            end if;
            if ce_46 = '1' then
               Cin_1_c46 <= Cin_1_c45;
            end if;
            if ce_47 = '1' then
               Cin_1_c47 <= Cin_1_c46;
            end if;
            if ce_48 = '1' then
               Cin_1_c48 <= Cin_1_c47;
            end if;
            if ce_49 = '1' then
               Cin_1_c49 <= Cin_1_c48;
            end if;
            if ce_50 = '1' then
               Cin_1_c50 <= Cin_1_c49;
            end if;
            if ce_51 = '1' then
               Cin_1_c51 <= Cin_1_c50;
            end if;
            if ce_52 = '1' then
               Cin_1_c52 <= Cin_1_c51;
            end if;
            if ce_53 = '1' then
               Cin_1_c53 <= Cin_1_c52;
            end if;
            if ce_54 = '1' then
               Cin_1_c54 <= Cin_1_c53;
            end if;
            if ce_55 = '1' then
               Cin_1_c55 <= Cin_1_c54;
            end if;
            if ce_56 = '1' then
               Cin_1_c56 <= Cin_1_c55;
            end if;
            if ce_57 = '1' then
               Cin_1_c57 <= Cin_1_c56;
            end if;
            if ce_58 = '1' then
               Cin_1_c58 <= Cin_1_c57;
            end if;
            if ce_59 = '1' then
               Cin_1_c59 <= Cin_1_c58;
            end if;
            if ce_60 = '1' then
               Cin_1_c60 <= Cin_1_c59;
            end if;
            if ce_61 = '1' then
               Cin_1_c61 <= Cin_1_c60;
            end if;
            if ce_62 = '1' then
               Cin_1_c62 <= Cin_1_c61;
               X_1_c62 <= X_1_c61;
               Y_1_c62 <= Y_1_c61;
               X_2_c62 <= X_2_c61;
               Y_2_c62 <= Y_2_c61;
               X_3_c62 <= X_3_c61;
               Y_3_c62 <= Y_3_c61;
               X_4_c62 <= X_4_c61;
               Y_4_c62 <= Y_4_c61;
               X_5_c62 <= X_5_c61;
               Y_5_c62 <= Y_5_c61;
               X_6_c62 <= X_6_c61;
               Y_6_c62 <= Y_6_c61;
               X_7_c62 <= X_7_c61;
               Y_7_c62 <= Y_7_c61;
               X_8_c62 <= X_8_c61;
               Y_8_c62 <= Y_8_c61;
               X_9_c62 <= X_9_c61;
               Y_9_c62 <= Y_9_c61;
               X_10_c62 <= X_10_c61;
               Y_10_c62 <= Y_10_c61;
               X_11_c62 <= X_11_c61;
               Y_11_c62 <= Y_11_c61;
            end if;
            if ce_63 = '1' then
               R_1_c63 <= R_1_c62;
               Cin_2_c63 <= Cin_2_c62;
               X_2_c63 <= X_2_c62;
               Y_2_c63 <= Y_2_c62;
               X_3_c63 <= X_3_c62;
               Y_3_c63 <= Y_3_c62;
               X_4_c63 <= X_4_c62;
               Y_4_c63 <= Y_4_c62;
               X_5_c63 <= X_5_c62;
               Y_5_c63 <= Y_5_c62;
               X_6_c63 <= X_6_c62;
               Y_6_c63 <= Y_6_c62;
               X_7_c63 <= X_7_c62;
               Y_7_c63 <= Y_7_c62;
               X_8_c63 <= X_8_c62;
               Y_8_c63 <= Y_8_c62;
               X_9_c63 <= X_9_c62;
               Y_9_c63 <= Y_9_c62;
               X_10_c63 <= X_10_c62;
               Y_10_c63 <= Y_10_c62;
               X_11_c63 <= X_11_c62;
               Y_11_c63 <= Y_11_c62;
            end if;
            if ce_64 = '1' then
               R_1_c64 <= R_1_c63;
               R_2_c64 <= R_2_c63;
               Cin_3_c64 <= Cin_3_c63;
               X_3_c64 <= X_3_c63;
               Y_3_c64 <= Y_3_c63;
               X_4_c64 <= X_4_c63;
               Y_4_c64 <= Y_4_c63;
               X_5_c64 <= X_5_c63;
               Y_5_c64 <= Y_5_c63;
               X_6_c64 <= X_6_c63;
               Y_6_c64 <= Y_6_c63;
               X_7_c64 <= X_7_c63;
               Y_7_c64 <= Y_7_c63;
               X_8_c64 <= X_8_c63;
               Y_8_c64 <= Y_8_c63;
               X_9_c64 <= X_9_c63;
               Y_9_c64 <= Y_9_c63;
               X_10_c64 <= X_10_c63;
               Y_10_c64 <= Y_10_c63;
               X_11_c64 <= X_11_c63;
               Y_11_c64 <= Y_11_c63;
            end if;
            if ce_65 = '1' then
               R_1_c65 <= R_1_c64;
               R_2_c65 <= R_2_c64;
               R_3_c65 <= R_3_c64;
               Cin_4_c65 <= Cin_4_c64;
               X_4_c65 <= X_4_c64;
               Y_4_c65 <= Y_4_c64;
               X_5_c65 <= X_5_c64;
               Y_5_c65 <= Y_5_c64;
               X_6_c65 <= X_6_c64;
               Y_6_c65 <= Y_6_c64;
               X_7_c65 <= X_7_c64;
               Y_7_c65 <= Y_7_c64;
               X_8_c65 <= X_8_c64;
               Y_8_c65 <= Y_8_c64;
               X_9_c65 <= X_9_c64;
               Y_9_c65 <= Y_9_c64;
               X_10_c65 <= X_10_c64;
               Y_10_c65 <= Y_10_c64;
               X_11_c65 <= X_11_c64;
               Y_11_c65 <= Y_11_c64;
            end if;
            if ce_66 = '1' then
               R_1_c66 <= R_1_c65;
               R_2_c66 <= R_2_c65;
               R_3_c66 <= R_3_c65;
               R_4_c66 <= R_4_c65;
               Cin_5_c66 <= Cin_5_c65;
               X_5_c66 <= X_5_c65;
               Y_5_c66 <= Y_5_c65;
               X_6_c66 <= X_6_c65;
               Y_6_c66 <= Y_6_c65;
               X_7_c66 <= X_7_c65;
               Y_7_c66 <= Y_7_c65;
               X_8_c66 <= X_8_c65;
               Y_8_c66 <= Y_8_c65;
               X_9_c66 <= X_9_c65;
               Y_9_c66 <= Y_9_c65;
               X_10_c66 <= X_10_c65;
               Y_10_c66 <= Y_10_c65;
               X_11_c66 <= X_11_c65;
               Y_11_c66 <= Y_11_c65;
            end if;
            if ce_67 = '1' then
               R_1_c67 <= R_1_c66;
               R_2_c67 <= R_2_c66;
               R_3_c67 <= R_3_c66;
               R_4_c67 <= R_4_c66;
               R_5_c67 <= R_5_c66;
               Cin_6_c67 <= Cin_6_c66;
               X_6_c67 <= X_6_c66;
               Y_6_c67 <= Y_6_c66;
               X_7_c67 <= X_7_c66;
               Y_7_c67 <= Y_7_c66;
               X_8_c67 <= X_8_c66;
               Y_8_c67 <= Y_8_c66;
               X_9_c67 <= X_9_c66;
               Y_9_c67 <= Y_9_c66;
               X_10_c67 <= X_10_c66;
               Y_10_c67 <= Y_10_c66;
               X_11_c67 <= X_11_c66;
               Y_11_c67 <= Y_11_c66;
            end if;
            if ce_68 = '1' then
               R_1_c68 <= R_1_c67;
               R_2_c68 <= R_2_c67;
               R_3_c68 <= R_3_c67;
               R_4_c68 <= R_4_c67;
               R_5_c68 <= R_5_c67;
               R_6_c68 <= R_6_c67;
               Cin_7_c68 <= Cin_7_c67;
               X_7_c68 <= X_7_c67;
               Y_7_c68 <= Y_7_c67;
               X_8_c68 <= X_8_c67;
               Y_8_c68 <= Y_8_c67;
               X_9_c68 <= X_9_c67;
               Y_9_c68 <= Y_9_c67;
               X_10_c68 <= X_10_c67;
               Y_10_c68 <= Y_10_c67;
               X_11_c68 <= X_11_c67;
               Y_11_c68 <= Y_11_c67;
            end if;
            if ce_69 = '1' then
               R_1_c69 <= R_1_c68;
               R_2_c69 <= R_2_c68;
               R_3_c69 <= R_3_c68;
               R_4_c69 <= R_4_c68;
               R_5_c69 <= R_5_c68;
               R_6_c69 <= R_6_c68;
               R_7_c69 <= R_7_c68;
               Cin_8_c69 <= Cin_8_c68;
               X_8_c69 <= X_8_c68;
               Y_8_c69 <= Y_8_c68;
               X_9_c69 <= X_9_c68;
               Y_9_c69 <= Y_9_c68;
               X_10_c69 <= X_10_c68;
               Y_10_c69 <= Y_10_c68;
               X_11_c69 <= X_11_c68;
               Y_11_c69 <= Y_11_c68;
            end if;
            if ce_70 = '1' then
               R_1_c70 <= R_1_c69;
               R_2_c70 <= R_2_c69;
               R_3_c70 <= R_3_c69;
               R_4_c70 <= R_4_c69;
               R_5_c70 <= R_5_c69;
               R_6_c70 <= R_6_c69;
               R_7_c70 <= R_7_c69;
               R_8_c70 <= R_8_c69;
               Cin_9_c70 <= Cin_9_c69;
               X_9_c70 <= X_9_c69;
               Y_9_c70 <= Y_9_c69;
               X_10_c70 <= X_10_c69;
               Y_10_c70 <= Y_10_c69;
               X_11_c70 <= X_11_c69;
               Y_11_c70 <= Y_11_c69;
            end if;
            if ce_71 = '1' then
               R_1_c71 <= R_1_c70;
               R_2_c71 <= R_2_c70;
               R_3_c71 <= R_3_c70;
               R_4_c71 <= R_4_c70;
               R_5_c71 <= R_5_c70;
               R_6_c71 <= R_6_c70;
               R_7_c71 <= R_7_c70;
               R_8_c71 <= R_8_c70;
               R_9_c71 <= R_9_c70;
               Cin_10_c71 <= Cin_10_c70;
               X_10_c71 <= X_10_c70;
               Y_10_c71 <= Y_10_c70;
               X_11_c71 <= X_11_c70;
               Y_11_c71 <= Y_11_c70;
            end if;
            if ce_72 = '1' then
               R_1_c72 <= R_1_c71;
               R_2_c72 <= R_2_c71;
               R_3_c72 <= R_3_c71;
               R_4_c72 <= R_4_c71;
               R_5_c72 <= R_5_c71;
               R_6_c72 <= R_6_c71;
               R_7_c72 <= R_7_c71;
               R_8_c72 <= R_8_c71;
               R_9_c72 <= R_9_c71;
               R_10_c72 <= R_10_c71;
               Cin_11_c72 <= Cin_11_c71;
               X_11_c72 <= X_11_c71;
               Y_11_c72 <= Y_11_c71;
            end if;
         end if;
      end process;
   Cin_1_c0 <= Cin;
   X_1_c61 <= '0' & X(2 downto 0);
   Y_1_c61 <= '0' & Y(2 downto 0);
   S_1_c62 <= X_1_c62 + Y_1_c62 + Cin_1_c62;
   R_1_c62 <= S_1_c62(2 downto 0);
   Cin_2_c62 <= S_1_c62(3);
   X_2_c61 <= '0' & X(5 downto 3);
   Y_2_c61 <= '0' & Y(5 downto 3);
   S_2_c63 <= X_2_c63 + Y_2_c63 + Cin_2_c63;
   R_2_c63 <= S_2_c63(2 downto 0);
   Cin_3_c63 <= S_2_c63(3);
   X_3_c61 <= '0' & X(8 downto 6);
   Y_3_c61 <= '0' & Y(8 downto 6);
   S_3_c64 <= X_3_c64 + Y_3_c64 + Cin_3_c64;
   R_3_c64 <= S_3_c64(2 downto 0);
   Cin_4_c64 <= S_3_c64(3);
   X_4_c61 <= '0' & X(11 downto 9);
   Y_4_c61 <= '0' & Y(11 downto 9);
   S_4_c65 <= X_4_c65 + Y_4_c65 + Cin_4_c65;
   R_4_c65 <= S_4_c65(2 downto 0);
   Cin_5_c65 <= S_4_c65(3);
   X_5_c61 <= '0' & X(14 downto 12);
   Y_5_c61 <= '0' & Y(14 downto 12);
   S_5_c66 <= X_5_c66 + Y_5_c66 + Cin_5_c66;
   R_5_c66 <= S_5_c66(2 downto 0);
   Cin_6_c66 <= S_5_c66(3);
   X_6_c61 <= '0' & X(17 downto 15);
   Y_6_c61 <= '0' & Y(17 downto 15);
   S_6_c67 <= X_6_c67 + Y_6_c67 + Cin_6_c67;
   R_6_c67 <= S_6_c67(2 downto 0);
   Cin_7_c67 <= S_6_c67(3);
   X_7_c61 <= '0' & X(20 downto 18);
   Y_7_c61 <= '0' & Y(20 downto 18);
   S_7_c68 <= X_7_c68 + Y_7_c68 + Cin_7_c68;
   R_7_c68 <= S_7_c68(2 downto 0);
   Cin_8_c68 <= S_7_c68(3);
   X_8_c61 <= '0' & X(23 downto 21);
   Y_8_c61 <= '0' & Y(23 downto 21);
   S_8_c69 <= X_8_c69 + Y_8_c69 + Cin_8_c69;
   R_8_c69 <= S_8_c69(2 downto 0);
   Cin_9_c69 <= S_8_c69(3);
   X_9_c61 <= '0' & X(26 downto 24);
   Y_9_c61 <= '0' & Y(26 downto 24);
   S_9_c70 <= X_9_c70 + Y_9_c70 + Cin_9_c70;
   R_9_c70 <= S_9_c70(2 downto 0);
   Cin_10_c70 <= S_9_c70(3);
   X_10_c61 <= '0' & X(29 downto 27);
   Y_10_c61 <= '0' & Y(29 downto 27);
   S_10_c71 <= X_10_c71 + Y_10_c71 + Cin_10_c71;
   R_10_c71 <= S_10_c71(2 downto 0);
   Cin_11_c71 <= S_10_c71(3);
   X_11_c61 <= '0' & X(32 downto 30);
   Y_11_c61 <= '0' & Y(32 downto 30);
   S_11_c72 <= X_11_c72 + Y_11_c72 + Cin_11_c72;
   R_11_c72 <= S_11_c72(2 downto 0);
   R <= R_11_c72 & R_10_c72 & R_9_c72 & R_8_c72 & R_7_c72 & R_6_c72 & R_5_c72 & R_4_c72 & R_3_c72 & R_2_c72 & R_1_c72 ;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointExponential
--                         (FPExp_8_23_Freq800_uid2)
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, Bogdan Pasca (2008-2021)
--------------------------------------------------------------------------------
-- Pipeline depth: 73 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointExponential is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56, ce_57, ce_58, ce_59, ce_60, ce_61, ce_62, ce_63, ce_64, ce_65, ce_66, ce_67, ce_68, ce_69, ce_70, ce_71, ce_72, ce_73 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointExponential is
   component LeftShifter24_by_max_33_Freq800_uid4 is
      port ( clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             S : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(56 downto 0)   );
   end component;

   component Exp_8_23_Freq800_uid6 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56, ce_57, ce_58, ce_59, ce_60, ce_61 : in std_logic;
             ufixX_i : in  std_logic_vector(33 downto 0);
             XSign : in  std_logic;
             expY : out  std_logic_vector(27 downto 0);
             K : out  std_logic_vector(8 downto 0)   );
   end component;

   component IntAdder_33_Freq800_uid447 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56, ce_57, ce_58, ce_59, ce_60, ce_61, ce_62, ce_63, ce_64, ce_65, ce_66, ce_67, ce_68, ce_69, ce_70, ce_71, ce_72 : in std_logic;
             X : in  std_logic_vector(32 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(32 downto 0)   );
   end component;

signal Xexn_c0, Xexn_c1, Xexn_c2, Xexn_c3, Xexn_c4, Xexn_c5, Xexn_c6, Xexn_c7, Xexn_c8, Xexn_c9, Xexn_c10, Xexn_c11, Xexn_c12, Xexn_c13, Xexn_c14, Xexn_c15, Xexn_c16, Xexn_c17, Xexn_c18, Xexn_c19, Xexn_c20, Xexn_c21, Xexn_c22, Xexn_c23, Xexn_c24, Xexn_c25, Xexn_c26, Xexn_c27, Xexn_c28, Xexn_c29, Xexn_c30, Xexn_c31, Xexn_c32, Xexn_c33, Xexn_c34, Xexn_c35, Xexn_c36, Xexn_c37, Xexn_c38, Xexn_c39, Xexn_c40, Xexn_c41, Xexn_c42, Xexn_c43, Xexn_c44, Xexn_c45, Xexn_c46, Xexn_c47, Xexn_c48, Xexn_c49, Xexn_c50, Xexn_c51, Xexn_c52, Xexn_c53, Xexn_c54, Xexn_c55, Xexn_c56, Xexn_c57, Xexn_c58, Xexn_c59, Xexn_c60, Xexn_c61, Xexn_c62, Xexn_c63, Xexn_c64, Xexn_c65, Xexn_c66, Xexn_c67, Xexn_c68, Xexn_c69, Xexn_c70, Xexn_c71, Xexn_c72, Xexn_c73 :  std_logic_vector(1 downto 0);
signal XSign_c0, XSign_c1, XSign_c2, XSign_c3, XSign_c4, XSign_c5, XSign_c6, XSign_c7, XSign_c8, XSign_c9, XSign_c10, XSign_c11, XSign_c12, XSign_c13, XSign_c14, XSign_c15, XSign_c16, XSign_c17, XSign_c18, XSign_c19, XSign_c20, XSign_c21, XSign_c22, XSign_c23, XSign_c24, XSign_c25, XSign_c26, XSign_c27, XSign_c28, XSign_c29, XSign_c30, XSign_c31, XSign_c32, XSign_c33, XSign_c34, XSign_c35, XSign_c36, XSign_c37, XSign_c38, XSign_c39, XSign_c40, XSign_c41, XSign_c42, XSign_c43, XSign_c44, XSign_c45, XSign_c46, XSign_c47, XSign_c48, XSign_c49, XSign_c50, XSign_c51, XSign_c52, XSign_c53, XSign_c54, XSign_c55, XSign_c56, XSign_c57, XSign_c58, XSign_c59, XSign_c60, XSign_c61, XSign_c62, XSign_c63, XSign_c64, XSign_c65, XSign_c66, XSign_c67, XSign_c68, XSign_c69, XSign_c70, XSign_c71, XSign_c72, XSign_c73 :  std_logic;
signal XexpField_c0, XexpField_c1 :  std_logic_vector(7 downto 0);
signal Xfrac_c0 :  unsigned(-1+23 downto 0);
signal e0_c0, e0_c1 :  std_logic_vector(9 downto 0);
signal shiftVal_c1, shiftVal_c2 :  std_logic_vector(9 downto 0);
signal resultWillBeOne_c1, resultWillBeOne_c2, resultWillBeOne_c3, resultWillBeOne_c4 :  std_logic;
signal mXu_c0 :  unsigned(0+23 downto 0);
signal maxShift_c0, maxShift_c1, maxShift_c2 :  std_logic_vector(8 downto 0);
signal overflow0_c2 :  std_logic;
signal shiftValIn_c1 :  std_logic_vector(5 downto 0);
signal fixX0_c4 :  std_logic_vector(56 downto 0);
signal ufixX_c4 :  unsigned(6+27 downto 0);
signal expY_c61 :  std_logic_vector(27 downto 0);
signal K_c11, K_c12, K_c13, K_c14, K_c15, K_c16, K_c17, K_c18, K_c19, K_c20, K_c21, K_c22, K_c23, K_c24, K_c25, K_c26, K_c27, K_c28, K_c29, K_c30, K_c31, K_c32, K_c33, K_c34, K_c35, K_c36, K_c37, K_c38, K_c39, K_c40, K_c41, K_c42, K_c43, K_c44, K_c45, K_c46, K_c47, K_c48, K_c49, K_c50, K_c51, K_c52, K_c53, K_c54, K_c55, K_c56, K_c57, K_c58, K_c59, K_c60, K_c61 :  std_logic_vector(8 downto 0);
signal needNoNorm_c61 :  std_logic;
signal preRoundBiasSig_c61 :  std_logic_vector(32 downto 0);
signal roundBit_c61 :  std_logic;
signal roundNormAddend_c61 :  std_logic_vector(32 downto 0);
signal roundedExpSigRes_c72, roundedExpSigRes_c73 :  std_logic_vector(32 downto 0);
signal roundedExpSig_c73 :  std_logic_vector(32 downto 0);
signal ofl1_c2, ofl1_c3, ofl1_c4, ofl1_c5, ofl1_c6, ofl1_c7, ofl1_c8, ofl1_c9, ofl1_c10, ofl1_c11, ofl1_c12, ofl1_c13, ofl1_c14, ofl1_c15, ofl1_c16, ofl1_c17, ofl1_c18, ofl1_c19, ofl1_c20, ofl1_c21, ofl1_c22, ofl1_c23, ofl1_c24, ofl1_c25, ofl1_c26, ofl1_c27, ofl1_c28, ofl1_c29, ofl1_c30, ofl1_c31, ofl1_c32, ofl1_c33, ofl1_c34, ofl1_c35, ofl1_c36, ofl1_c37, ofl1_c38, ofl1_c39, ofl1_c40, ofl1_c41, ofl1_c42, ofl1_c43, ofl1_c44, ofl1_c45, ofl1_c46, ofl1_c47, ofl1_c48, ofl1_c49, ofl1_c50, ofl1_c51, ofl1_c52, ofl1_c53, ofl1_c54, ofl1_c55, ofl1_c56, ofl1_c57, ofl1_c58, ofl1_c59, ofl1_c60, ofl1_c61, ofl1_c62, ofl1_c63, ofl1_c64, ofl1_c65, ofl1_c66, ofl1_c67, ofl1_c68, ofl1_c69, ofl1_c70, ofl1_c71, ofl1_c72, ofl1_c73 :  std_logic;
signal ofl2_c73 :  std_logic;
signal ofl3_c0, ofl3_c1, ofl3_c2, ofl3_c3, ofl3_c4, ofl3_c5, ofl3_c6, ofl3_c7, ofl3_c8, ofl3_c9, ofl3_c10, ofl3_c11, ofl3_c12, ofl3_c13, ofl3_c14, ofl3_c15, ofl3_c16, ofl3_c17, ofl3_c18, ofl3_c19, ofl3_c20, ofl3_c21, ofl3_c22, ofl3_c23, ofl3_c24, ofl3_c25, ofl3_c26, ofl3_c27, ofl3_c28, ofl3_c29, ofl3_c30, ofl3_c31, ofl3_c32, ofl3_c33, ofl3_c34, ofl3_c35, ofl3_c36, ofl3_c37, ofl3_c38, ofl3_c39, ofl3_c40, ofl3_c41, ofl3_c42, ofl3_c43, ofl3_c44, ofl3_c45, ofl3_c46, ofl3_c47, ofl3_c48, ofl3_c49, ofl3_c50, ofl3_c51, ofl3_c52, ofl3_c53, ofl3_c54, ofl3_c55, ofl3_c56, ofl3_c57, ofl3_c58, ofl3_c59, ofl3_c60, ofl3_c61, ofl3_c62, ofl3_c63, ofl3_c64, ofl3_c65, ofl3_c66, ofl3_c67, ofl3_c68, ofl3_c69, ofl3_c70, ofl3_c71, ofl3_c72, ofl3_c73 :  std_logic;
signal ofl_c73 :  std_logic;
signal ufl1_c73 :  std_logic;
signal ufl2_c0, ufl2_c1, ufl2_c2, ufl2_c3, ufl2_c4, ufl2_c5, ufl2_c6, ufl2_c7, ufl2_c8, ufl2_c9, ufl2_c10, ufl2_c11, ufl2_c12, ufl2_c13, ufl2_c14, ufl2_c15, ufl2_c16, ufl2_c17, ufl2_c18, ufl2_c19, ufl2_c20, ufl2_c21, ufl2_c22, ufl2_c23, ufl2_c24, ufl2_c25, ufl2_c26, ufl2_c27, ufl2_c28, ufl2_c29, ufl2_c30, ufl2_c31, ufl2_c32, ufl2_c33, ufl2_c34, ufl2_c35, ufl2_c36, ufl2_c37, ufl2_c38, ufl2_c39, ufl2_c40, ufl2_c41, ufl2_c42, ufl2_c43, ufl2_c44, ufl2_c45, ufl2_c46, ufl2_c47, ufl2_c48, ufl2_c49, ufl2_c50, ufl2_c51, ufl2_c52, ufl2_c53, ufl2_c54, ufl2_c55, ufl2_c56, ufl2_c57, ufl2_c58, ufl2_c59, ufl2_c60, ufl2_c61, ufl2_c62, ufl2_c63, ufl2_c64, ufl2_c65, ufl2_c66, ufl2_c67, ufl2_c68, ufl2_c69, ufl2_c70, ufl2_c71, ufl2_c72, ufl2_c73 :  std_logic;
signal ufl3_c2, ufl3_c3, ufl3_c4, ufl3_c5, ufl3_c6, ufl3_c7, ufl3_c8, ufl3_c9, ufl3_c10, ufl3_c11, ufl3_c12, ufl3_c13, ufl3_c14, ufl3_c15, ufl3_c16, ufl3_c17, ufl3_c18, ufl3_c19, ufl3_c20, ufl3_c21, ufl3_c22, ufl3_c23, ufl3_c24, ufl3_c25, ufl3_c26, ufl3_c27, ufl3_c28, ufl3_c29, ufl3_c30, ufl3_c31, ufl3_c32, ufl3_c33, ufl3_c34, ufl3_c35, ufl3_c36, ufl3_c37, ufl3_c38, ufl3_c39, ufl3_c40, ufl3_c41, ufl3_c42, ufl3_c43, ufl3_c44, ufl3_c45, ufl3_c46, ufl3_c47, ufl3_c48, ufl3_c49, ufl3_c50, ufl3_c51, ufl3_c52, ufl3_c53, ufl3_c54, ufl3_c55, ufl3_c56, ufl3_c57, ufl3_c58, ufl3_c59, ufl3_c60, ufl3_c61, ufl3_c62, ufl3_c63, ufl3_c64, ufl3_c65, ufl3_c66, ufl3_c67, ufl3_c68, ufl3_c69, ufl3_c70, ufl3_c71, ufl3_c72, ufl3_c73 :  std_logic;
signal ufl_c73 :  std_logic;
signal Rexn_c73 :  std_logic_vector(1 downto 0);
constant g: positive := 4;
constant wE: positive := 8;
constant wF: positive := 23;
constant wFIn: positive := 23;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Xexn_c1 <= Xexn_c0;
               XSign_c1 <= XSign_c0;
               XexpField_c1 <= XexpField_c0;
               e0_c1 <= e0_c0;
               maxShift_c1 <= maxShift_c0;
               ofl3_c1 <= ofl3_c0;
               ufl2_c1 <= ufl2_c0;
            end if;
            if ce_2 = '1' then
               Xexn_c2 <= Xexn_c1;
               XSign_c2 <= XSign_c1;
               shiftVal_c2 <= shiftVal_c1;
               resultWillBeOne_c2 <= resultWillBeOne_c1;
               maxShift_c2 <= maxShift_c1;
               ofl3_c2 <= ofl3_c1;
               ufl2_c2 <= ufl2_c1;
            end if;
            if ce_3 = '1' then
               Xexn_c3 <= Xexn_c2;
               XSign_c3 <= XSign_c2;
               resultWillBeOne_c3 <= resultWillBeOne_c2;
               ofl1_c3 <= ofl1_c2;
               ofl3_c3 <= ofl3_c2;
               ufl2_c3 <= ufl2_c2;
               ufl3_c3 <= ufl3_c2;
            end if;
            if ce_4 = '1' then
               Xexn_c4 <= Xexn_c3;
               XSign_c4 <= XSign_c3;
               resultWillBeOne_c4 <= resultWillBeOne_c3;
               ofl1_c4 <= ofl1_c3;
               ofl3_c4 <= ofl3_c3;
               ufl2_c4 <= ufl2_c3;
               ufl3_c4 <= ufl3_c3;
            end if;
            if ce_5 = '1' then
               Xexn_c5 <= Xexn_c4;
               XSign_c5 <= XSign_c4;
               ofl1_c5 <= ofl1_c4;
               ofl3_c5 <= ofl3_c4;
               ufl2_c5 <= ufl2_c4;
               ufl3_c5 <= ufl3_c4;
            end if;
            if ce_6 = '1' then
               Xexn_c6 <= Xexn_c5;
               XSign_c6 <= XSign_c5;
               ofl1_c6 <= ofl1_c5;
               ofl3_c6 <= ofl3_c5;
               ufl2_c6 <= ufl2_c5;
               ufl3_c6 <= ufl3_c5;
            end if;
            if ce_7 = '1' then
               Xexn_c7 <= Xexn_c6;
               XSign_c7 <= XSign_c6;
               ofl1_c7 <= ofl1_c6;
               ofl3_c7 <= ofl3_c6;
               ufl2_c7 <= ufl2_c6;
               ufl3_c7 <= ufl3_c6;
            end if;
            if ce_8 = '1' then
               Xexn_c8 <= Xexn_c7;
               XSign_c8 <= XSign_c7;
               ofl1_c8 <= ofl1_c7;
               ofl3_c8 <= ofl3_c7;
               ufl2_c8 <= ufl2_c7;
               ufl3_c8 <= ufl3_c7;
            end if;
            if ce_9 = '1' then
               Xexn_c9 <= Xexn_c8;
               XSign_c9 <= XSign_c8;
               ofl1_c9 <= ofl1_c8;
               ofl3_c9 <= ofl3_c8;
               ufl2_c9 <= ufl2_c8;
               ufl3_c9 <= ufl3_c8;
            end if;
            if ce_10 = '1' then
               Xexn_c10 <= Xexn_c9;
               XSign_c10 <= XSign_c9;
               ofl1_c10 <= ofl1_c9;
               ofl3_c10 <= ofl3_c9;
               ufl2_c10 <= ufl2_c9;
               ufl3_c10 <= ufl3_c9;
            end if;
            if ce_11 = '1' then
               Xexn_c11 <= Xexn_c10;
               XSign_c11 <= XSign_c10;
               ofl1_c11 <= ofl1_c10;
               ofl3_c11 <= ofl3_c10;
               ufl2_c11 <= ufl2_c10;
               ufl3_c11 <= ufl3_c10;
            end if;
            if ce_12 = '1' then
               Xexn_c12 <= Xexn_c11;
               XSign_c12 <= XSign_c11;
               K_c12 <= K_c11;
               ofl1_c12 <= ofl1_c11;
               ofl3_c12 <= ofl3_c11;
               ufl2_c12 <= ufl2_c11;
               ufl3_c12 <= ufl3_c11;
            end if;
            if ce_13 = '1' then
               Xexn_c13 <= Xexn_c12;
               XSign_c13 <= XSign_c12;
               K_c13 <= K_c12;
               ofl1_c13 <= ofl1_c12;
               ofl3_c13 <= ofl3_c12;
               ufl2_c13 <= ufl2_c12;
               ufl3_c13 <= ufl3_c12;
            end if;
            if ce_14 = '1' then
               Xexn_c14 <= Xexn_c13;
               XSign_c14 <= XSign_c13;
               K_c14 <= K_c13;
               ofl1_c14 <= ofl1_c13;
               ofl3_c14 <= ofl3_c13;
               ufl2_c14 <= ufl2_c13;
               ufl3_c14 <= ufl3_c13;
            end if;
            if ce_15 = '1' then
               Xexn_c15 <= Xexn_c14;
               XSign_c15 <= XSign_c14;
               K_c15 <= K_c14;
               ofl1_c15 <= ofl1_c14;
               ofl3_c15 <= ofl3_c14;
               ufl2_c15 <= ufl2_c14;
               ufl3_c15 <= ufl3_c14;
            end if;
            if ce_16 = '1' then
               Xexn_c16 <= Xexn_c15;
               XSign_c16 <= XSign_c15;
               K_c16 <= K_c15;
               ofl1_c16 <= ofl1_c15;
               ofl3_c16 <= ofl3_c15;
               ufl2_c16 <= ufl2_c15;
               ufl3_c16 <= ufl3_c15;
            end if;
            if ce_17 = '1' then
               Xexn_c17 <= Xexn_c16;
               XSign_c17 <= XSign_c16;
               K_c17 <= K_c16;
               ofl1_c17 <= ofl1_c16;
               ofl3_c17 <= ofl3_c16;
               ufl2_c17 <= ufl2_c16;
               ufl3_c17 <= ufl3_c16;
            end if;
            if ce_18 = '1' then
               Xexn_c18 <= Xexn_c17;
               XSign_c18 <= XSign_c17;
               K_c18 <= K_c17;
               ofl1_c18 <= ofl1_c17;
               ofl3_c18 <= ofl3_c17;
               ufl2_c18 <= ufl2_c17;
               ufl3_c18 <= ufl3_c17;
            end if;
            if ce_19 = '1' then
               Xexn_c19 <= Xexn_c18;
               XSign_c19 <= XSign_c18;
               K_c19 <= K_c18;
               ofl1_c19 <= ofl1_c18;
               ofl3_c19 <= ofl3_c18;
               ufl2_c19 <= ufl2_c18;
               ufl3_c19 <= ufl3_c18;
            end if;
            if ce_20 = '1' then
               Xexn_c20 <= Xexn_c19;
               XSign_c20 <= XSign_c19;
               K_c20 <= K_c19;
               ofl1_c20 <= ofl1_c19;
               ofl3_c20 <= ofl3_c19;
               ufl2_c20 <= ufl2_c19;
               ufl3_c20 <= ufl3_c19;
            end if;
            if ce_21 = '1' then
               Xexn_c21 <= Xexn_c20;
               XSign_c21 <= XSign_c20;
               K_c21 <= K_c20;
               ofl1_c21 <= ofl1_c20;
               ofl3_c21 <= ofl3_c20;
               ufl2_c21 <= ufl2_c20;
               ufl3_c21 <= ufl3_c20;
            end if;
            if ce_22 = '1' then
               Xexn_c22 <= Xexn_c21;
               XSign_c22 <= XSign_c21;
               K_c22 <= K_c21;
               ofl1_c22 <= ofl1_c21;
               ofl3_c22 <= ofl3_c21;
               ufl2_c22 <= ufl2_c21;
               ufl3_c22 <= ufl3_c21;
            end if;
            if ce_23 = '1' then
               Xexn_c23 <= Xexn_c22;
               XSign_c23 <= XSign_c22;
               K_c23 <= K_c22;
               ofl1_c23 <= ofl1_c22;
               ofl3_c23 <= ofl3_c22;
               ufl2_c23 <= ufl2_c22;
               ufl3_c23 <= ufl3_c22;
            end if;
            if ce_24 = '1' then
               Xexn_c24 <= Xexn_c23;
               XSign_c24 <= XSign_c23;
               K_c24 <= K_c23;
               ofl1_c24 <= ofl1_c23;
               ofl3_c24 <= ofl3_c23;
               ufl2_c24 <= ufl2_c23;
               ufl3_c24 <= ufl3_c23;
            end if;
            if ce_25 = '1' then
               Xexn_c25 <= Xexn_c24;
               XSign_c25 <= XSign_c24;
               K_c25 <= K_c24;
               ofl1_c25 <= ofl1_c24;
               ofl3_c25 <= ofl3_c24;
               ufl2_c25 <= ufl2_c24;
               ufl3_c25 <= ufl3_c24;
            end if;
            if ce_26 = '1' then
               Xexn_c26 <= Xexn_c25;
               XSign_c26 <= XSign_c25;
               K_c26 <= K_c25;
               ofl1_c26 <= ofl1_c25;
               ofl3_c26 <= ofl3_c25;
               ufl2_c26 <= ufl2_c25;
               ufl3_c26 <= ufl3_c25;
            end if;
            if ce_27 = '1' then
               Xexn_c27 <= Xexn_c26;
               XSign_c27 <= XSign_c26;
               K_c27 <= K_c26;
               ofl1_c27 <= ofl1_c26;
               ofl3_c27 <= ofl3_c26;
               ufl2_c27 <= ufl2_c26;
               ufl3_c27 <= ufl3_c26;
            end if;
            if ce_28 = '1' then
               Xexn_c28 <= Xexn_c27;
               XSign_c28 <= XSign_c27;
               K_c28 <= K_c27;
               ofl1_c28 <= ofl1_c27;
               ofl3_c28 <= ofl3_c27;
               ufl2_c28 <= ufl2_c27;
               ufl3_c28 <= ufl3_c27;
            end if;
            if ce_29 = '1' then
               Xexn_c29 <= Xexn_c28;
               XSign_c29 <= XSign_c28;
               K_c29 <= K_c28;
               ofl1_c29 <= ofl1_c28;
               ofl3_c29 <= ofl3_c28;
               ufl2_c29 <= ufl2_c28;
               ufl3_c29 <= ufl3_c28;
            end if;
            if ce_30 = '1' then
               Xexn_c30 <= Xexn_c29;
               XSign_c30 <= XSign_c29;
               K_c30 <= K_c29;
               ofl1_c30 <= ofl1_c29;
               ofl3_c30 <= ofl3_c29;
               ufl2_c30 <= ufl2_c29;
               ufl3_c30 <= ufl3_c29;
            end if;
            if ce_31 = '1' then
               Xexn_c31 <= Xexn_c30;
               XSign_c31 <= XSign_c30;
               K_c31 <= K_c30;
               ofl1_c31 <= ofl1_c30;
               ofl3_c31 <= ofl3_c30;
               ufl2_c31 <= ufl2_c30;
               ufl3_c31 <= ufl3_c30;
            end if;
            if ce_32 = '1' then
               Xexn_c32 <= Xexn_c31;
               XSign_c32 <= XSign_c31;
               K_c32 <= K_c31;
               ofl1_c32 <= ofl1_c31;
               ofl3_c32 <= ofl3_c31;
               ufl2_c32 <= ufl2_c31;
               ufl3_c32 <= ufl3_c31;
            end if;
            if ce_33 = '1' then
               Xexn_c33 <= Xexn_c32;
               XSign_c33 <= XSign_c32;
               K_c33 <= K_c32;
               ofl1_c33 <= ofl1_c32;
               ofl3_c33 <= ofl3_c32;
               ufl2_c33 <= ufl2_c32;
               ufl3_c33 <= ufl3_c32;
            end if;
            if ce_34 = '1' then
               Xexn_c34 <= Xexn_c33;
               XSign_c34 <= XSign_c33;
               K_c34 <= K_c33;
               ofl1_c34 <= ofl1_c33;
               ofl3_c34 <= ofl3_c33;
               ufl2_c34 <= ufl2_c33;
               ufl3_c34 <= ufl3_c33;
            end if;
            if ce_35 = '1' then
               Xexn_c35 <= Xexn_c34;
               XSign_c35 <= XSign_c34;
               K_c35 <= K_c34;
               ofl1_c35 <= ofl1_c34;
               ofl3_c35 <= ofl3_c34;
               ufl2_c35 <= ufl2_c34;
               ufl3_c35 <= ufl3_c34;
            end if;
            if ce_36 = '1' then
               Xexn_c36 <= Xexn_c35;
               XSign_c36 <= XSign_c35;
               K_c36 <= K_c35;
               ofl1_c36 <= ofl1_c35;
               ofl3_c36 <= ofl3_c35;
               ufl2_c36 <= ufl2_c35;
               ufl3_c36 <= ufl3_c35;
            end if;
            if ce_37 = '1' then
               Xexn_c37 <= Xexn_c36;
               XSign_c37 <= XSign_c36;
               K_c37 <= K_c36;
               ofl1_c37 <= ofl1_c36;
               ofl3_c37 <= ofl3_c36;
               ufl2_c37 <= ufl2_c36;
               ufl3_c37 <= ufl3_c36;
            end if;
            if ce_38 = '1' then
               Xexn_c38 <= Xexn_c37;
               XSign_c38 <= XSign_c37;
               K_c38 <= K_c37;
               ofl1_c38 <= ofl1_c37;
               ofl3_c38 <= ofl3_c37;
               ufl2_c38 <= ufl2_c37;
               ufl3_c38 <= ufl3_c37;
            end if;
            if ce_39 = '1' then
               Xexn_c39 <= Xexn_c38;
               XSign_c39 <= XSign_c38;
               K_c39 <= K_c38;
               ofl1_c39 <= ofl1_c38;
               ofl3_c39 <= ofl3_c38;
               ufl2_c39 <= ufl2_c38;
               ufl3_c39 <= ufl3_c38;
            end if;
            if ce_40 = '1' then
               Xexn_c40 <= Xexn_c39;
               XSign_c40 <= XSign_c39;
               K_c40 <= K_c39;
               ofl1_c40 <= ofl1_c39;
               ofl3_c40 <= ofl3_c39;
               ufl2_c40 <= ufl2_c39;
               ufl3_c40 <= ufl3_c39;
            end if;
            if ce_41 = '1' then
               Xexn_c41 <= Xexn_c40;
               XSign_c41 <= XSign_c40;
               K_c41 <= K_c40;
               ofl1_c41 <= ofl1_c40;
               ofl3_c41 <= ofl3_c40;
               ufl2_c41 <= ufl2_c40;
               ufl3_c41 <= ufl3_c40;
            end if;
            if ce_42 = '1' then
               Xexn_c42 <= Xexn_c41;
               XSign_c42 <= XSign_c41;
               K_c42 <= K_c41;
               ofl1_c42 <= ofl1_c41;
               ofl3_c42 <= ofl3_c41;
               ufl2_c42 <= ufl2_c41;
               ufl3_c42 <= ufl3_c41;
            end if;
            if ce_43 = '1' then
               Xexn_c43 <= Xexn_c42;
               XSign_c43 <= XSign_c42;
               K_c43 <= K_c42;
               ofl1_c43 <= ofl1_c42;
               ofl3_c43 <= ofl3_c42;
               ufl2_c43 <= ufl2_c42;
               ufl3_c43 <= ufl3_c42;
            end if;
            if ce_44 = '1' then
               Xexn_c44 <= Xexn_c43;
               XSign_c44 <= XSign_c43;
               K_c44 <= K_c43;
               ofl1_c44 <= ofl1_c43;
               ofl3_c44 <= ofl3_c43;
               ufl2_c44 <= ufl2_c43;
               ufl3_c44 <= ufl3_c43;
            end if;
            if ce_45 = '1' then
               Xexn_c45 <= Xexn_c44;
               XSign_c45 <= XSign_c44;
               K_c45 <= K_c44;
               ofl1_c45 <= ofl1_c44;
               ofl3_c45 <= ofl3_c44;
               ufl2_c45 <= ufl2_c44;
               ufl3_c45 <= ufl3_c44;
            end if;
            if ce_46 = '1' then
               Xexn_c46 <= Xexn_c45;
               XSign_c46 <= XSign_c45;
               K_c46 <= K_c45;
               ofl1_c46 <= ofl1_c45;
               ofl3_c46 <= ofl3_c45;
               ufl2_c46 <= ufl2_c45;
               ufl3_c46 <= ufl3_c45;
            end if;
            if ce_47 = '1' then
               Xexn_c47 <= Xexn_c46;
               XSign_c47 <= XSign_c46;
               K_c47 <= K_c46;
               ofl1_c47 <= ofl1_c46;
               ofl3_c47 <= ofl3_c46;
               ufl2_c47 <= ufl2_c46;
               ufl3_c47 <= ufl3_c46;
            end if;
            if ce_48 = '1' then
               Xexn_c48 <= Xexn_c47;
               XSign_c48 <= XSign_c47;
               K_c48 <= K_c47;
               ofl1_c48 <= ofl1_c47;
               ofl3_c48 <= ofl3_c47;
               ufl2_c48 <= ufl2_c47;
               ufl3_c48 <= ufl3_c47;
            end if;
            if ce_49 = '1' then
               Xexn_c49 <= Xexn_c48;
               XSign_c49 <= XSign_c48;
               K_c49 <= K_c48;
               ofl1_c49 <= ofl1_c48;
               ofl3_c49 <= ofl3_c48;
               ufl2_c49 <= ufl2_c48;
               ufl3_c49 <= ufl3_c48;
            end if;
            if ce_50 = '1' then
               Xexn_c50 <= Xexn_c49;
               XSign_c50 <= XSign_c49;
               K_c50 <= K_c49;
               ofl1_c50 <= ofl1_c49;
               ofl3_c50 <= ofl3_c49;
               ufl2_c50 <= ufl2_c49;
               ufl3_c50 <= ufl3_c49;
            end if;
            if ce_51 = '1' then
               Xexn_c51 <= Xexn_c50;
               XSign_c51 <= XSign_c50;
               K_c51 <= K_c50;
               ofl1_c51 <= ofl1_c50;
               ofl3_c51 <= ofl3_c50;
               ufl2_c51 <= ufl2_c50;
               ufl3_c51 <= ufl3_c50;
            end if;
            if ce_52 = '1' then
               Xexn_c52 <= Xexn_c51;
               XSign_c52 <= XSign_c51;
               K_c52 <= K_c51;
               ofl1_c52 <= ofl1_c51;
               ofl3_c52 <= ofl3_c51;
               ufl2_c52 <= ufl2_c51;
               ufl3_c52 <= ufl3_c51;
            end if;
            if ce_53 = '1' then
               Xexn_c53 <= Xexn_c52;
               XSign_c53 <= XSign_c52;
               K_c53 <= K_c52;
               ofl1_c53 <= ofl1_c52;
               ofl3_c53 <= ofl3_c52;
               ufl2_c53 <= ufl2_c52;
               ufl3_c53 <= ufl3_c52;
            end if;
            if ce_54 = '1' then
               Xexn_c54 <= Xexn_c53;
               XSign_c54 <= XSign_c53;
               K_c54 <= K_c53;
               ofl1_c54 <= ofl1_c53;
               ofl3_c54 <= ofl3_c53;
               ufl2_c54 <= ufl2_c53;
               ufl3_c54 <= ufl3_c53;
            end if;
            if ce_55 = '1' then
               Xexn_c55 <= Xexn_c54;
               XSign_c55 <= XSign_c54;
               K_c55 <= K_c54;
               ofl1_c55 <= ofl1_c54;
               ofl3_c55 <= ofl3_c54;
               ufl2_c55 <= ufl2_c54;
               ufl3_c55 <= ufl3_c54;
            end if;
            if ce_56 = '1' then
               Xexn_c56 <= Xexn_c55;
               XSign_c56 <= XSign_c55;
               K_c56 <= K_c55;
               ofl1_c56 <= ofl1_c55;
               ofl3_c56 <= ofl3_c55;
               ufl2_c56 <= ufl2_c55;
               ufl3_c56 <= ufl3_c55;
            end if;
            if ce_57 = '1' then
               Xexn_c57 <= Xexn_c56;
               XSign_c57 <= XSign_c56;
               K_c57 <= K_c56;
               ofl1_c57 <= ofl1_c56;
               ofl3_c57 <= ofl3_c56;
               ufl2_c57 <= ufl2_c56;
               ufl3_c57 <= ufl3_c56;
            end if;
            if ce_58 = '1' then
               Xexn_c58 <= Xexn_c57;
               XSign_c58 <= XSign_c57;
               K_c58 <= K_c57;
               ofl1_c58 <= ofl1_c57;
               ofl3_c58 <= ofl3_c57;
               ufl2_c58 <= ufl2_c57;
               ufl3_c58 <= ufl3_c57;
            end if;
            if ce_59 = '1' then
               Xexn_c59 <= Xexn_c58;
               XSign_c59 <= XSign_c58;
               K_c59 <= K_c58;
               ofl1_c59 <= ofl1_c58;
               ofl3_c59 <= ofl3_c58;
               ufl2_c59 <= ufl2_c58;
               ufl3_c59 <= ufl3_c58;
            end if;
            if ce_60 = '1' then
               Xexn_c60 <= Xexn_c59;
               XSign_c60 <= XSign_c59;
               K_c60 <= K_c59;
               ofl1_c60 <= ofl1_c59;
               ofl3_c60 <= ofl3_c59;
               ufl2_c60 <= ufl2_c59;
               ufl3_c60 <= ufl3_c59;
            end if;
            if ce_61 = '1' then
               Xexn_c61 <= Xexn_c60;
               XSign_c61 <= XSign_c60;
               K_c61 <= K_c60;
               ofl1_c61 <= ofl1_c60;
               ofl3_c61 <= ofl3_c60;
               ufl2_c61 <= ufl2_c60;
               ufl3_c61 <= ufl3_c60;
            end if;
            if ce_62 = '1' then
               Xexn_c62 <= Xexn_c61;
               XSign_c62 <= XSign_c61;
               ofl1_c62 <= ofl1_c61;
               ofl3_c62 <= ofl3_c61;
               ufl2_c62 <= ufl2_c61;
               ufl3_c62 <= ufl3_c61;
            end if;
            if ce_63 = '1' then
               Xexn_c63 <= Xexn_c62;
               XSign_c63 <= XSign_c62;
               ofl1_c63 <= ofl1_c62;
               ofl3_c63 <= ofl3_c62;
               ufl2_c63 <= ufl2_c62;
               ufl3_c63 <= ufl3_c62;
            end if;
            if ce_64 = '1' then
               Xexn_c64 <= Xexn_c63;
               XSign_c64 <= XSign_c63;
               ofl1_c64 <= ofl1_c63;
               ofl3_c64 <= ofl3_c63;
               ufl2_c64 <= ufl2_c63;
               ufl3_c64 <= ufl3_c63;
            end if;
            if ce_65 = '1' then
               Xexn_c65 <= Xexn_c64;
               XSign_c65 <= XSign_c64;
               ofl1_c65 <= ofl1_c64;
               ofl3_c65 <= ofl3_c64;
               ufl2_c65 <= ufl2_c64;
               ufl3_c65 <= ufl3_c64;
            end if;
            if ce_66 = '1' then
               Xexn_c66 <= Xexn_c65;
               XSign_c66 <= XSign_c65;
               ofl1_c66 <= ofl1_c65;
               ofl3_c66 <= ofl3_c65;
               ufl2_c66 <= ufl2_c65;
               ufl3_c66 <= ufl3_c65;
            end if;
            if ce_67 = '1' then
               Xexn_c67 <= Xexn_c66;
               XSign_c67 <= XSign_c66;
               ofl1_c67 <= ofl1_c66;
               ofl3_c67 <= ofl3_c66;
               ufl2_c67 <= ufl2_c66;
               ufl3_c67 <= ufl3_c66;
            end if;
            if ce_68 = '1' then
               Xexn_c68 <= Xexn_c67;
               XSign_c68 <= XSign_c67;
               ofl1_c68 <= ofl1_c67;
               ofl3_c68 <= ofl3_c67;
               ufl2_c68 <= ufl2_c67;
               ufl3_c68 <= ufl3_c67;
            end if;
            if ce_69 = '1' then
               Xexn_c69 <= Xexn_c68;
               XSign_c69 <= XSign_c68;
               ofl1_c69 <= ofl1_c68;
               ofl3_c69 <= ofl3_c68;
               ufl2_c69 <= ufl2_c68;
               ufl3_c69 <= ufl3_c68;
            end if;
            if ce_70 = '1' then
               Xexn_c70 <= Xexn_c69;
               XSign_c70 <= XSign_c69;
               ofl1_c70 <= ofl1_c69;
               ofl3_c70 <= ofl3_c69;
               ufl2_c70 <= ufl2_c69;
               ufl3_c70 <= ufl3_c69;
            end if;
            if ce_71 = '1' then
               Xexn_c71 <= Xexn_c70;
               XSign_c71 <= XSign_c70;
               ofl1_c71 <= ofl1_c70;
               ofl3_c71 <= ofl3_c70;
               ufl2_c71 <= ufl2_c70;
               ufl3_c71 <= ufl3_c70;
            end if;
            if ce_72 = '1' then
               Xexn_c72 <= Xexn_c71;
               XSign_c72 <= XSign_c71;
               ofl1_c72 <= ofl1_c71;
               ofl3_c72 <= ofl3_c71;
               ufl2_c72 <= ufl2_c71;
               ufl3_c72 <= ufl3_c71;
            end if;
            if ce_73 = '1' then
               Xexn_c73 <= Xexn_c72;
               XSign_c73 <= XSign_c72;
               roundedExpSigRes_c73 <= roundedExpSigRes_c72;
               ofl1_c73 <= ofl1_c72;
               ofl3_c73 <= ofl3_c72;
               ufl2_c73 <= ufl2_c72;
               ufl3_c73 <= ufl3_c72;
            end if;
         end if;
      end process;
   Xexn_c0 <= X(wE+wFIn+2 downto wE+wFIn+1);
   XSign_c0 <= X(wE+wFIn);
   XexpField_c0 <= X(wE+wFIn-1 downto wFIn);
   Xfrac_c0 <= unsigned(X(wFIn-1 downto 0));
   e0_c0 <= conv_std_logic_vector(100, wE+2);  -- bias - (wF+g)
   shiftVal_c1 <= ("00" & XexpField_c1) - e0_c1; -- for a left shift
   -- underflow when input is shifted to zero (shiftval<0), in which case exp = 1
   resultWillBeOne_c1 <= shiftVal_c1(wE+1);
   --  mantissa with implicit bit
   mXu_c0 <= "1" & Xfrac_c0;
   -- Partial overflow detection
   maxShift_c0 <= conv_std_logic_vector(33, wE+1);  -- wE-2 + wF+g
   overflow0_c2 <= not shiftVal_c2(wE+1) when shiftVal_c2(wE downto 0) > maxShift_c2 else '0';
   shiftValIn_c1 <= shiftVal_c1(5 downto 0);
   mantissa_shift: LeftShifter24_by_max_33_Freq800_uid4
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 S => shiftValIn_c1,
                 X => std_logic_vector(mXu_c0),
                 R => fixX0_c4);
   ufixX_c4 <=  unsigned(fixX0_c4(56 downto 23)) when resultWillBeOne_c4='0' else "0000000000000000000000000000000000";
   exp_helper: Exp_8_23_Freq800_uid6
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 ce_36=> ce_36,
                 ce_37=> ce_37,
                 ce_38=> ce_38,
                 ce_39=> ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 ce_42=> ce_42,
                 ce_43=> ce_43,
                 ce_44=> ce_44,
                 ce_45=> ce_45,
                 ce_46=> ce_46,
                 ce_47=> ce_47,
                 ce_48=> ce_48,
                 ce_49=> ce_49,
                 ce_50=> ce_50,
                 ce_51=> ce_51,
                 ce_52=> ce_52,
                 ce_53=> ce_53,
                 ce_54=> ce_54,
                 ce_55=> ce_55,
                 ce_56=> ce_56,
                 ce_57=> ce_57,
                 ce_58=> ce_58,
                 ce_59=> ce_59,
                 ce_60=> ce_60,
                 ce_61=> ce_61,
                 XSign => XSign_c0,
                 ufixX_i => std_logic_vector(ufixX_c4),
                 K => K_c11,
                 expY => expY_c61);
   needNoNorm_c61 <= expY_c61(27);
   -- Rounding: all this should consume one row of LUTs
   preRoundBiasSig_c61 <= conv_std_logic_vector(127, wE+2)  & expY_c61(26 downto 4) when needNoNorm_c61 = '1'
      else conv_std_logic_vector(126, wE+2)  & expY_c61(25 downto 3) ;
   roundBit_c61 <= expY_c61(3)  when needNoNorm_c61 = '1'    else expY_c61(2) ;
   roundNormAddend_c61 <= K_c61(8) & K_c61 & (22 downto 1 => '0') & roundBit_c61;
   roundedExpSigOperandAdder: IntAdder_33_Freq800_uid447
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 ce_36=> ce_36,
                 ce_37=> ce_37,
                 ce_38=> ce_38,
                 ce_39=> ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 ce_42=> ce_42,
                 ce_43=> ce_43,
                 ce_44=> ce_44,
                 ce_45=> ce_45,
                 ce_46=> ce_46,
                 ce_47=> ce_47,
                 ce_48=> ce_48,
                 ce_49=> ce_49,
                 ce_50=> ce_50,
                 ce_51=> ce_51,
                 ce_52=> ce_52,
                 ce_53=> ce_53,
                 ce_54=> ce_54,
                 ce_55=> ce_55,
                 ce_56=> ce_56,
                 ce_57=> ce_57,
                 ce_58=> ce_58,
                 ce_59=> ce_59,
                 ce_60=> ce_60,
                 ce_61=> ce_61,
                 ce_62=> ce_62,
                 ce_63=> ce_63,
                 ce_64=> ce_64,
                 ce_65=> ce_65,
                 ce_66=> ce_66,
                 ce_67=> ce_67,
                 ce_68=> ce_68,
                 ce_69=> ce_69,
                 ce_70=> ce_70,
                 ce_71=> ce_71,
                 ce_72=> ce_72,
                 Cin => '0',
                 X => preRoundBiasSig_c61,
                 Y => roundNormAddend_c61,
                 R => roundedExpSigRes_c72);
   roundedExpSig_c73 <= roundedExpSigRes_c73 when Xexn_c73="01" else  "000" & (wE-2 downto 0 => '1') & (wF-1 downto 0 => '0');
   ofl1_c2 <= not XSign_c2 and overflow0_c2 and (not Xexn_c2(1) and Xexn_c2(0)); -- input positive, normal,  very large
   ofl2_c73 <= not XSign_c73 and (roundedExpSig_c73(wE+wF) and not roundedExpSig_c73(wE+wF+1)) and (not Xexn_c73(1) and Xexn_c73(0)); -- input positive, normal, overflowed
   ofl3_c0 <= not XSign_c0 and Xexn_c0(1) and not Xexn_c0(0);  -- input was -infty
   ofl_c73 <= ofl1_c73 or ofl2_c73 or ofl3_c73;
   ufl1_c73 <= (roundedExpSig_c73(wE+wF) and roundedExpSig_c73(wE+wF+1))  and (not Xexn_c73(1) and Xexn_c73(0)); -- input normal
   ufl2_c0 <= XSign_c0 and Xexn_c0(1) and not Xexn_c0(0);  -- input was -infty
   ufl3_c2 <= XSign_c2 and overflow0_c2  and (not Xexn_c2(1) and Xexn_c2(0)); -- input negative, normal,  very large
   ufl_c73 <= ufl1_c73 or ufl2_c73 or ufl3_c73;
   Rexn_c73 <= "11" when Xexn_c73 = "11"
      else "10" when ofl_c73='1'
      else "00" when ufl_c73='1'
      else "01";
   R <= Rexn_c73 & '0' & roundedExpSig_c73(30 downto 0);
end architecture;



