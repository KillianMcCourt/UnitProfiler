--------------------------------------------------------------------------------
--                RightShifterSticky53_by_max_55_Freq500_uid4
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifterSticky53_by_max_55_Freq500_uid4 is
    port (clk, ce_2, ce_3, ce_4, ce_5 : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          S : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(54 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of RightShifterSticky53_by_max_55_Freq500_uid4 is
signal ps_c1, ps_c2, ps_c3, ps_c4, ps_c5 :  std_logic_vector(5 downto 0);
signal Xpadded_c1 :  std_logic_vector(54 downto 0);
signal level6_c1, level6_c2 :  std_logic_vector(54 downto 0);
signal stk5_c2, stk5_c3 :  std_logic;
signal level5_c1, level5_c2, level5_c3 :  std_logic_vector(54 downto 0);
signal stk4_c3 :  std_logic;
signal level4_c2, level4_c3 :  std_logic_vector(54 downto 0);
signal stk3_c3, stk3_c4 :  std_logic;
signal level3_c2, level3_c3, level3_c4 :  std_logic_vector(54 downto 0);
signal stk2_c4 :  std_logic;
signal level2_c2, level2_c3, level2_c4 :  std_logic_vector(54 downto 0);
signal stk1_c4, stk1_c5 :  std_logic;
signal level1_c2, level1_c3, level1_c4, level1_c5 :  std_logic_vector(54 downto 0);
signal stk0_c5 :  std_logic;
signal level0_c2 :  std_logic_vector(54 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_2 = '1' then
               ps_c2 <= ps_c1;
               level6_c2 <= level6_c1;
               level5_c2 <= level5_c1;
            end if;
            if ce_3 = '1' then
               ps_c3 <= ps_c2;
               stk5_c3 <= stk5_c2;
               level5_c3 <= level5_c2;
               level4_c3 <= level4_c2;
               level3_c3 <= level3_c2;
               level2_c3 <= level2_c2;
               level1_c3 <= level1_c2;
            end if;
            if ce_4 = '1' then
               ps_c4 <= ps_c3;
               stk3_c4 <= stk3_c3;
               level3_c4 <= level3_c3;
               level2_c4 <= level2_c3;
               level1_c4 <= level1_c3;
            end if;
            if ce_5 = '1' then
               ps_c5 <= ps_c4;
               stk1_c5 <= stk1_c4;
               level1_c5 <= level1_c4;
            end if;
         end if;
      end process;
   ps_c1<= S;
   Xpadded_c1 <= X&(1 downto 0 => '0');
   level6_c1<= Xpadded_c1;
   stk5_c2 <= '1' when (level6_c2(31 downto 0)/="00000000000000000000000000000000" and ps_c2(5)='1')   else '0';
   level5_c1 <=  level6_c1 when  ps_c1(5)='0'    else (31 downto 0 => '0') & level6_c1(54 downto 32);
   stk4_c3 <= '1' when (level5_c3(15 downto 0)/="0000000000000000" and ps_c3(4)='1') or stk5_c3 ='1'   else '0';
   level4_c2 <=  level5_c2 when  ps_c2(4)='0'    else (15 downto 0 => '0') & level5_c2(54 downto 16);
   stk3_c3 <= '1' when (level4_c3(7 downto 0)/="00000000" and ps_c3(3)='1') or stk4_c3 ='1'   else '0';
   level3_c2 <=  level4_c2 when  ps_c2(3)='0'    else (7 downto 0 => '0') & level4_c2(54 downto 8);
   stk2_c4 <= '1' when (level3_c4(3 downto 0)/="0000" and ps_c4(2)='1') or stk3_c4 ='1'   else '0';
   level2_c2 <=  level3_c2 when  ps_c2(2)='0'    else (3 downto 0 => '0') & level3_c2(54 downto 4);
   stk1_c4 <= '1' when (level2_c4(1 downto 0)/="00" and ps_c4(1)='1') or stk2_c4 ='1'   else '0';
   level1_c2 <=  level2_c2 when  ps_c2(1)='0'    else (1 downto 0 => '0') & level2_c2(54 downto 2);
   stk0_c5 <= '1' when (level1_c5(0 downto 0)/="0" and ps_c5(0)='1') or stk1_c5 ='1'   else '0';
   level0_c2 <=  level1_c2 when  ps_c2(0)='0'    else (0 downto 0 => '0') & level1_c2(54 downto 1);
   R <= level0_c2;
   Sticky <= stk0_c5;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_56_Freq500_uid6
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_56_Freq500_uid6 is
    port (clk, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntAdder_56_Freq500_uid6 is
signal Cin_1_c5, Cin_1_c6 :  std_logic;
signal X_1_c1, X_1_c2, X_1_c3, X_1_c4, X_1_c5, X_1_c6 :  std_logic_vector(56 downto 0);
signal Y_1_c2, Y_1_c3, Y_1_c4, Y_1_c5, Y_1_c6 :  std_logic_vector(56 downto 0);
signal S_1_c6 :  std_logic_vector(56 downto 0);
signal R_1_c6 :  std_logic_vector(55 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_2 = '1' then
               X_1_c2 <= X_1_c1;
            end if;
            if ce_3 = '1' then
               X_1_c3 <= X_1_c2;
               Y_1_c3 <= Y_1_c2;
            end if;
            if ce_4 = '1' then
               X_1_c4 <= X_1_c3;
               Y_1_c4 <= Y_1_c3;
            end if;
            if ce_5 = '1' then
               X_1_c5 <= X_1_c4;
               Y_1_c5 <= Y_1_c4;
            end if;
            if ce_6 = '1' then
               Cin_1_c6 <= Cin_1_c5;
               X_1_c6 <= X_1_c5;
               Y_1_c6 <= Y_1_c5;
            end if;
         end if;
      end process;
   Cin_1_c5 <= Cin;
   X_1_c1 <= '0' & X(55 downto 0);
   Y_1_c2 <= '0' & Y(55 downto 0);
   S_1_c6 <= X_1_c6 + Y_1_c6 + Cin_1_c6;
   R_1_c6 <= S_1_c6(55 downto 0);
   R <= R_1_c6 ;
end architecture;

--------------------------------------------------------------------------------
--                     Normalizer_Z_57_57_57_Freq500_uid8
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_57_57_57_Freq500_uid8 is
    port (clk, ce_7, ce_8, ce_9, ce_10 : in std_logic;
          X : in  std_logic_vector(56 downto 0);
          Count : out  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of Normalizer_Z_57_57_57_Freq500_uid8 is
signal level6_c6, level6_c7 :  std_logic_vector(56 downto 0);
signal count5_c7, count5_c8, count5_c9, count5_c10 :  std_logic;
signal level5_c7, level5_c8 :  std_logic_vector(56 downto 0);
signal count4_c7, count4_c8, count4_c9, count4_c10 :  std_logic;
signal level4_c8 :  std_logic_vector(56 downto 0);
signal count3_c8, count3_c9, count3_c10 :  std_logic;
signal level3_c8, level3_c9 :  std_logic_vector(56 downto 0);
signal count2_c8, count2_c9, count2_c10 :  std_logic;
signal level2_c9 :  std_logic_vector(56 downto 0);
signal count1_c9, count1_c10 :  std_logic;
signal level1_c9, level1_c10 :  std_logic_vector(56 downto 0);
signal count0_c10 :  std_logic;
signal level0_c10 :  std_logic_vector(56 downto 0);
signal sCount_c10 :  std_logic_vector(5 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_7 = '1' then
               level6_c7 <= level6_c6;
            end if;
            if ce_8 = '1' then
               count5_c8 <= count5_c7;
               level5_c8 <= level5_c7;
               count4_c8 <= count4_c7;
            end if;
            if ce_9 = '1' then
               count5_c9 <= count5_c8;
               count4_c9 <= count4_c8;
               count3_c9 <= count3_c8;
               level3_c9 <= level3_c8;
               count2_c9 <= count2_c8;
            end if;
            if ce_10 = '1' then
               count5_c10 <= count5_c9;
               count4_c10 <= count4_c9;
               count3_c10 <= count3_c9;
               count2_c10 <= count2_c9;
               count1_c10 <= count1_c9;
               level1_c10 <= level1_c9;
            end if;
         end if;
      end process;
   level6_c6 <= X ;
   count5_c7<= '1' when level6_c7(56 downto 25) = (56 downto 25=>'0') else '0';
   level5_c7<= level6_c7(56 downto 0) when count5_c7='0' else level6_c7(24 downto 0) & (31 downto 0 => '0');

   count4_c7<= '1' when level5_c7(56 downto 41) = (56 downto 41=>'0') else '0';
   level4_c8<= level5_c8(56 downto 0) when count4_c8='0' else level5_c8(40 downto 0) & (15 downto 0 => '0');

   count3_c8<= '1' when level4_c8(56 downto 49) = (56 downto 49=>'0') else '0';
   level3_c8<= level4_c8(56 downto 0) when count3_c8='0' else level4_c8(48 downto 0) & (7 downto 0 => '0');

   count2_c8<= '1' when level3_c8(56 downto 53) = (56 downto 53=>'0') else '0';
   level2_c9<= level3_c9(56 downto 0) when count2_c9='0' else level3_c9(52 downto 0) & (3 downto 0 => '0');

   count1_c9<= '1' when level2_c9(56 downto 55) = (56 downto 55=>'0') else '0';
   level1_c9<= level2_c9(56 downto 0) when count1_c9='0' else level2_c9(54 downto 0) & (1 downto 0 => '0');

   count0_c10<= '1' when level1_c10(56 downto 56) = (56 downto 56=>'0') else '0';
   level0_c10<= level1_c10(56 downto 0) when count0_c10='0' else level1_c10(55 downto 0) & (0 downto 0 => '0');

   R <= level0_c10;
   sCount_c10 <= count5_c10 & count4_c10 & count3_c10 & count2_c10 & count1_c10 & count0_c10;
   Count <= sCount_c10;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_66_Freq500_uid11
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 11 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_66_Freq500_uid11 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
          X : in  std_logic_vector(65 downto 0);
          Y : in  std_logic_vector(65 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of IntAdder_66_Freq500_uid11 is
signal Cin_1_c10, Cin_1_c11 :  std_logic;
signal X_1_c10, X_1_c11 :  std_logic_vector(66 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3, Y_1_c4, Y_1_c5, Y_1_c6, Y_1_c7, Y_1_c8, Y_1_c9, Y_1_c10, Y_1_c11 :  std_logic_vector(66 downto 0);
signal S_1_c11 :  std_logic_vector(66 downto 0);
signal R_1_c11 :  std_logic_vector(65 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_1_c1 <= Y_1_c0;
            end if;
            if ce_2 = '1' then
               Y_1_c2 <= Y_1_c1;
            end if;
            if ce_3 = '1' then
               Y_1_c3 <= Y_1_c2;
            end if;
            if ce_4 = '1' then
               Y_1_c4 <= Y_1_c3;
            end if;
            if ce_5 = '1' then
               Y_1_c5 <= Y_1_c4;
            end if;
            if ce_6 = '1' then
               Y_1_c6 <= Y_1_c5;
            end if;
            if ce_7 = '1' then
               Y_1_c7 <= Y_1_c6;
            end if;
            if ce_8 = '1' then
               Y_1_c8 <= Y_1_c7;
            end if;
            if ce_9 = '1' then
               Y_1_c9 <= Y_1_c8;
            end if;
            if ce_10 = '1' then
               Y_1_c10 <= Y_1_c9;
            end if;
            if ce_11 = '1' then
               Cin_1_c11 <= Cin_1_c10;
               X_1_c11 <= X_1_c10;
               Y_1_c11 <= Y_1_c10;
            end if;
         end if;
      end process;
   Cin_1_c10 <= Cin;
   X_1_c10 <= '0' & X(65 downto 0);
   Y_1_c0 <= '0' & Y(65 downto 0);
   S_1_c11 <= X_1_c11 + Y_1_c11 + Cin_1_c11;
   R_1_c11 <= S_1_c11(65 downto 0);
   R <= R_1_c11 ;
end architecture;

--------------------------------------------------------------------------------
--                             FloatingPointAdder
--                         (FPAdd_11_52_Freq500_uid2)
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2010-2017)
--------------------------------------------------------------------------------
-- Pipeline depth: 12 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointAdder_64_2_705000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointAdder_64_2_705000 is
   component RightShifterSticky53_by_max_55_Freq500_uid4 is
      port ( clk, ce_2, ce_3, ce_4, ce_5 : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             S : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(54 downto 0);
             Sticky : out  std_logic   );
   end component;

   component IntAdder_56_Freq500_uid6 is
      port ( clk, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(55 downto 0)   );
   end component;

   component Normalizer_Z_57_57_57_Freq500_uid8 is
      port ( clk, ce_7, ce_8, ce_9, ce_10 : in std_logic;
             X : in  std_logic_vector(56 downto 0);
             Count : out  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(56 downto 0)   );
   end component;

   component IntAdder_66_Freq500_uid11 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11 : in std_logic;
             X : in  std_logic_vector(65 downto 0);
             Y : in  std_logic_vector(65 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(65 downto 0)   );
   end component;

signal excExpFracX_c0 :  std_logic_vector(64 downto 0);
signal excExpFracY_c0 :  std_logic_vector(64 downto 0);
signal swap_c0, swap_c1 :  std_logic;
signal eXmeY_c0, eXmeY_c1 :  std_logic_vector(10 downto 0);
signal eYmeX_c0, eYmeX_c1 :  std_logic_vector(10 downto 0);
signal expDiff_c1 :  std_logic_vector(10 downto 0);
signal newX_c1 :  std_logic_vector(65 downto 0);
signal newY_c1 :  std_logic_vector(65 downto 0);
signal expX_c1 :  std_logic_vector(10 downto 0);
signal excX_c1 :  std_logic_vector(1 downto 0);
signal excY_c1 :  std_logic_vector(1 downto 0);
signal signX_c1 :  std_logic;
signal signY_c1 :  std_logic;
signal EffSub_c1, EffSub_c2, EffSub_c3, EffSub_c4, EffSub_c5, EffSub_c6, EffSub_c7, EffSub_c8, EffSub_c9, EffSub_c10, EffSub_c11, EffSub_c12 :  std_logic;
signal sXsYExnXY_c1 :  std_logic_vector(5 downto 0);
signal sdExnXY_c1 :  std_logic_vector(3 downto 0);
signal fracY_c1 :  std_logic_vector(52 downto 0);
signal excRt_c1, excRt_c2, excRt_c3, excRt_c4, excRt_c5, excRt_c6, excRt_c7, excRt_c8, excRt_c9, excRt_c10, excRt_c11, excRt_c12 :  std_logic_vector(1 downto 0);
signal signR_c1, signR_c2, signR_c3, signR_c4, signR_c5, signR_c6, signR_c7, signR_c8, signR_c9, signR_c10 :  std_logic;
signal shiftedOut_c1 :  std_logic;
signal shiftVal_c1 :  std_logic_vector(5 downto 0);
signal shiftedFracY_c2 :  std_logic_vector(54 downto 0);
signal sticky_c5, sticky_c6 :  std_logic;
signal fracYpad_c2 :  std_logic_vector(55 downto 0);
signal EffSubVector_c1, EffSubVector_c2 :  std_logic_vector(55 downto 0);
signal fracYpadXorOp_c2 :  std_logic_vector(55 downto 0);
signal fracXpad_c1 :  std_logic_vector(55 downto 0);
signal cInSigAdd_c5 :  std_logic;
signal fracAddResult_c6 :  std_logic_vector(55 downto 0);
signal fracSticky_c6 :  std_logic_vector(56 downto 0);
signal nZerosNew_c10 :  std_logic_vector(5 downto 0);
signal shiftedFrac_c10 :  std_logic_vector(56 downto 0);
signal extendedExpInc_c1, extendedExpInc_c2, extendedExpInc_c3, extendedExpInc_c4, extendedExpInc_c5, extendedExpInc_c6, extendedExpInc_c7, extendedExpInc_c8, extendedExpInc_c9, extendedExpInc_c10 :  std_logic_vector(11 downto 0);
signal updatedExp_c10 :  std_logic_vector(12 downto 0);
signal eqdiffsign_c10, eqdiffsign_c11, eqdiffsign_c12 :  std_logic;
signal expFrac_c10 :  std_logic_vector(65 downto 0);
signal stk_c10 :  std_logic;
signal rnd_c10 :  std_logic;
signal lsb_c10 :  std_logic;
signal needToRound_c10 :  std_logic;
signal RoundedExpFrac_c11 :  std_logic_vector(65 downto 0);
signal upExc_c11 :  std_logic_vector(1 downto 0);
signal fracR_c11, fracR_c12 :  std_logic_vector(51 downto 0);
signal expR_c11, expR_c12 :  std_logic_vector(10 downto 0);
signal exExpExc_c11, exExpExc_c12 :  std_logic_vector(3 downto 0);
signal excRt2_c12 :  std_logic_vector(1 downto 0);
signal excR_c12 :  std_logic_vector(1 downto 0);
signal signR2_c10, signR2_c11, signR2_c12 :  std_logic;
signal computedR_c12 :  std_logic_vector(65 downto 0);
signal X_c1 :  std_logic_vector(11+52+2 downto 0);
signal Y_c1 :  std_logic_vector(11+52+2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               swap_c1 <= swap_c0;
               eXmeY_c1 <= eXmeY_c0;
               eYmeX_c1 <= eYmeX_c0;
               X_c1 <= X;
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               EffSub_c2 <= EffSub_c1;
               excRt_c2 <= excRt_c1;
               signR_c2 <= signR_c1;
               EffSubVector_c2 <= EffSubVector_c1;
               extendedExpInc_c2 <= extendedExpInc_c1;
            end if;
            if ce_3 = '1' then
               EffSub_c3 <= EffSub_c2;
               excRt_c3 <= excRt_c2;
               signR_c3 <= signR_c2;
               extendedExpInc_c3 <= extendedExpInc_c2;
            end if;
            if ce_4 = '1' then
               EffSub_c4 <= EffSub_c3;
               excRt_c4 <= excRt_c3;
               signR_c4 <= signR_c3;
               extendedExpInc_c4 <= extendedExpInc_c3;
            end if;
            if ce_5 = '1' then
               EffSub_c5 <= EffSub_c4;
               excRt_c5 <= excRt_c4;
               signR_c5 <= signR_c4;
               extendedExpInc_c5 <= extendedExpInc_c4;
            end if;
            if ce_6 = '1' then
               EffSub_c6 <= EffSub_c5;
               excRt_c6 <= excRt_c5;
               signR_c6 <= signR_c5;
               sticky_c6 <= sticky_c5;
               extendedExpInc_c6 <= extendedExpInc_c5;
            end if;
            if ce_7 = '1' then
               EffSub_c7 <= EffSub_c6;
               excRt_c7 <= excRt_c6;
               signR_c7 <= signR_c6;
               extendedExpInc_c7 <= extendedExpInc_c6;
            end if;
            if ce_8 = '1' then
               EffSub_c8 <= EffSub_c7;
               excRt_c8 <= excRt_c7;
               signR_c8 <= signR_c7;
               extendedExpInc_c8 <= extendedExpInc_c7;
            end if;
            if ce_9 = '1' then
               EffSub_c9 <= EffSub_c8;
               excRt_c9 <= excRt_c8;
               signR_c9 <= signR_c8;
               extendedExpInc_c9 <= extendedExpInc_c8;
            end if;
            if ce_10 = '1' then
               EffSub_c10 <= EffSub_c9;
               excRt_c10 <= excRt_c9;
               signR_c10 <= signR_c9;
               extendedExpInc_c10 <= extendedExpInc_c9;
            end if;
            if ce_11 = '1' then
               EffSub_c11 <= EffSub_c10;
               excRt_c11 <= excRt_c10;
               eqdiffsign_c11 <= eqdiffsign_c10;
               signR2_c11 <= signR2_c10;
            end if;
            if ce_12 = '1' then
               EffSub_c12 <= EffSub_c11;
               excRt_c12 <= excRt_c11;
               eqdiffsign_c12 <= eqdiffsign_c11;
               fracR_c12 <= fracR_c11;
               expR_c12 <= expR_c11;
               exExpExc_c12 <= exExpExc_c11;
               signR2_c12 <= signR2_c11;
            end if;
         end if;
      end process;
   excExpFracX_c0 <= X(65 downto 64) & X(62 downto 0);
   excExpFracY_c0 <= Y(65 downto 64) & Y(62 downto 0);
   swap_c0 <= '1' when excExpFracX_c0 < excExpFracY_c0 else '0';
   -- exponent difference
   eXmeY_c0 <= (X(62 downto 52)) - (Y(62 downto 52));
   eYmeX_c0 <= (Y(62 downto 52)) - (X(62 downto 52));
   expDiff_c1 <= eXmeY_c1 when swap_c1 = '0' else eYmeX_c1;
   -- input swap so that |X|>|Y|
   newX_c1 <= X_c1 when swap_c1 = '0' else Y_c1;
   newY_c1 <= Y_c1 when swap_c1 = '0' else X_c1;
   -- now we decompose the inputs into their sign, exponent, fraction
   expX_c1<= newX_c1(62 downto 52);
   excX_c1<= newX_c1(65 downto 64);
   excY_c1<= newY_c1(65 downto 64);
   signX_c1<= newX_c1(63);
   signY_c1<= newY_c1(63);
   EffSub_c1 <= signX_c1 xor signY_c1;
   sXsYExnXY_c1 <= signX_c1 & signY_c1 & excX_c1 & excY_c1;
   sdExnXY_c1 <= excX_c1 & excY_c1;
   fracY_c1 <= "00000000000000000000000000000000000000000000000000000" when excY_c1="00" else ('1' & newY_c1(51 downto 0));
   -- Exception management logic
   with sXsYExnXY_c1  select  
   excRt_c1 <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR_c1<= '0' when (sXsYExnXY_c1="100000" or sXsYExnXY_c1="010000") else signX_c1;
   shiftedOut_c1 <= '1' when (expDiff_c1 > 54) else '0';
   shiftVal_c1 <= expDiff_c1(5 downto 0) when shiftedOut_c1='0' else CONV_STD_LOGIC_VECTOR(55,6);
   RightShifterComponent: RightShifterSticky53_by_max_55_Freq500_uid4
      port map ( clk  => clk,
                 ce_2 => ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 S => shiftVal_c1,
                 X => fracY_c1,
                 R => shiftedFracY_c2,
                 Sticky => sticky_c5);
   fracYpad_c2 <= "0" & shiftedFracY_c2;
   EffSubVector_c1 <= (55 downto 0 => EffSub_c1);
   fracYpadXorOp_c2 <= fracYpad_c2 xor EffSubVector_c2;
   fracXpad_c1 <= "01" & (newX_c1(51 downto 0)) & "00";
   cInSigAdd_c5 <= EffSub_c5 and not sticky_c5; -- if we subtract and the sticky was one, some of the negated sticky bits would have absorbed this carry 
   fracAdder: IntAdder_56_Freq500_uid6
      port map ( clk  => clk,
                 ce_2 => ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 Cin => cInSigAdd_c5,
                 X => fracXpad_c1,
                 Y => fracYpadXorOp_c2,
                 R => fracAddResult_c6);
   fracSticky_c6<= fracAddResult_c6 & sticky_c6; 
   LZCAndShifter: Normalizer_Z_57_57_57_Freq500_uid8
      port map ( clk  => clk,
                 ce_7 => ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 X => fracSticky_c6,
                 Count => nZerosNew_c10,
                 R => shiftedFrac_c10);
   extendedExpInc_c1<= ("0" & expX_c1) + '1';
   updatedExp_c10 <= ("0" &extendedExpInc_c10) - ("0000000" & nZerosNew_c10);
   eqdiffsign_c10 <= '1' when nZerosNew_c10="111111" else '0';
   expFrac_c10<= updatedExp_c10 & shiftedFrac_c10(55 downto 3);
   stk_c10<= shiftedFrac_c10(2) or shiftedFrac_c10(1) or shiftedFrac_c10(0);
   rnd_c10<= shiftedFrac_c10(3);
   lsb_c10<= shiftedFrac_c10(4);
   needToRound_c10<= '1' when (rnd_c10='1' and stk_c10='1') or (rnd_c10='1' and stk_c10='0' and lsb_c10='1')
  else '0';
   roundingAdder: IntAdder_66_Freq500_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 Cin => needToRound_c10,
                 X => expFrac_c10,
                 Y => "000000000000000000000000000000000000000000000000000000000000000000",
                 R => RoundedExpFrac_c11);
   -- possible update to exception bits
   upExc_c11 <= RoundedExpFrac_c11(65 downto 64);
   fracR_c11 <= RoundedExpFrac_c11(52 downto 1);
   expR_c11 <= RoundedExpFrac_c11(63 downto 53);
   exExpExc_c11 <= upExc_c11 & excRt_c11;
   with exExpExc_c12  select  
   excRt2_c12<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR_c12 <= "00" when (eqdiffsign_c12='1' and EffSub_c12='1'  and not(excRt_c12="11")) else excRt2_c12;
   signR2_c10 <= '0' when (eqdiffsign_c10='1' and EffSub_c10='1') else signR_c10;
   computedR_c12 <= excR_c12 & signR2_c12 & expR_c12 & fracR_c12;
   R <= computedR_c12;
end architecture;




--------------------------------------------------------------------------------
--                RightShifterSticky53_by_max_55_Freq300_uid4
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X S
-- Output signals: R Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifterSticky53_by_max_55_Freq300_uid4 is
    port (clk, ce_1, ce_2, ce_3 : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          S : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(54 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of RightShifterSticky53_by_max_55_Freq300_uid4 is
signal ps_c0, ps_c1, ps_c2, ps_c3 :  std_logic_vector(5 downto 0);
signal Xpadded_c0 :  std_logic_vector(54 downto 0);
signal level6_c0, level6_c1 :  std_logic_vector(54 downto 0);
signal stk5_c1 :  std_logic;
signal level5_c0, level5_c1 :  std_logic_vector(54 downto 0);
signal stk4_c1, stk4_c2 :  std_logic;
signal level4_c1, level4_c2 :  std_logic_vector(54 downto 0);
signal stk3_c2 :  std_logic;
signal level3_c1, level3_c2 :  std_logic_vector(54 downto 0);
signal stk2_c2 :  std_logic;
signal level2_c1, level2_c2 :  std_logic_vector(54 downto 0);
signal stk1_c2, stk1_c3 :  std_logic;
signal level1_c1, level1_c2, level1_c3 :  std_logic_vector(54 downto 0);
signal stk0_c3 :  std_logic;
signal level0_c1 :  std_logic_vector(54 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               ps_c1 <= ps_c0;
               level6_c1 <= level6_c0;
               level5_c1 <= level5_c0;
            end if;
            if ce_2 = '1' then
               ps_c2 <= ps_c1;
               stk4_c2 <= stk4_c1;
               level4_c2 <= level4_c1;
               level3_c2 <= level3_c1;
               level2_c2 <= level2_c1;
               level1_c2 <= level1_c1;
            end if;
            if ce_3 = '1' then
               ps_c3 <= ps_c2;
               stk1_c3 <= stk1_c2;
               level1_c3 <= level1_c2;
            end if;
         end if;
      end process;
   ps_c0<= S;
   Xpadded_c0 <= X&(1 downto 0 => '0');
   level6_c0<= Xpadded_c0;
   stk5_c1 <= '1' when (level6_c1(31 downto 0)/="00000000000000000000000000000000" and ps_c1(5)='1')   else '0';
   level5_c0 <=  level6_c0 when  ps_c0(5)='0'    else (31 downto 0 => '0') & level6_c0(54 downto 32);
   stk4_c1 <= '1' when (level5_c1(15 downto 0)/="0000000000000000" and ps_c1(4)='1') or stk5_c1 ='1'   else '0';
   level4_c1 <=  level5_c1 when  ps_c1(4)='0'    else (15 downto 0 => '0') & level5_c1(54 downto 16);
   stk3_c2 <= '1' when (level4_c2(7 downto 0)/="00000000" and ps_c2(3)='1') or stk4_c2 ='1'   else '0';
   level3_c1 <=  level4_c1 when  ps_c1(3)='0'    else (7 downto 0 => '0') & level4_c1(54 downto 8);
   stk2_c2 <= '1' when (level3_c2(3 downto 0)/="0000" and ps_c2(2)='1') or stk3_c2 ='1'   else '0';
   level2_c1 <=  level3_c1 when  ps_c1(2)='0'    else (3 downto 0 => '0') & level3_c1(54 downto 4);
   stk1_c2 <= '1' when (level2_c2(1 downto 0)/="00" and ps_c2(1)='1') or stk2_c2 ='1'   else '0';
   level1_c1 <=  level2_c1 when  ps_c1(1)='0'    else (1 downto 0 => '0') & level2_c1(54 downto 2);
   stk0_c3 <= '1' when (level1_c3(0 downto 0)/="0" and ps_c3(0)='1') or stk1_c3 ='1'   else '0';
   level0_c1 <=  level1_c1 when  ps_c1(0)='0'    else (0 downto 0 => '0') & level1_c1(54 downto 1);
   R <= level0_c1;
   Sticky <= stk0_c3;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_56_Freq300_uid6
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_56_Freq300_uid6 is
    port (clk, ce_1, ce_2, ce_3 : in std_logic;
          X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntAdder_56_Freq300_uid6 is
signal Rtmp_c3 :  std_logic_vector(55 downto 0);
signal X_c1, X_c2, X_c3 :  std_logic_vector(55 downto 0);
signal Y_c2, Y_c3 :  std_logic_vector(55 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               X_c1 <= X;
            end if;
            if ce_2 = '1' then
               X_c2 <= X_c1;
               Y_c2 <= Y;
            end if;
            if ce_3 = '1' then
               X_c3 <= X_c2;
               Y_c3 <= Y_c2;
            end if;
         end if;
      end process;
   Rtmp_c3 <= X_c3 + Y_c3 + Cin;
   R <= Rtmp_c3;
end architecture;

--------------------------------------------------------------------------------
--                     Normalizer_Z_57_57_57_Freq300_uid8
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_57_57_57_Freq300_uid8 is
    port (clk, ce_4, ce_5 : in std_logic;
          X : in  std_logic_vector(56 downto 0);
          Count : out  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of Normalizer_Z_57_57_57_Freq300_uid8 is
signal level6_c3, level6_c4 :  std_logic_vector(56 downto 0);
signal count5_c4, count5_c5 :  std_logic;
signal level5_c4 :  std_logic_vector(56 downto 0);
signal count4_c4, count4_c5 :  std_logic;
signal level4_c4 :  std_logic_vector(56 downto 0);
signal count3_c4, count3_c5 :  std_logic;
signal level3_c4, level3_c5 :  std_logic_vector(56 downto 0);
signal count2_c5 :  std_logic;
signal level2_c5 :  std_logic_vector(56 downto 0);
signal count1_c5 :  std_logic;
signal level1_c5 :  std_logic_vector(56 downto 0);
signal count0_c5 :  std_logic;
signal level0_c5 :  std_logic_vector(56 downto 0);
signal sCount_c5 :  std_logic_vector(5 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_4 = '1' then
               level6_c4 <= level6_c3;
            end if;
            if ce_5 = '1' then
               count5_c5 <= count5_c4;
               count4_c5 <= count4_c4;
               count3_c5 <= count3_c4;
               level3_c5 <= level3_c4;
            end if;
         end if;
      end process;
   level6_c3 <= X ;
   count5_c4<= '1' when level6_c4(56 downto 25) = (56 downto 25=>'0') else '0';
   level5_c4<= level6_c4(56 downto 0) when count5_c4='0' else level6_c4(24 downto 0) & (31 downto 0 => '0');

   count4_c4<= '1' when level5_c4(56 downto 41) = (56 downto 41=>'0') else '0';
   level4_c4<= level5_c4(56 downto 0) when count4_c4='0' else level5_c4(40 downto 0) & (15 downto 0 => '0');

   count3_c4<= '1' when level4_c4(56 downto 49) = (56 downto 49=>'0') else '0';
   level3_c4<= level4_c4(56 downto 0) when count3_c4='0' else level4_c4(48 downto 0) & (7 downto 0 => '0');

   count2_c5<= '1' when level3_c5(56 downto 53) = (56 downto 53=>'0') else '0';
   level2_c5<= level3_c5(56 downto 0) when count2_c5='0' else level3_c5(52 downto 0) & (3 downto 0 => '0');

   count1_c5<= '1' when level2_c5(56 downto 55) = (56 downto 55=>'0') else '0';
   level1_c5<= level2_c5(56 downto 0) when count1_c5='0' else level2_c5(54 downto 0) & (1 downto 0 => '0');

   count0_c5<= '1' when level1_c5(56 downto 56) = (56 downto 56=>'0') else '0';
   level0_c5<= level1_c5(56 downto 0) when count0_c5='0' else level1_c5(55 downto 0) & (0 downto 0 => '0');

   R <= level0_c5;
   sCount_c5 <= count5_c5 & count4_c5 & count3_c5 & count2_c5 & count1_c5 & count0_c5;
   Count <= sCount_c5;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_66_Freq300_uid11
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_66_Freq300_uid11 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(65 downto 0);
          Y : in  std_logic_vector(65 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of IntAdder_66_Freq300_uid11 is
signal Rtmp_c6 :  std_logic_vector(65 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6 :  std_logic_vector(65 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
         end if;
      end process;
   Rtmp_c6 <= X + Y_c6 + Cin;
   R <= Rtmp_c6;
end architecture;

--------------------------------------------------------------------------------
--                             FloatingPointAdder
--                         (FPAdd_11_52_Freq300_uid2)
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2010-2017)
--------------------------------------------------------------------------------
-- Pipeline depth: 7 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointAdder_64_5_091333 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointAdder_64_5_091333 is
   component RightShifterSticky53_by_max_55_Freq300_uid4 is
      port ( clk, ce_1, ce_2, ce_3 : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             S : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(54 downto 0);
             Sticky : out  std_logic   );
   end component;

   component IntAdder_56_Freq300_uid6 is
      port ( clk, ce_1, ce_2, ce_3 : in std_logic;
             X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(55 downto 0)   );
   end component;

   component Normalizer_Z_57_57_57_Freq300_uid8 is
      port ( clk, ce_4, ce_5 : in std_logic;
             X : in  std_logic_vector(56 downto 0);
             Count : out  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(56 downto 0)   );
   end component;

   component IntAdder_66_Freq300_uid11 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(65 downto 0);
             Y : in  std_logic_vector(65 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(65 downto 0)   );
   end component;

signal excExpFracX_c0 :  std_logic_vector(64 downto 0);
signal excExpFracY_c0 :  std_logic_vector(64 downto 0);
signal swap_c0 :  std_logic;
signal eXmeY_c0 :  std_logic_vector(10 downto 0);
signal eYmeX_c0 :  std_logic_vector(10 downto 0);
signal expDiff_c0 :  std_logic_vector(10 downto 0);
signal newX_c0 :  std_logic_vector(65 downto 0);
signal newY_c0 :  std_logic_vector(65 downto 0);
signal expX_c0 :  std_logic_vector(10 downto 0);
signal excX_c0 :  std_logic_vector(1 downto 0);
signal excY_c0 :  std_logic_vector(1 downto 0);
signal signX_c0 :  std_logic;
signal signY_c0 :  std_logic;
signal EffSub_c0, EffSub_c1, EffSub_c2, EffSub_c3, EffSub_c4, EffSub_c5, EffSub_c6, EffSub_c7 :  std_logic;
signal sXsYExnXY_c0 :  std_logic_vector(5 downto 0);
signal sdExnXY_c0 :  std_logic_vector(3 downto 0);
signal fracY_c0 :  std_logic_vector(52 downto 0);
signal excRt_c0, excRt_c1, excRt_c2, excRt_c3, excRt_c4, excRt_c5, excRt_c6, excRt_c7 :  std_logic_vector(1 downto 0);
signal signR_c0, signR_c1, signR_c2, signR_c3, signR_c4, signR_c5 :  std_logic;
signal shiftedOut_c0 :  std_logic;
signal shiftVal_c0 :  std_logic_vector(5 downto 0);
signal shiftedFracY_c1 :  std_logic_vector(54 downto 0);
signal sticky_c3 :  std_logic;
signal fracYpad_c1 :  std_logic_vector(55 downto 0);
signal EffSubVector_c0, EffSubVector_c1 :  std_logic_vector(55 downto 0);
signal fracYpadXorOp_c1 :  std_logic_vector(55 downto 0);
signal fracXpad_c0 :  std_logic_vector(55 downto 0);
signal cInSigAdd_c3 :  std_logic;
signal fracAddResult_c3 :  std_logic_vector(55 downto 0);
signal fracSticky_c3 :  std_logic_vector(56 downto 0);
signal nZerosNew_c5, nZerosNew_c6 :  std_logic_vector(5 downto 0);
signal shiftedFrac_c5, shiftedFrac_c6 :  std_logic_vector(56 downto 0);
signal extendedExpInc_c0, extendedExpInc_c1, extendedExpInc_c2, extendedExpInc_c3, extendedExpInc_c4, extendedExpInc_c5, extendedExpInc_c6 :  std_logic_vector(11 downto 0);
signal updatedExp_c6 :  std_logic_vector(12 downto 0);
signal eqdiffsign_c5, eqdiffsign_c6, eqdiffsign_c7 :  std_logic;
signal expFrac_c6 :  std_logic_vector(65 downto 0);
signal stk_c5, stk_c6 :  std_logic;
signal rnd_c5, rnd_c6 :  std_logic;
signal lsb_c5, lsb_c6 :  std_logic;
signal needToRound_c6 :  std_logic;
signal RoundedExpFrac_c6 :  std_logic_vector(65 downto 0);
signal upExc_c6 :  std_logic_vector(1 downto 0);
signal fracR_c6, fracR_c7 :  std_logic_vector(51 downto 0);
signal expR_c6, expR_c7 :  std_logic_vector(10 downto 0);
signal exExpExc_c6 :  std_logic_vector(3 downto 0);
signal excRt2_c6, excRt2_c7 :  std_logic_vector(1 downto 0);
signal excR_c7 :  std_logic_vector(1 downto 0);
signal signR2_c5, signR2_c6, signR2_c7 :  std_logic;
signal computedR_c7 :  std_logic_vector(65 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               EffSub_c1 <= EffSub_c0;
               excRt_c1 <= excRt_c0;
               signR_c1 <= signR_c0;
               EffSubVector_c1 <= EffSubVector_c0;
               extendedExpInc_c1 <= extendedExpInc_c0;
            end if;
            if ce_2 = '1' then
               EffSub_c2 <= EffSub_c1;
               excRt_c2 <= excRt_c1;
               signR_c2 <= signR_c1;
               extendedExpInc_c2 <= extendedExpInc_c1;
            end if;
            if ce_3 = '1' then
               EffSub_c3 <= EffSub_c2;
               excRt_c3 <= excRt_c2;
               signR_c3 <= signR_c2;
               extendedExpInc_c3 <= extendedExpInc_c2;
            end if;
            if ce_4 = '1' then
               EffSub_c4 <= EffSub_c3;
               excRt_c4 <= excRt_c3;
               signR_c4 <= signR_c3;
               extendedExpInc_c4 <= extendedExpInc_c3;
            end if;
            if ce_5 = '1' then
               EffSub_c5 <= EffSub_c4;
               excRt_c5 <= excRt_c4;
               signR_c5 <= signR_c4;
               extendedExpInc_c5 <= extendedExpInc_c4;
            end if;
            if ce_6 = '1' then
               EffSub_c6 <= EffSub_c5;
               excRt_c6 <= excRt_c5;
               nZerosNew_c6 <= nZerosNew_c5;
               shiftedFrac_c6 <= shiftedFrac_c5;
               extendedExpInc_c6 <= extendedExpInc_c5;
               eqdiffsign_c6 <= eqdiffsign_c5;
               stk_c6 <= stk_c5;
               rnd_c6 <= rnd_c5;
               lsb_c6 <= lsb_c5;
               signR2_c6 <= signR2_c5;
            end if;
            if ce_7 = '1' then
               EffSub_c7 <= EffSub_c6;
               excRt_c7 <= excRt_c6;
               eqdiffsign_c7 <= eqdiffsign_c6;
               fracR_c7 <= fracR_c6;
               expR_c7 <= expR_c6;
               excRt2_c7 <= excRt2_c6;
               signR2_c7 <= signR2_c6;
            end if;
         end if;
      end process;
   excExpFracX_c0 <= X(65 downto 64) & X(62 downto 0);
   excExpFracY_c0 <= Y(65 downto 64) & Y(62 downto 0);
   swap_c0 <= '1' when excExpFracX_c0 < excExpFracY_c0 else '0';
   -- exponent difference
   eXmeY_c0 <= (X(62 downto 52)) - (Y(62 downto 52));
   eYmeX_c0 <= (Y(62 downto 52)) - (X(62 downto 52));
   expDiff_c0 <= eXmeY_c0 when swap_c0 = '0' else eYmeX_c0;
   -- input swap so that |X|>|Y|
   newX_c0 <= X when swap_c0 = '0' else Y;
   newY_c0 <= Y when swap_c0 = '0' else X;
   -- now we decompose the inputs into their sign, exponent, fraction
   expX_c0<= newX_c0(62 downto 52);
   excX_c0<= newX_c0(65 downto 64);
   excY_c0<= newY_c0(65 downto 64);
   signX_c0<= newX_c0(63);
   signY_c0<= newY_c0(63);
   EffSub_c0 <= signX_c0 xor signY_c0;
   sXsYExnXY_c0 <= signX_c0 & signY_c0 & excX_c0 & excY_c0;
   sdExnXY_c0 <= excX_c0 & excY_c0;
   fracY_c0 <= "00000000000000000000000000000000000000000000000000000" when excY_c0="00" else ('1' & newY_c0(51 downto 0));
   -- Exception management logic
   with sXsYExnXY_c0  select  
   excRt_c0 <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR_c0<= '0' when (sXsYExnXY_c0="100000" or sXsYExnXY_c0="010000") else signX_c0;
   shiftedOut_c0 <= '1' when (expDiff_c0 > 54) else '0';
   shiftVal_c0 <= expDiff_c0(5 downto 0) when shiftedOut_c0='0' else CONV_STD_LOGIC_VECTOR(55,6);
   RightShifterComponent: RightShifterSticky53_by_max_55_Freq300_uid4
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 S => shiftVal_c0,
                 X => fracY_c0,
                 R => shiftedFracY_c1,
                 Sticky => sticky_c3);
   fracYpad_c1 <= "0" & shiftedFracY_c1;
   EffSubVector_c0 <= (55 downto 0 => EffSub_c0);
   fracYpadXorOp_c1 <= fracYpad_c1 xor EffSubVector_c1;
   fracXpad_c0 <= "01" & (newX_c0(51 downto 0)) & "00";
   cInSigAdd_c3 <= EffSub_c3 and not sticky_c3; -- if we subtract and the sticky was one, some of the negated sticky bits would have absorbed this carry 
   fracAdder: IntAdder_56_Freq300_uid6
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 Cin => cInSigAdd_c3,
                 X => fracXpad_c0,
                 Y => fracYpadXorOp_c1,
                 R => fracAddResult_c3);
   fracSticky_c3<= fracAddResult_c3 & sticky_c3; 
   LZCAndShifter: Normalizer_Z_57_57_57_Freq300_uid8
      port map ( clk  => clk,
                 ce_4 => ce_4,
                 ce_5=> ce_5,
                 X => fracSticky_c3,
                 Count => nZerosNew_c5,
                 R => shiftedFrac_c5);
   extendedExpInc_c0<= ("0" & expX_c0) + '1';
   updatedExp_c6 <= ("0" &extendedExpInc_c6) - ("0000000" & nZerosNew_c6);
   eqdiffsign_c5 <= '1' when nZerosNew_c5="111111" else '0';
   expFrac_c6<= updatedExp_c6 & shiftedFrac_c6(55 downto 3);
   stk_c5<= shiftedFrac_c5(2) or shiftedFrac_c5(1) or shiftedFrac_c5(0);
   rnd_c5<= shiftedFrac_c5(3);
   lsb_c5<= shiftedFrac_c5(4);
   needToRound_c6<= '1' when (rnd_c6='1' and stk_c6='1') or (rnd_c6='1' and stk_c6='0' and lsb_c6='1')
  else '0';
   roundingAdder: IntAdder_66_Freq300_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 Cin => needToRound_c6,
                 X => expFrac_c6,
                 Y => "000000000000000000000000000000000000000000000000000000000000000000",
                 R => RoundedExpFrac_c6);
   -- possible update to exception bits
   upExc_c6 <= RoundedExpFrac_c6(65 downto 64);
   fracR_c6 <= RoundedExpFrac_c6(52 downto 1);
   expR_c6 <= RoundedExpFrac_c6(63 downto 53);
   exExpExc_c6 <= upExc_c6 & excRt_c6;
   with exExpExc_c6  select  
   excRt2_c6<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR_c7 <= "00" when (eqdiffsign_c7='1' and EffSub_c7='1'  and not(excRt_c7="11")) else excRt2_c7;
   signR2_c5 <= '0' when (eqdiffsign_c5='1' and EffSub_c5='1') else signR_c5;
   computedR_c7 <= excR_c7 & signR2_c7 & expR_c7 & fracR_c7;
   R <= computedR_c7;
end architecture;




--------------------------------------------------------------------------------
--                RightShifterSticky53_by_max_55_Freq100_uid4
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X S
-- Output signals: R Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifterSticky53_by_max_55_Freq100_uid4 is
    port (clk : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          S : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(54 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of RightShifterSticky53_by_max_55_Freq100_uid4 is
signal ps_c0 :  std_logic_vector(5 downto 0);
signal Xpadded_c0 :  std_logic_vector(54 downto 0);
signal level6_c0 :  std_logic_vector(54 downto 0);
signal stk5_c0 :  std_logic;
signal level5_c0 :  std_logic_vector(54 downto 0);
signal stk4_c0 :  std_logic;
signal level4_c0 :  std_logic_vector(54 downto 0);
signal stk3_c0 :  std_logic;
signal level3_c0 :  std_logic_vector(54 downto 0);
signal stk2_c0 :  std_logic;
signal level2_c0 :  std_logic_vector(54 downto 0);
signal stk1_c0 :  std_logic;
signal level1_c0 :  std_logic_vector(54 downto 0);
signal stk0_c0 :  std_logic;
signal level0_c0 :  std_logic_vector(54 downto 0);
begin
   ps_c0<= S;
   Xpadded_c0 <= X&(1 downto 0 => '0');
   level6_c0<= Xpadded_c0;
   stk5_c0 <= '1' when (level6_c0(31 downto 0)/="00000000000000000000000000000000" and ps_c0(5)='1')   else '0';
   level5_c0 <=  level6_c0 when  ps_c0(5)='0'    else (31 downto 0 => '0') & level6_c0(54 downto 32);
   stk4_c0 <= '1' when (level5_c0(15 downto 0)/="0000000000000000" and ps_c0(4)='1') or stk5_c0 ='1'   else '0';
   level4_c0 <=  level5_c0 when  ps_c0(4)='0'    else (15 downto 0 => '0') & level5_c0(54 downto 16);
   stk3_c0 <= '1' when (level4_c0(7 downto 0)/="00000000" and ps_c0(3)='1') or stk4_c0 ='1'   else '0';
   level3_c0 <=  level4_c0 when  ps_c0(3)='0'    else (7 downto 0 => '0') & level4_c0(54 downto 8);
   stk2_c0 <= '1' when (level3_c0(3 downto 0)/="0000" and ps_c0(2)='1') or stk3_c0 ='1'   else '0';
   level2_c0 <=  level3_c0 when  ps_c0(2)='0'    else (3 downto 0 => '0') & level3_c0(54 downto 4);
   stk1_c0 <= '1' when (level2_c0(1 downto 0)/="00" and ps_c0(1)='1') or stk2_c0 ='1'   else '0';
   level1_c0 <=  level2_c0 when  ps_c0(1)='0'    else (1 downto 0 => '0') & level2_c0(54 downto 2);
   stk0_c0 <= '1' when (level1_c0(0 downto 0)/="0" and ps_c0(0)='1') or stk1_c0 ='1'   else '0';
   level0_c0 <=  level1_c0 when  ps_c0(0)='0'    else (0 downto 0 => '0') & level1_c0(54 downto 1);
   R <= level0_c0;
   Sticky <= stk0_c0;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_56_Freq100_uid6
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_56_Freq100_uid6 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntAdder_56_Freq100_uid6 is
signal Rtmp_c1 :  std_logic_vector(55 downto 0);
signal X_c1 :  std_logic_vector(55 downto 0);
signal Y_c1 :  std_logic_vector(55 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               X_c1 <= X;
               Y_c1 <= Y;
            end if;
         end if;
      end process;
   Rtmp_c1 <= X_c1 + Y_c1 + Cin;
   R <= Rtmp_c1;
end architecture;

--------------------------------------------------------------------------------
--                     Normalizer_Z_57_57_57_Freq100_uid8
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_57_57_57_Freq100_uid8 is
    port (clk : in std_logic;
          X : in  std_logic_vector(56 downto 0);
          Count : out  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(56 downto 0)   );
end entity;

architecture arch of Normalizer_Z_57_57_57_Freq100_uid8 is
signal level6_c1 :  std_logic_vector(56 downto 0);
signal count5_c1 :  std_logic;
signal level5_c1 :  std_logic_vector(56 downto 0);
signal count4_c1 :  std_logic;
signal level4_c1 :  std_logic_vector(56 downto 0);
signal count3_c1 :  std_logic;
signal level3_c1 :  std_logic_vector(56 downto 0);
signal count2_c1 :  std_logic;
signal level2_c1 :  std_logic_vector(56 downto 0);
signal count1_c1 :  std_logic;
signal level1_c1 :  std_logic_vector(56 downto 0);
signal count0_c1 :  std_logic;
signal level0_c1 :  std_logic_vector(56 downto 0);
signal sCount_c1 :  std_logic_vector(5 downto 0);
begin
   level6_c1 <= X ;
   count5_c1<= '1' when level6_c1(56 downto 25) = (56 downto 25=>'0') else '0';
   level5_c1<= level6_c1(56 downto 0) when count5_c1='0' else level6_c1(24 downto 0) & (31 downto 0 => '0');

   count4_c1<= '1' when level5_c1(56 downto 41) = (56 downto 41=>'0') else '0';
   level4_c1<= level5_c1(56 downto 0) when count4_c1='0' else level5_c1(40 downto 0) & (15 downto 0 => '0');

   count3_c1<= '1' when level4_c1(56 downto 49) = (56 downto 49=>'0') else '0';
   level3_c1<= level4_c1(56 downto 0) when count3_c1='0' else level4_c1(48 downto 0) & (7 downto 0 => '0');

   count2_c1<= '1' when level3_c1(56 downto 53) = (56 downto 53=>'0') else '0';
   level2_c1<= level3_c1(56 downto 0) when count2_c1='0' else level3_c1(52 downto 0) & (3 downto 0 => '0');

   count1_c1<= '1' when level2_c1(56 downto 55) = (56 downto 55=>'0') else '0';
   level1_c1<= level2_c1(56 downto 0) when count1_c1='0' else level2_c1(54 downto 0) & (1 downto 0 => '0');

   count0_c1<= '1' when level1_c1(56 downto 56) = (56 downto 56=>'0') else '0';
   level0_c1<= level1_c1(56 downto 0) when count0_c1='0' else level1_c1(55 downto 0) & (0 downto 0 => '0');

   R <= level0_c1;
   sCount_c1 <= count5_c1 & count4_c1 & count3_c1 & count2_c1 & count1_c1 & count0_c1;
   Count <= sCount_c1;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_66_Freq100_uid11
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_66_Freq100_uid11 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(65 downto 0);
          Y : in  std_logic_vector(65 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of IntAdder_66_Freq100_uid11 is
signal Cin_1_c1, Cin_1_c2 :  std_logic;
signal X_1_c1, X_1_c2 :  std_logic_vector(66 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2 :  std_logic_vector(66 downto 0);
signal S_1_c2 :  std_logic_vector(66 downto 0);
signal R_1_c2 :  std_logic_vector(65 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_1_c1 <= Y_1_c0;
            end if;
            if ce_2 = '1' then
               Cin_1_c2 <= Cin_1_c1;
               X_1_c2 <= X_1_c1;
               Y_1_c2 <= Y_1_c1;
            end if;
         end if;
      end process;
   Cin_1_c1 <= Cin;
   X_1_c1 <= '0' & X(65 downto 0);
   Y_1_c0 <= '0' & Y(65 downto 0);
   S_1_c2 <= X_1_c2 + Y_1_c2 + Cin_1_c2;
   R_1_c2 <= S_1_c2(65 downto 0);
   R <= R_1_c2 ;
end architecture;

--------------------------------------------------------------------------------
--                             FloatingPointAdder
--                         (FPAdd_11_52_Freq100_uid2)
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2010-2017)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointAdder_64_9_068000 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointAdder_64_9_068000 is
   component RightShifterSticky53_by_max_55_Freq100_uid4 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             S : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(54 downto 0);
             Sticky : out  std_logic   );
   end component;

   component IntAdder_56_Freq100_uid6 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(55 downto 0)   );
   end component;

   component Normalizer_Z_57_57_57_Freq100_uid8 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(56 downto 0);
             Count : out  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(56 downto 0)   );
   end component;

   component IntAdder_66_Freq100_uid11 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(65 downto 0);
             Y : in  std_logic_vector(65 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(65 downto 0)   );
   end component;

signal excExpFracX_c0 :  std_logic_vector(64 downto 0);
signal excExpFracY_c0 :  std_logic_vector(64 downto 0);
signal swap_c0 :  std_logic;
signal eXmeY_c0 :  std_logic_vector(10 downto 0);
signal eYmeX_c0 :  std_logic_vector(10 downto 0);
signal expDiff_c0 :  std_logic_vector(10 downto 0);
signal newX_c0 :  std_logic_vector(65 downto 0);
signal newY_c0 :  std_logic_vector(65 downto 0);
signal expX_c0 :  std_logic_vector(10 downto 0);
signal excX_c0 :  std_logic_vector(1 downto 0);
signal excY_c0 :  std_logic_vector(1 downto 0);
signal signX_c0 :  std_logic;
signal signY_c0 :  std_logic;
signal EffSub_c0, EffSub_c1, EffSub_c2 :  std_logic;
signal sXsYExnXY_c0 :  std_logic_vector(5 downto 0);
signal sdExnXY_c0 :  std_logic_vector(3 downto 0);
signal fracY_c0 :  std_logic_vector(52 downto 0);
signal excRt_c0, excRt_c1, excRt_c2 :  std_logic_vector(1 downto 0);
signal signR_c0, signR_c1 :  std_logic;
signal shiftedOut_c0 :  std_logic;
signal shiftVal_c0 :  std_logic_vector(5 downto 0);
signal shiftedFracY_c0 :  std_logic_vector(54 downto 0);
signal sticky_c0, sticky_c1 :  std_logic;
signal fracYpad_c0 :  std_logic_vector(55 downto 0);
signal EffSubVector_c0 :  std_logic_vector(55 downto 0);
signal fracYpadXorOp_c0 :  std_logic_vector(55 downto 0);
signal fracXpad_c0 :  std_logic_vector(55 downto 0);
signal cInSigAdd_c1 :  std_logic;
signal fracAddResult_c1 :  std_logic_vector(55 downto 0);
signal fracSticky_c1 :  std_logic_vector(56 downto 0);
signal nZerosNew_c1 :  std_logic_vector(5 downto 0);
signal shiftedFrac_c1 :  std_logic_vector(56 downto 0);
signal extendedExpInc_c0, extendedExpInc_c1 :  std_logic_vector(11 downto 0);
signal updatedExp_c1 :  std_logic_vector(12 downto 0);
signal eqdiffsign_c1, eqdiffsign_c2 :  std_logic;
signal expFrac_c1 :  std_logic_vector(65 downto 0);
signal stk_c1 :  std_logic;
signal rnd_c1 :  std_logic;
signal lsb_c1 :  std_logic;
signal needToRound_c1 :  std_logic;
signal RoundedExpFrac_c2 :  std_logic_vector(65 downto 0);
signal upExc_c2 :  std_logic_vector(1 downto 0);
signal fracR_c2 :  std_logic_vector(51 downto 0);
signal expR_c2 :  std_logic_vector(10 downto 0);
signal exExpExc_c2 :  std_logic_vector(3 downto 0);
signal excRt2_c2 :  std_logic_vector(1 downto 0);
signal excR_c2 :  std_logic_vector(1 downto 0);
signal signR2_c1, signR2_c2 :  std_logic;
signal computedR_c2 :  std_logic_vector(65 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               EffSub_c1 <= EffSub_c0;
               excRt_c1 <= excRt_c0;
               signR_c1 <= signR_c0;
               sticky_c1 <= sticky_c0;
               extendedExpInc_c1 <= extendedExpInc_c0;
            end if;
            if ce_2 = '1' then
               EffSub_c2 <= EffSub_c1;
               excRt_c2 <= excRt_c1;
               eqdiffsign_c2 <= eqdiffsign_c1;
               signR2_c2 <= signR2_c1;
            end if;
         end if;
      end process;
   excExpFracX_c0 <= X(65 downto 64) & X(62 downto 0);
   excExpFracY_c0 <= Y(65 downto 64) & Y(62 downto 0);
   swap_c0 <= '1' when excExpFracX_c0 < excExpFracY_c0 else '0';
   -- exponent difference
   eXmeY_c0 <= (X(62 downto 52)) - (Y(62 downto 52));
   eYmeX_c0 <= (Y(62 downto 52)) - (X(62 downto 52));
   expDiff_c0 <= eXmeY_c0 when swap_c0 = '0' else eYmeX_c0;
   -- input swap so that |X|>|Y|
   newX_c0 <= X when swap_c0 = '0' else Y;
   newY_c0 <= Y when swap_c0 = '0' else X;
   -- now we decompose the inputs into their sign, exponent, fraction
   expX_c0<= newX_c0(62 downto 52);
   excX_c0<= newX_c0(65 downto 64);
   excY_c0<= newY_c0(65 downto 64);
   signX_c0<= newX_c0(63);
   signY_c0<= newY_c0(63);
   EffSub_c0 <= signX_c0 xor signY_c0;
   sXsYExnXY_c0 <= signX_c0 & signY_c0 & excX_c0 & excY_c0;
   sdExnXY_c0 <= excX_c0 & excY_c0;
   fracY_c0 <= "00000000000000000000000000000000000000000000000000000" when excY_c0="00" else ('1' & newY_c0(51 downto 0));
   -- Exception management logic
   with sXsYExnXY_c0  select  
   excRt_c0 <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR_c0<= '0' when (sXsYExnXY_c0="100000" or sXsYExnXY_c0="010000") else signX_c0;
   shiftedOut_c0 <= '1' when (expDiff_c0 > 54) else '0';
   shiftVal_c0 <= expDiff_c0(5 downto 0) when shiftedOut_c0='0' else CONV_STD_LOGIC_VECTOR(55,6);
   RightShifterComponent: RightShifterSticky53_by_max_55_Freq100_uid4
      port map ( clk  => clk,
                 S => shiftVal_c0,
                 X => fracY_c0,
                 R => shiftedFracY_c0,
                 Sticky => sticky_c0);
   fracYpad_c0 <= "0" & shiftedFracY_c0;
   EffSubVector_c0 <= (55 downto 0 => EffSub_c0);
   fracYpadXorOp_c0 <= fracYpad_c0 xor EffSubVector_c0;
   fracXpad_c0 <= "01" & (newX_c0(51 downto 0)) & "00";
   cInSigAdd_c1 <= EffSub_c1 and not sticky_c1; -- if we subtract and the sticky was one, some of the negated sticky bits would have absorbed this carry 
   fracAdder: IntAdder_56_Freq100_uid6
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 Cin => cInSigAdd_c1,
                 X => fracXpad_c0,
                 Y => fracYpadXorOp_c0,
                 R => fracAddResult_c1);
   fracSticky_c1<= fracAddResult_c1 & sticky_c1; 
   LZCAndShifter: Normalizer_Z_57_57_57_Freq100_uid8
      port map ( clk  => clk,
                 X => fracSticky_c1,
                 Count => nZerosNew_c1,
                 R => shiftedFrac_c1);
   extendedExpInc_c0<= ("0" & expX_c0) + '1';
   updatedExp_c1 <= ("0" &extendedExpInc_c1) - ("0000000" & nZerosNew_c1);
   eqdiffsign_c1 <= '1' when nZerosNew_c1="111111" else '0';
   expFrac_c1<= updatedExp_c1 & shiftedFrac_c1(55 downto 3);
   stk_c1<= shiftedFrac_c1(2) or shiftedFrac_c1(1) or shiftedFrac_c1(0);
   rnd_c1<= shiftedFrac_c1(3);
   lsb_c1<= shiftedFrac_c1(4);
   needToRound_c1<= '1' when (rnd_c1='1' and stk_c1='1') or (rnd_c1='1' and stk_c1='0' and lsb_c1='1')
  else '0';
   roundingAdder: IntAdder_66_Freq100_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 Cin => needToRound_c1,
                 X => expFrac_c1,
                 Y => "000000000000000000000000000000000000000000000000000000000000000000",
                 R => RoundedExpFrac_c2);
   -- possible update to exception bits
   upExc_c2 <= RoundedExpFrac_c2(65 downto 64);
   fracR_c2 <= RoundedExpFrac_c2(52 downto 1);
   expR_c2 <= RoundedExpFrac_c2(63 downto 53);
   exExpExc_c2 <= upExc_c2 & excRt_c2;
   with exExpExc_c2  select  
   excRt2_c2<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR_c2 <= "00" when (eqdiffsign_c2='1' and EffSub_c2='1'  and not(excRt_c2="11")) else excRt2_c2;
   signR2_c1 <= '0' when (eqdiffsign_c1='1' and EffSub_c1='1') else signR_c1;
   computedR_c2 <= excR_c2 & signR2_c2 & expR_c2 & fracR_c2;
   R <= computedR_c2;
end architecture;




--------------------------------------------------------------------------------
--                RightShifterSticky24_by_max_26_Freq800_uid4
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X S
-- Output signals: R Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifterSticky24_by_max_26_Freq800_uid4 is
    port (clk, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(25 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of RightShifterSticky24_by_max_26_Freq800_uid4 is
signal ps_c2, ps_c3, ps_c4, ps_c5, ps_c6, ps_c7, ps_c8 :  std_logic_vector(4 downto 0);
signal Xpadded_c2 :  std_logic_vector(25 downto 0);
signal level5_c2, level5_c3 :  std_logic_vector(25 downto 0);
signal stk4_c3, stk4_c4 :  std_logic;
signal level4_c2, level4_c3, level4_c4 :  std_logic_vector(25 downto 0);
signal stk3_c4, stk3_c5 :  std_logic;
signal level3_c3, level3_c4, level3_c5 :  std_logic_vector(25 downto 0);
signal stk2_c5, stk2_c6, stk2_c7 :  std_logic;
signal level2_c3, level2_c4, level2_c5, level2_c6, level2_c7 :  std_logic_vector(25 downto 0);
signal stk1_c7, stk1_c8 :  std_logic;
signal level1_c3, level1_c4, level1_c5, level1_c6, level1_c7, level1_c8 :  std_logic_vector(25 downto 0);
signal stk0_c8 :  std_logic;
signal level0_c3 :  std_logic_vector(25 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_3 = '1' then
               ps_c3 <= ps_c2;
               level5_c3 <= level5_c2;
               level4_c3 <= level4_c2;
            end if;
            if ce_4 = '1' then
               ps_c4 <= ps_c3;
               stk4_c4 <= stk4_c3;
               level4_c4 <= level4_c3;
               level3_c4 <= level3_c3;
               level2_c4 <= level2_c3;
               level1_c4 <= level1_c3;
            end if;
            if ce_5 = '1' then
               ps_c5 <= ps_c4;
               stk3_c5 <= stk3_c4;
               level3_c5 <= level3_c4;
               level2_c5 <= level2_c4;
               level1_c5 <= level1_c4;
            end if;
            if ce_6 = '1' then
               ps_c6 <= ps_c5;
               stk2_c6 <= stk2_c5;
               level2_c6 <= level2_c5;
               level1_c6 <= level1_c5;
            end if;
            if ce_7 = '1' then
               ps_c7 <= ps_c6;
               stk2_c7 <= stk2_c6;
               level2_c7 <= level2_c6;
               level1_c7 <= level1_c6;
            end if;
            if ce_8 = '1' then
               ps_c8 <= ps_c7;
               stk1_c8 <= stk1_c7;
               level1_c8 <= level1_c7;
            end if;
         end if;
      end process;
   ps_c2<= S;
   Xpadded_c2 <= X&(1 downto 0 => '0');
   level5_c2<= Xpadded_c2;
   stk4_c3 <= '1' when (level5_c3(15 downto 0)/="0000000000000000" and ps_c3(4)='1')   else '0';
   level4_c2 <=  level5_c2 when  ps_c2(4)='0'    else (15 downto 0 => '0') & level5_c2(25 downto 16);
   stk3_c4 <= '1' when (level4_c4(7 downto 0)/="00000000" and ps_c4(3)='1') or stk4_c4 ='1'   else '0';
   level3_c3 <=  level4_c3 when  ps_c3(3)='0'    else (7 downto 0 => '0') & level4_c3(25 downto 8);
   stk2_c5 <= '1' when (level3_c5(3 downto 0)/="0000" and ps_c5(2)='1') or stk3_c5 ='1'   else '0';
   level2_c3 <=  level3_c3 when  ps_c3(2)='0'    else (3 downto 0 => '0') & level3_c3(25 downto 4);
   stk1_c7 <= '1' when (level2_c7(1 downto 0)/="00" and ps_c7(1)='1') or stk2_c7 ='1'   else '0';
   level1_c3 <=  level2_c3 when  ps_c3(1)='0'    else (1 downto 0 => '0') & level2_c3(25 downto 2);
   stk0_c8 <= '1' when (level1_c8(0 downto 0)/="0" and ps_c8(0)='1') or stk1_c8 ='1'   else '0';
   level0_c3 <=  level1_c3 when  ps_c3(0)='0'    else (0 downto 0 => '0') & level1_c3(25 downto 1);
   R <= level0_c3;
   Sticky <= stk0_c8;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_27_Freq800_uid6
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 16 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_Freq800_uid6 is
    port (clk, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17 : in std_logic;
          X : in  std_logic_vector(26 downto 0);
          Y : in  std_logic_vector(26 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_Freq800_uid6 is
signal Cin_1_c8, Cin_1_c9 :  std_logic;
signal X_1_c1, X_1_c2, X_1_c3, X_1_c4, X_1_c5, X_1_c6, X_1_c7, X_1_c8, X_1_c9 :  std_logic_vector(3 downto 0);
signal Y_1_c4, Y_1_c5, Y_1_c6, Y_1_c7, Y_1_c8, Y_1_c9 :  std_logic_vector(3 downto 0);
signal S_1_c9 :  std_logic_vector(3 downto 0);
signal R_1_c9, R_1_c10, R_1_c11, R_1_c12, R_1_c13, R_1_c14, R_1_c15, R_1_c16, R_1_c17 :  std_logic_vector(2 downto 0);
signal Cin_2_c9, Cin_2_c10 :  std_logic;
signal X_2_c1, X_2_c2, X_2_c3, X_2_c4, X_2_c5, X_2_c6, X_2_c7, X_2_c8, X_2_c9, X_2_c10 :  std_logic_vector(3 downto 0);
signal Y_2_c4, Y_2_c5, Y_2_c6, Y_2_c7, Y_2_c8, Y_2_c9, Y_2_c10 :  std_logic_vector(3 downto 0);
signal S_2_c10 :  std_logic_vector(3 downto 0);
signal R_2_c10, R_2_c11, R_2_c12, R_2_c13, R_2_c14, R_2_c15, R_2_c16, R_2_c17 :  std_logic_vector(2 downto 0);
signal Cin_3_c10, Cin_3_c11 :  std_logic;
signal X_3_c1, X_3_c2, X_3_c3, X_3_c4, X_3_c5, X_3_c6, X_3_c7, X_3_c8, X_3_c9, X_3_c10, X_3_c11 :  std_logic_vector(3 downto 0);
signal Y_3_c4, Y_3_c5, Y_3_c6, Y_3_c7, Y_3_c8, Y_3_c9, Y_3_c10, Y_3_c11 :  std_logic_vector(3 downto 0);
signal S_3_c11 :  std_logic_vector(3 downto 0);
signal R_3_c11, R_3_c12, R_3_c13, R_3_c14, R_3_c15, R_3_c16, R_3_c17 :  std_logic_vector(2 downto 0);
signal Cin_4_c11, Cin_4_c12 :  std_logic;
signal X_4_c1, X_4_c2, X_4_c3, X_4_c4, X_4_c5, X_4_c6, X_4_c7, X_4_c8, X_4_c9, X_4_c10, X_4_c11, X_4_c12 :  std_logic_vector(3 downto 0);
signal Y_4_c4, Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8, Y_4_c9, Y_4_c10, Y_4_c11, Y_4_c12 :  std_logic_vector(3 downto 0);
signal S_4_c12 :  std_logic_vector(3 downto 0);
signal R_4_c12, R_4_c13, R_4_c14, R_4_c15, R_4_c16, R_4_c17 :  std_logic_vector(2 downto 0);
signal Cin_5_c12, Cin_5_c13 :  std_logic;
signal X_5_c1, X_5_c2, X_5_c3, X_5_c4, X_5_c5, X_5_c6, X_5_c7, X_5_c8, X_5_c9, X_5_c10, X_5_c11, X_5_c12, X_5_c13 :  std_logic_vector(3 downto 0);
signal Y_5_c4, Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9, Y_5_c10, Y_5_c11, Y_5_c12, Y_5_c13 :  std_logic_vector(3 downto 0);
signal S_5_c13 :  std_logic_vector(3 downto 0);
signal R_5_c13, R_5_c14, R_5_c15, R_5_c16, R_5_c17 :  std_logic_vector(2 downto 0);
signal Cin_6_c13, Cin_6_c14 :  std_logic;
signal X_6_c1, X_6_c2, X_6_c3, X_6_c4, X_6_c5, X_6_c6, X_6_c7, X_6_c8, X_6_c9, X_6_c10, X_6_c11, X_6_c12, X_6_c13, X_6_c14 :  std_logic_vector(3 downto 0);
signal Y_6_c4, Y_6_c5, Y_6_c6, Y_6_c7, Y_6_c8, Y_6_c9, Y_6_c10, Y_6_c11, Y_6_c12, Y_6_c13, Y_6_c14 :  std_logic_vector(3 downto 0);
signal S_6_c14 :  std_logic_vector(3 downto 0);
signal R_6_c14, R_6_c15, R_6_c16, R_6_c17 :  std_logic_vector(2 downto 0);
signal Cin_7_c14, Cin_7_c15 :  std_logic;
signal X_7_c1, X_7_c2, X_7_c3, X_7_c4, X_7_c5, X_7_c6, X_7_c7, X_7_c8, X_7_c9, X_7_c10, X_7_c11, X_7_c12, X_7_c13, X_7_c14, X_7_c15 :  std_logic_vector(3 downto 0);
signal Y_7_c4, Y_7_c5, Y_7_c6, Y_7_c7, Y_7_c8, Y_7_c9, Y_7_c10, Y_7_c11, Y_7_c12, Y_7_c13, Y_7_c14, Y_7_c15 :  std_logic_vector(3 downto 0);
signal S_7_c15 :  std_logic_vector(3 downto 0);
signal R_7_c15, R_7_c16, R_7_c17 :  std_logic_vector(2 downto 0);
signal Cin_8_c15, Cin_8_c16 :  std_logic;
signal X_8_c1, X_8_c2, X_8_c3, X_8_c4, X_8_c5, X_8_c6, X_8_c7, X_8_c8, X_8_c9, X_8_c10, X_8_c11, X_8_c12, X_8_c13, X_8_c14, X_8_c15, X_8_c16 :  std_logic_vector(3 downto 0);
signal Y_8_c4, Y_8_c5, Y_8_c6, Y_8_c7, Y_8_c8, Y_8_c9, Y_8_c10, Y_8_c11, Y_8_c12, Y_8_c13, Y_8_c14, Y_8_c15, Y_8_c16 :  std_logic_vector(3 downto 0);
signal S_8_c16 :  std_logic_vector(3 downto 0);
signal R_8_c16, R_8_c17 :  std_logic_vector(2 downto 0);
signal Cin_9_c16, Cin_9_c17 :  std_logic;
signal X_9_c1, X_9_c2, X_9_c3, X_9_c4, X_9_c5, X_9_c6, X_9_c7, X_9_c8, X_9_c9, X_9_c10, X_9_c11, X_9_c12, X_9_c13, X_9_c14, X_9_c15, X_9_c16, X_9_c17 :  std_logic_vector(3 downto 0);
signal Y_9_c4, Y_9_c5, Y_9_c6, Y_9_c7, Y_9_c8, Y_9_c9, Y_9_c10, Y_9_c11, Y_9_c12, Y_9_c13, Y_9_c14, Y_9_c15, Y_9_c16, Y_9_c17 :  std_logic_vector(3 downto 0);
signal S_9_c17 :  std_logic_vector(3 downto 0);
signal R_9_c17 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_2 = '1' then
               X_1_c2 <= X_1_c1;
               X_2_c2 <= X_2_c1;
               X_3_c2 <= X_3_c1;
               X_4_c2 <= X_4_c1;
               X_5_c2 <= X_5_c1;
               X_6_c2 <= X_6_c1;
               X_7_c2 <= X_7_c1;
               X_8_c2 <= X_8_c1;
               X_9_c2 <= X_9_c1;
            end if;
            if ce_3 = '1' then
               X_1_c3 <= X_1_c2;
               X_2_c3 <= X_2_c2;
               X_3_c3 <= X_3_c2;
               X_4_c3 <= X_4_c2;
               X_5_c3 <= X_5_c2;
               X_6_c3 <= X_6_c2;
               X_7_c3 <= X_7_c2;
               X_8_c3 <= X_8_c2;
               X_9_c3 <= X_9_c2;
            end if;
            if ce_4 = '1' then
               X_1_c4 <= X_1_c3;
               X_2_c4 <= X_2_c3;
               X_3_c4 <= X_3_c3;
               X_4_c4 <= X_4_c3;
               X_5_c4 <= X_5_c3;
               X_6_c4 <= X_6_c3;
               X_7_c4 <= X_7_c3;
               X_8_c4 <= X_8_c3;
               X_9_c4 <= X_9_c3;
            end if;
            if ce_5 = '1' then
               X_1_c5 <= X_1_c4;
               Y_1_c5 <= Y_1_c4;
               X_2_c5 <= X_2_c4;
               Y_2_c5 <= Y_2_c4;
               X_3_c5 <= X_3_c4;
               Y_3_c5 <= Y_3_c4;
               X_4_c5 <= X_4_c4;
               Y_4_c5 <= Y_4_c4;
               X_5_c5 <= X_5_c4;
               Y_5_c5 <= Y_5_c4;
               X_6_c5 <= X_6_c4;
               Y_6_c5 <= Y_6_c4;
               X_7_c5 <= X_7_c4;
               Y_7_c5 <= Y_7_c4;
               X_8_c5 <= X_8_c4;
               Y_8_c5 <= Y_8_c4;
               X_9_c5 <= X_9_c4;
               Y_9_c5 <= Y_9_c4;
            end if;
            if ce_6 = '1' then
               X_1_c6 <= X_1_c5;
               Y_1_c6 <= Y_1_c5;
               X_2_c6 <= X_2_c5;
               Y_2_c6 <= Y_2_c5;
               X_3_c6 <= X_3_c5;
               Y_3_c6 <= Y_3_c5;
               X_4_c6 <= X_4_c5;
               Y_4_c6 <= Y_4_c5;
               X_5_c6 <= X_5_c5;
               Y_5_c6 <= Y_5_c5;
               X_6_c6 <= X_6_c5;
               Y_6_c6 <= Y_6_c5;
               X_7_c6 <= X_7_c5;
               Y_7_c6 <= Y_7_c5;
               X_8_c6 <= X_8_c5;
               Y_8_c6 <= Y_8_c5;
               X_9_c6 <= X_9_c5;
               Y_9_c6 <= Y_9_c5;
            end if;
            if ce_7 = '1' then
               X_1_c7 <= X_1_c6;
               Y_1_c7 <= Y_1_c6;
               X_2_c7 <= X_2_c6;
               Y_2_c7 <= Y_2_c6;
               X_3_c7 <= X_3_c6;
               Y_3_c7 <= Y_3_c6;
               X_4_c7 <= X_4_c6;
               Y_4_c7 <= Y_4_c6;
               X_5_c7 <= X_5_c6;
               Y_5_c7 <= Y_5_c6;
               X_6_c7 <= X_6_c6;
               Y_6_c7 <= Y_6_c6;
               X_7_c7 <= X_7_c6;
               Y_7_c7 <= Y_7_c6;
               X_8_c7 <= X_8_c6;
               Y_8_c7 <= Y_8_c6;
               X_9_c7 <= X_9_c6;
               Y_9_c7 <= Y_9_c6;
            end if;
            if ce_8 = '1' then
               X_1_c8 <= X_1_c7;
               Y_1_c8 <= Y_1_c7;
               X_2_c8 <= X_2_c7;
               Y_2_c8 <= Y_2_c7;
               X_3_c8 <= X_3_c7;
               Y_3_c8 <= Y_3_c7;
               X_4_c8 <= X_4_c7;
               Y_4_c8 <= Y_4_c7;
               X_5_c8 <= X_5_c7;
               Y_5_c8 <= Y_5_c7;
               X_6_c8 <= X_6_c7;
               Y_6_c8 <= Y_6_c7;
               X_7_c8 <= X_7_c7;
               Y_7_c8 <= Y_7_c7;
               X_8_c8 <= X_8_c7;
               Y_8_c8 <= Y_8_c7;
               X_9_c8 <= X_9_c7;
               Y_9_c8 <= Y_9_c7;
            end if;
            if ce_9 = '1' then
               Cin_1_c9 <= Cin_1_c8;
               X_1_c9 <= X_1_c8;
               Y_1_c9 <= Y_1_c8;
               X_2_c9 <= X_2_c8;
               Y_2_c9 <= Y_2_c8;
               X_3_c9 <= X_3_c8;
               Y_3_c9 <= Y_3_c8;
               X_4_c9 <= X_4_c8;
               Y_4_c9 <= Y_4_c8;
               X_5_c9 <= X_5_c8;
               Y_5_c9 <= Y_5_c8;
               X_6_c9 <= X_6_c8;
               Y_6_c9 <= Y_6_c8;
               X_7_c9 <= X_7_c8;
               Y_7_c9 <= Y_7_c8;
               X_8_c9 <= X_8_c8;
               Y_8_c9 <= Y_8_c8;
               X_9_c9 <= X_9_c8;
               Y_9_c9 <= Y_9_c8;
            end if;
            if ce_10 = '1' then
               R_1_c10 <= R_1_c9;
               Cin_2_c10 <= Cin_2_c9;
               X_2_c10 <= X_2_c9;
               Y_2_c10 <= Y_2_c9;
               X_3_c10 <= X_3_c9;
               Y_3_c10 <= Y_3_c9;
               X_4_c10 <= X_4_c9;
               Y_4_c10 <= Y_4_c9;
               X_5_c10 <= X_5_c9;
               Y_5_c10 <= Y_5_c9;
               X_6_c10 <= X_6_c9;
               Y_6_c10 <= Y_6_c9;
               X_7_c10 <= X_7_c9;
               Y_7_c10 <= Y_7_c9;
               X_8_c10 <= X_8_c9;
               Y_8_c10 <= Y_8_c9;
               X_9_c10 <= X_9_c9;
               Y_9_c10 <= Y_9_c9;
            end if;
            if ce_11 = '1' then
               R_1_c11 <= R_1_c10;
               R_2_c11 <= R_2_c10;
               Cin_3_c11 <= Cin_3_c10;
               X_3_c11 <= X_3_c10;
               Y_3_c11 <= Y_3_c10;
               X_4_c11 <= X_4_c10;
               Y_4_c11 <= Y_4_c10;
               X_5_c11 <= X_5_c10;
               Y_5_c11 <= Y_5_c10;
               X_6_c11 <= X_6_c10;
               Y_6_c11 <= Y_6_c10;
               X_7_c11 <= X_7_c10;
               Y_7_c11 <= Y_7_c10;
               X_8_c11 <= X_8_c10;
               Y_8_c11 <= Y_8_c10;
               X_9_c11 <= X_9_c10;
               Y_9_c11 <= Y_9_c10;
            end if;
            if ce_12 = '1' then
               R_1_c12 <= R_1_c11;
               R_2_c12 <= R_2_c11;
               R_3_c12 <= R_3_c11;
               Cin_4_c12 <= Cin_4_c11;
               X_4_c12 <= X_4_c11;
               Y_4_c12 <= Y_4_c11;
               X_5_c12 <= X_5_c11;
               Y_5_c12 <= Y_5_c11;
               X_6_c12 <= X_6_c11;
               Y_6_c12 <= Y_6_c11;
               X_7_c12 <= X_7_c11;
               Y_7_c12 <= Y_7_c11;
               X_8_c12 <= X_8_c11;
               Y_8_c12 <= Y_8_c11;
               X_9_c12 <= X_9_c11;
               Y_9_c12 <= Y_9_c11;
            end if;
            if ce_13 = '1' then
               R_1_c13 <= R_1_c12;
               R_2_c13 <= R_2_c12;
               R_3_c13 <= R_3_c12;
               R_4_c13 <= R_4_c12;
               Cin_5_c13 <= Cin_5_c12;
               X_5_c13 <= X_5_c12;
               Y_5_c13 <= Y_5_c12;
               X_6_c13 <= X_6_c12;
               Y_6_c13 <= Y_6_c12;
               X_7_c13 <= X_7_c12;
               Y_7_c13 <= Y_7_c12;
               X_8_c13 <= X_8_c12;
               Y_8_c13 <= Y_8_c12;
               X_9_c13 <= X_9_c12;
               Y_9_c13 <= Y_9_c12;
            end if;
            if ce_14 = '1' then
               R_1_c14 <= R_1_c13;
               R_2_c14 <= R_2_c13;
               R_3_c14 <= R_3_c13;
               R_4_c14 <= R_4_c13;
               R_5_c14 <= R_5_c13;
               Cin_6_c14 <= Cin_6_c13;
               X_6_c14 <= X_6_c13;
               Y_6_c14 <= Y_6_c13;
               X_7_c14 <= X_7_c13;
               Y_7_c14 <= Y_7_c13;
               X_8_c14 <= X_8_c13;
               Y_8_c14 <= Y_8_c13;
               X_9_c14 <= X_9_c13;
               Y_9_c14 <= Y_9_c13;
            end if;
            if ce_15 = '1' then
               R_1_c15 <= R_1_c14;
               R_2_c15 <= R_2_c14;
               R_3_c15 <= R_3_c14;
               R_4_c15 <= R_4_c14;
               R_5_c15 <= R_5_c14;
               R_6_c15 <= R_6_c14;
               Cin_7_c15 <= Cin_7_c14;
               X_7_c15 <= X_7_c14;
               Y_7_c15 <= Y_7_c14;
               X_8_c15 <= X_8_c14;
               Y_8_c15 <= Y_8_c14;
               X_9_c15 <= X_9_c14;
               Y_9_c15 <= Y_9_c14;
            end if;
            if ce_16 = '1' then
               R_1_c16 <= R_1_c15;
               R_2_c16 <= R_2_c15;
               R_3_c16 <= R_3_c15;
               R_4_c16 <= R_4_c15;
               R_5_c16 <= R_5_c15;
               R_6_c16 <= R_6_c15;
               R_7_c16 <= R_7_c15;
               Cin_8_c16 <= Cin_8_c15;
               X_8_c16 <= X_8_c15;
               Y_8_c16 <= Y_8_c15;
               X_9_c16 <= X_9_c15;
               Y_9_c16 <= Y_9_c15;
            end if;
            if ce_17 = '1' then
               R_1_c17 <= R_1_c16;
               R_2_c17 <= R_2_c16;
               R_3_c17 <= R_3_c16;
               R_4_c17 <= R_4_c16;
               R_5_c17 <= R_5_c16;
               R_6_c17 <= R_6_c16;
               R_7_c17 <= R_7_c16;
               R_8_c17 <= R_8_c16;
               Cin_9_c17 <= Cin_9_c16;
               X_9_c17 <= X_9_c16;
               Y_9_c17 <= Y_9_c16;
            end if;
         end if;
      end process;
   Cin_1_c8 <= Cin;
   X_1_c1 <= '0' & X(2 downto 0);
   Y_1_c4 <= '0' & Y(2 downto 0);
   S_1_c9 <= X_1_c9 + Y_1_c9 + Cin_1_c9;
   R_1_c9 <= S_1_c9(2 downto 0);
   Cin_2_c9 <= S_1_c9(3);
   X_2_c1 <= '0' & X(5 downto 3);
   Y_2_c4 <= '0' & Y(5 downto 3);
   S_2_c10 <= X_2_c10 + Y_2_c10 + Cin_2_c10;
   R_2_c10 <= S_2_c10(2 downto 0);
   Cin_3_c10 <= S_2_c10(3);
   X_3_c1 <= '0' & X(8 downto 6);
   Y_3_c4 <= '0' & Y(8 downto 6);
   S_3_c11 <= X_3_c11 + Y_3_c11 + Cin_3_c11;
   R_3_c11 <= S_3_c11(2 downto 0);
   Cin_4_c11 <= S_3_c11(3);
   X_4_c1 <= '0' & X(11 downto 9);
   Y_4_c4 <= '0' & Y(11 downto 9);
   S_4_c12 <= X_4_c12 + Y_4_c12 + Cin_4_c12;
   R_4_c12 <= S_4_c12(2 downto 0);
   Cin_5_c12 <= S_4_c12(3);
   X_5_c1 <= '0' & X(14 downto 12);
   Y_5_c4 <= '0' & Y(14 downto 12);
   S_5_c13 <= X_5_c13 + Y_5_c13 + Cin_5_c13;
   R_5_c13 <= S_5_c13(2 downto 0);
   Cin_6_c13 <= S_5_c13(3);
   X_6_c1 <= '0' & X(17 downto 15);
   Y_6_c4 <= '0' & Y(17 downto 15);
   S_6_c14 <= X_6_c14 + Y_6_c14 + Cin_6_c14;
   R_6_c14 <= S_6_c14(2 downto 0);
   Cin_7_c14 <= S_6_c14(3);
   X_7_c1 <= '0' & X(20 downto 18);
   Y_7_c4 <= '0' & Y(20 downto 18);
   S_7_c15 <= X_7_c15 + Y_7_c15 + Cin_7_c15;
   R_7_c15 <= S_7_c15(2 downto 0);
   Cin_8_c15 <= S_7_c15(3);
   X_8_c1 <= '0' & X(23 downto 21);
   Y_8_c4 <= '0' & Y(23 downto 21);
   S_8_c16 <= X_8_c16 + Y_8_c16 + Cin_8_c16;
   R_8_c16 <= S_8_c16(2 downto 0);
   Cin_9_c16 <= S_8_c16(3);
   X_9_c1 <= '0' & X(26 downto 24);
   Y_9_c4 <= '0' & Y(26 downto 24);
   S_9_c17 <= X_9_c17 + Y_9_c17 + Cin_9_c17;
   R_9_c17 <= S_9_c17(2 downto 0);
   R <= R_9_c17 & R_8_c17 & R_7_c17 & R_6_c17 & R_5_c17 & R_4_c17 & R_3_c17 & R_2_c17 & R_1_c17 ;
end architecture;

--------------------------------------------------------------------------------
--                     Normalizer_Z_28_28_28_Freq800_uid8
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_28_28_28_Freq800_uid8 is
    port (clk, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23 : in std_logic;
          X : in  std_logic_vector(27 downto 0);
          Count : out  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of Normalizer_Z_28_28_28_Freq800_uid8 is
signal level5_c17, level5_c18 :  std_logic_vector(27 downto 0);
signal count4_c18, count4_c19, count4_c20, count4_c21, count4_c22 :  std_logic;
signal level4_c18, level4_c19 :  std_logic_vector(27 downto 0);
signal count3_c19, count3_c20, count3_c21, count3_c22 :  std_logic;
signal level3_c19, level3_c20 :  std_logic_vector(27 downto 0);
signal count2_c20, count2_c21, count2_c22 :  std_logic;
signal level2_c20, level2_c21, level2_c22 :  std_logic_vector(27 downto 0);
signal count1_c21, count1_c22 :  std_logic;
signal level1_c22, level1_c23 :  std_logic_vector(27 downto 0);
signal count0_c22, count0_c23 :  std_logic;
signal level0_c23 :  std_logic_vector(27 downto 0);
signal sCount_c22 :  std_logic_vector(4 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_18 = '1' then
               level5_c18 <= level5_c17;
            end if;
            if ce_19 = '1' then
               count4_c19 <= count4_c18;
               level4_c19 <= level4_c18;
            end if;
            if ce_20 = '1' then
               count4_c20 <= count4_c19;
               count3_c20 <= count3_c19;
               level3_c20 <= level3_c19;
            end if;
            if ce_21 = '1' then
               count4_c21 <= count4_c20;
               count3_c21 <= count3_c20;
               count2_c21 <= count2_c20;
               level2_c21 <= level2_c20;
            end if;
            if ce_22 = '1' then
               count4_c22 <= count4_c21;
               count3_c22 <= count3_c21;
               count2_c22 <= count2_c21;
               level2_c22 <= level2_c21;
               count1_c22 <= count1_c21;
            end if;
            if ce_23 = '1' then
               level1_c23 <= level1_c22;
               count0_c23 <= count0_c22;
            end if;
         end if;
      end process;
   level5_c17 <= X ;
   count4_c18<= '1' when level5_c18(27 downto 12) = (27 downto 12=>'0') else '0';
   level4_c18<= level5_c18(27 downto 0) when count4_c18='0' else level5_c18(11 downto 0) & (15 downto 0 => '0');

   count3_c19<= '1' when level4_c19(27 downto 20) = (27 downto 20=>'0') else '0';
   level3_c19<= level4_c19(27 downto 0) when count3_c19='0' else level4_c19(19 downto 0) & (7 downto 0 => '0');

   count2_c20<= '1' when level3_c20(27 downto 24) = (27 downto 24=>'0') else '0';
   level2_c20<= level3_c20(27 downto 0) when count2_c20='0' else level3_c20(23 downto 0) & (3 downto 0 => '0');

   count1_c21<= '1' when level2_c21(27 downto 26) = (27 downto 26=>'0') else '0';
   level1_c22<= level2_c22(27 downto 0) when count1_c22='0' else level2_c22(25 downto 0) & (1 downto 0 => '0');

   count0_c22<= '1' when level1_c22(27 downto 27) = (27 downto 27=>'0') else '0';
   level0_c23<= level1_c23(27 downto 0) when count0_c23='0' else level1_c23(26 downto 0) & (0 downto 0 => '0');

   R <= level0_c23;
   sCount_c22 <= count4_c22 & count3_c22 & count2_c22 & count1_c22 & count0_c22;
   Count <= sCount_c22;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_Freq800_uid11
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 35 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_Freq800_uid11 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35 : in std_logic;
          X : in  std_logic_vector(33 downto 0);
          Y : in  std_logic_vector(33 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_Freq800_uid11 is
signal Cin_1_c23, Cin_1_c24 :  std_logic;
signal X_1_c23, X_1_c24 :  std_logic_vector(3 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3, Y_1_c4, Y_1_c5, Y_1_c6, Y_1_c7, Y_1_c8, Y_1_c9, Y_1_c10, Y_1_c11, Y_1_c12, Y_1_c13, Y_1_c14, Y_1_c15, Y_1_c16, Y_1_c17, Y_1_c18, Y_1_c19, Y_1_c20, Y_1_c21, Y_1_c22, Y_1_c23, Y_1_c24 :  std_logic_vector(3 downto 0);
signal S_1_c24 :  std_logic_vector(3 downto 0);
signal R_1_c24, R_1_c25, R_1_c26, R_1_c27, R_1_c28, R_1_c29, R_1_c30, R_1_c31, R_1_c32, R_1_c33, R_1_c34, R_1_c35 :  std_logic_vector(2 downto 0);
signal Cin_2_c24, Cin_2_c25 :  std_logic;
signal X_2_c23, X_2_c24, X_2_c25 :  std_logic_vector(3 downto 0);
signal Y_2_c0, Y_2_c1, Y_2_c2, Y_2_c3, Y_2_c4, Y_2_c5, Y_2_c6, Y_2_c7, Y_2_c8, Y_2_c9, Y_2_c10, Y_2_c11, Y_2_c12, Y_2_c13, Y_2_c14, Y_2_c15, Y_2_c16, Y_2_c17, Y_2_c18, Y_2_c19, Y_2_c20, Y_2_c21, Y_2_c22, Y_2_c23, Y_2_c24, Y_2_c25 :  std_logic_vector(3 downto 0);
signal S_2_c25 :  std_logic_vector(3 downto 0);
signal R_2_c25, R_2_c26, R_2_c27, R_2_c28, R_2_c29, R_2_c30, R_2_c31, R_2_c32, R_2_c33, R_2_c34, R_2_c35 :  std_logic_vector(2 downto 0);
signal Cin_3_c25, Cin_3_c26 :  std_logic;
signal X_3_c23, X_3_c24, X_3_c25, X_3_c26 :  std_logic_vector(3 downto 0);
signal Y_3_c0, Y_3_c1, Y_3_c2, Y_3_c3, Y_3_c4, Y_3_c5, Y_3_c6, Y_3_c7, Y_3_c8, Y_3_c9, Y_3_c10, Y_3_c11, Y_3_c12, Y_3_c13, Y_3_c14, Y_3_c15, Y_3_c16, Y_3_c17, Y_3_c18, Y_3_c19, Y_3_c20, Y_3_c21, Y_3_c22, Y_3_c23, Y_3_c24, Y_3_c25, Y_3_c26 :  std_logic_vector(3 downto 0);
signal S_3_c26 :  std_logic_vector(3 downto 0);
signal R_3_c26, R_3_c27, R_3_c28, R_3_c29, R_3_c30, R_3_c31, R_3_c32, R_3_c33, R_3_c34, R_3_c35 :  std_logic_vector(2 downto 0);
signal Cin_4_c26, Cin_4_c27 :  std_logic;
signal X_4_c23, X_4_c24, X_4_c25, X_4_c26, X_4_c27 :  std_logic_vector(3 downto 0);
signal Y_4_c0, Y_4_c1, Y_4_c2, Y_4_c3, Y_4_c4, Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8, Y_4_c9, Y_4_c10, Y_4_c11, Y_4_c12, Y_4_c13, Y_4_c14, Y_4_c15, Y_4_c16, Y_4_c17, Y_4_c18, Y_4_c19, Y_4_c20, Y_4_c21, Y_4_c22, Y_4_c23, Y_4_c24, Y_4_c25, Y_4_c26, Y_4_c27 :  std_logic_vector(3 downto 0);
signal S_4_c27 :  std_logic_vector(3 downto 0);
signal R_4_c27, R_4_c28, R_4_c29, R_4_c30, R_4_c31, R_4_c32, R_4_c33, R_4_c34, R_4_c35 :  std_logic_vector(2 downto 0);
signal Cin_5_c27, Cin_5_c28 :  std_logic;
signal X_5_c23, X_5_c24, X_5_c25, X_5_c26, X_5_c27, X_5_c28 :  std_logic_vector(3 downto 0);
signal Y_5_c0, Y_5_c1, Y_5_c2, Y_5_c3, Y_5_c4, Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9, Y_5_c10, Y_5_c11, Y_5_c12, Y_5_c13, Y_5_c14, Y_5_c15, Y_5_c16, Y_5_c17, Y_5_c18, Y_5_c19, Y_5_c20, Y_5_c21, Y_5_c22, Y_5_c23, Y_5_c24, Y_5_c25, Y_5_c26, Y_5_c27, Y_5_c28 :  std_logic_vector(3 downto 0);
signal S_5_c28 :  std_logic_vector(3 downto 0);
signal R_5_c28, R_5_c29, R_5_c30, R_5_c31, R_5_c32, R_5_c33, R_5_c34, R_5_c35 :  std_logic_vector(2 downto 0);
signal Cin_6_c28, Cin_6_c29 :  std_logic;
signal X_6_c23, X_6_c24, X_6_c25, X_6_c26, X_6_c27, X_6_c28, X_6_c29 :  std_logic_vector(3 downto 0);
signal Y_6_c0, Y_6_c1, Y_6_c2, Y_6_c3, Y_6_c4, Y_6_c5, Y_6_c6, Y_6_c7, Y_6_c8, Y_6_c9, Y_6_c10, Y_6_c11, Y_6_c12, Y_6_c13, Y_6_c14, Y_6_c15, Y_6_c16, Y_6_c17, Y_6_c18, Y_6_c19, Y_6_c20, Y_6_c21, Y_6_c22, Y_6_c23, Y_6_c24, Y_6_c25, Y_6_c26, Y_6_c27, Y_6_c28, Y_6_c29 :  std_logic_vector(3 downto 0);
signal S_6_c29 :  std_logic_vector(3 downto 0);
signal R_6_c29, R_6_c30, R_6_c31, R_6_c32, R_6_c33, R_6_c34, R_6_c35 :  std_logic_vector(2 downto 0);
signal Cin_7_c29, Cin_7_c30 :  std_logic;
signal X_7_c23, X_7_c24, X_7_c25, X_7_c26, X_7_c27, X_7_c28, X_7_c29, X_7_c30 :  std_logic_vector(3 downto 0);
signal Y_7_c0, Y_7_c1, Y_7_c2, Y_7_c3, Y_7_c4, Y_7_c5, Y_7_c6, Y_7_c7, Y_7_c8, Y_7_c9, Y_7_c10, Y_7_c11, Y_7_c12, Y_7_c13, Y_7_c14, Y_7_c15, Y_7_c16, Y_7_c17, Y_7_c18, Y_7_c19, Y_7_c20, Y_7_c21, Y_7_c22, Y_7_c23, Y_7_c24, Y_7_c25, Y_7_c26, Y_7_c27, Y_7_c28, Y_7_c29, Y_7_c30 :  std_logic_vector(3 downto 0);
signal S_7_c30 :  std_logic_vector(3 downto 0);
signal R_7_c30, R_7_c31, R_7_c32, R_7_c33, R_7_c34, R_7_c35 :  std_logic_vector(2 downto 0);
signal Cin_8_c30, Cin_8_c31 :  std_logic;
signal X_8_c23, X_8_c24, X_8_c25, X_8_c26, X_8_c27, X_8_c28, X_8_c29, X_8_c30, X_8_c31 :  std_logic_vector(3 downto 0);
signal Y_8_c0, Y_8_c1, Y_8_c2, Y_8_c3, Y_8_c4, Y_8_c5, Y_8_c6, Y_8_c7, Y_8_c8, Y_8_c9, Y_8_c10, Y_8_c11, Y_8_c12, Y_8_c13, Y_8_c14, Y_8_c15, Y_8_c16, Y_8_c17, Y_8_c18, Y_8_c19, Y_8_c20, Y_8_c21, Y_8_c22, Y_8_c23, Y_8_c24, Y_8_c25, Y_8_c26, Y_8_c27, Y_8_c28, Y_8_c29, Y_8_c30, Y_8_c31 :  std_logic_vector(3 downto 0);
signal S_8_c31 :  std_logic_vector(3 downto 0);
signal R_8_c31, R_8_c32, R_8_c33, R_8_c34, R_8_c35 :  std_logic_vector(2 downto 0);
signal Cin_9_c31, Cin_9_c32 :  std_logic;
signal X_9_c23, X_9_c24, X_9_c25, X_9_c26, X_9_c27, X_9_c28, X_9_c29, X_9_c30, X_9_c31, X_9_c32 :  std_logic_vector(3 downto 0);
signal Y_9_c0, Y_9_c1, Y_9_c2, Y_9_c3, Y_9_c4, Y_9_c5, Y_9_c6, Y_9_c7, Y_9_c8, Y_9_c9, Y_9_c10, Y_9_c11, Y_9_c12, Y_9_c13, Y_9_c14, Y_9_c15, Y_9_c16, Y_9_c17, Y_9_c18, Y_9_c19, Y_9_c20, Y_9_c21, Y_9_c22, Y_9_c23, Y_9_c24, Y_9_c25, Y_9_c26, Y_9_c27, Y_9_c28, Y_9_c29, Y_9_c30, Y_9_c31, Y_9_c32 :  std_logic_vector(3 downto 0);
signal S_9_c32 :  std_logic_vector(3 downto 0);
signal R_9_c32, R_9_c33, R_9_c34, R_9_c35 :  std_logic_vector(2 downto 0);
signal Cin_10_c32, Cin_10_c33 :  std_logic;
signal X_10_c23, X_10_c24, X_10_c25, X_10_c26, X_10_c27, X_10_c28, X_10_c29, X_10_c30, X_10_c31, X_10_c32, X_10_c33 :  std_logic_vector(3 downto 0);
signal Y_10_c0, Y_10_c1, Y_10_c2, Y_10_c3, Y_10_c4, Y_10_c5, Y_10_c6, Y_10_c7, Y_10_c8, Y_10_c9, Y_10_c10, Y_10_c11, Y_10_c12, Y_10_c13, Y_10_c14, Y_10_c15, Y_10_c16, Y_10_c17, Y_10_c18, Y_10_c19, Y_10_c20, Y_10_c21, Y_10_c22, Y_10_c23, Y_10_c24, Y_10_c25, Y_10_c26, Y_10_c27, Y_10_c28, Y_10_c29, Y_10_c30, Y_10_c31, Y_10_c32, Y_10_c33 :  std_logic_vector(3 downto 0);
signal S_10_c33 :  std_logic_vector(3 downto 0);
signal R_10_c33, R_10_c34, R_10_c35 :  std_logic_vector(2 downto 0);
signal Cin_11_c33, Cin_11_c34 :  std_logic;
signal X_11_c23, X_11_c24, X_11_c25, X_11_c26, X_11_c27, X_11_c28, X_11_c29, X_11_c30, X_11_c31, X_11_c32, X_11_c33, X_11_c34 :  std_logic_vector(3 downto 0);
signal Y_11_c0, Y_11_c1, Y_11_c2, Y_11_c3, Y_11_c4, Y_11_c5, Y_11_c6, Y_11_c7, Y_11_c8, Y_11_c9, Y_11_c10, Y_11_c11, Y_11_c12, Y_11_c13, Y_11_c14, Y_11_c15, Y_11_c16, Y_11_c17, Y_11_c18, Y_11_c19, Y_11_c20, Y_11_c21, Y_11_c22, Y_11_c23, Y_11_c24, Y_11_c25, Y_11_c26, Y_11_c27, Y_11_c28, Y_11_c29, Y_11_c30, Y_11_c31, Y_11_c32, Y_11_c33, Y_11_c34 :  std_logic_vector(3 downto 0);
signal S_11_c34 :  std_logic_vector(3 downto 0);
signal R_11_c34, R_11_c35 :  std_logic_vector(2 downto 0);
signal Cin_12_c34, Cin_12_c35 :  std_logic;
signal X_12_c23, X_12_c24, X_12_c25, X_12_c26, X_12_c27, X_12_c28, X_12_c29, X_12_c30, X_12_c31, X_12_c32, X_12_c33, X_12_c34, X_12_c35 :  std_logic_vector(1 downto 0);
signal Y_12_c0, Y_12_c1, Y_12_c2, Y_12_c3, Y_12_c4, Y_12_c5, Y_12_c6, Y_12_c7, Y_12_c8, Y_12_c9, Y_12_c10, Y_12_c11, Y_12_c12, Y_12_c13, Y_12_c14, Y_12_c15, Y_12_c16, Y_12_c17, Y_12_c18, Y_12_c19, Y_12_c20, Y_12_c21, Y_12_c22, Y_12_c23, Y_12_c24, Y_12_c25, Y_12_c26, Y_12_c27, Y_12_c28, Y_12_c29, Y_12_c30, Y_12_c31, Y_12_c32, Y_12_c33, Y_12_c34, Y_12_c35 :  std_logic_vector(1 downto 0);
signal S_12_c35 :  std_logic_vector(1 downto 0);
signal R_12_c35 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_1_c1 <= Y_1_c0;
               Y_2_c1 <= Y_2_c0;
               Y_3_c1 <= Y_3_c0;
               Y_4_c1 <= Y_4_c0;
               Y_5_c1 <= Y_5_c0;
               Y_6_c1 <= Y_6_c0;
               Y_7_c1 <= Y_7_c0;
               Y_8_c1 <= Y_8_c0;
               Y_9_c1 <= Y_9_c0;
               Y_10_c1 <= Y_10_c0;
               Y_11_c1 <= Y_11_c0;
               Y_12_c1 <= Y_12_c0;
            end if;
            if ce_2 = '1' then
               Y_1_c2 <= Y_1_c1;
               Y_2_c2 <= Y_2_c1;
               Y_3_c2 <= Y_3_c1;
               Y_4_c2 <= Y_4_c1;
               Y_5_c2 <= Y_5_c1;
               Y_6_c2 <= Y_6_c1;
               Y_7_c2 <= Y_7_c1;
               Y_8_c2 <= Y_8_c1;
               Y_9_c2 <= Y_9_c1;
               Y_10_c2 <= Y_10_c1;
               Y_11_c2 <= Y_11_c1;
               Y_12_c2 <= Y_12_c1;
            end if;
            if ce_3 = '1' then
               Y_1_c3 <= Y_1_c2;
               Y_2_c3 <= Y_2_c2;
               Y_3_c3 <= Y_3_c2;
               Y_4_c3 <= Y_4_c2;
               Y_5_c3 <= Y_5_c2;
               Y_6_c3 <= Y_6_c2;
               Y_7_c3 <= Y_7_c2;
               Y_8_c3 <= Y_8_c2;
               Y_9_c3 <= Y_9_c2;
               Y_10_c3 <= Y_10_c2;
               Y_11_c3 <= Y_11_c2;
               Y_12_c3 <= Y_12_c2;
            end if;
            if ce_4 = '1' then
               Y_1_c4 <= Y_1_c3;
               Y_2_c4 <= Y_2_c3;
               Y_3_c4 <= Y_3_c3;
               Y_4_c4 <= Y_4_c3;
               Y_5_c4 <= Y_5_c3;
               Y_6_c4 <= Y_6_c3;
               Y_7_c4 <= Y_7_c3;
               Y_8_c4 <= Y_8_c3;
               Y_9_c4 <= Y_9_c3;
               Y_10_c4 <= Y_10_c3;
               Y_11_c4 <= Y_11_c3;
               Y_12_c4 <= Y_12_c3;
            end if;
            if ce_5 = '1' then
               Y_1_c5 <= Y_1_c4;
               Y_2_c5 <= Y_2_c4;
               Y_3_c5 <= Y_3_c4;
               Y_4_c5 <= Y_4_c4;
               Y_5_c5 <= Y_5_c4;
               Y_6_c5 <= Y_6_c4;
               Y_7_c5 <= Y_7_c4;
               Y_8_c5 <= Y_8_c4;
               Y_9_c5 <= Y_9_c4;
               Y_10_c5 <= Y_10_c4;
               Y_11_c5 <= Y_11_c4;
               Y_12_c5 <= Y_12_c4;
            end if;
            if ce_6 = '1' then
               Y_1_c6 <= Y_1_c5;
               Y_2_c6 <= Y_2_c5;
               Y_3_c6 <= Y_3_c5;
               Y_4_c6 <= Y_4_c5;
               Y_5_c6 <= Y_5_c5;
               Y_6_c6 <= Y_6_c5;
               Y_7_c6 <= Y_7_c5;
               Y_8_c6 <= Y_8_c5;
               Y_9_c6 <= Y_9_c5;
               Y_10_c6 <= Y_10_c5;
               Y_11_c6 <= Y_11_c5;
               Y_12_c6 <= Y_12_c5;
            end if;
            if ce_7 = '1' then
               Y_1_c7 <= Y_1_c6;
               Y_2_c7 <= Y_2_c6;
               Y_3_c7 <= Y_3_c6;
               Y_4_c7 <= Y_4_c6;
               Y_5_c7 <= Y_5_c6;
               Y_6_c7 <= Y_6_c6;
               Y_7_c7 <= Y_7_c6;
               Y_8_c7 <= Y_8_c6;
               Y_9_c7 <= Y_9_c6;
               Y_10_c7 <= Y_10_c6;
               Y_11_c7 <= Y_11_c6;
               Y_12_c7 <= Y_12_c6;
            end if;
            if ce_8 = '1' then
               Y_1_c8 <= Y_1_c7;
               Y_2_c8 <= Y_2_c7;
               Y_3_c8 <= Y_3_c7;
               Y_4_c8 <= Y_4_c7;
               Y_5_c8 <= Y_5_c7;
               Y_6_c8 <= Y_6_c7;
               Y_7_c8 <= Y_7_c7;
               Y_8_c8 <= Y_8_c7;
               Y_9_c8 <= Y_9_c7;
               Y_10_c8 <= Y_10_c7;
               Y_11_c8 <= Y_11_c7;
               Y_12_c8 <= Y_12_c7;
            end if;
            if ce_9 = '1' then
               Y_1_c9 <= Y_1_c8;
               Y_2_c9 <= Y_2_c8;
               Y_3_c9 <= Y_3_c8;
               Y_4_c9 <= Y_4_c8;
               Y_5_c9 <= Y_5_c8;
               Y_6_c9 <= Y_6_c8;
               Y_7_c9 <= Y_7_c8;
               Y_8_c9 <= Y_8_c8;
               Y_9_c9 <= Y_9_c8;
               Y_10_c9 <= Y_10_c8;
               Y_11_c9 <= Y_11_c8;
               Y_12_c9 <= Y_12_c8;
            end if;
            if ce_10 = '1' then
               Y_1_c10 <= Y_1_c9;
               Y_2_c10 <= Y_2_c9;
               Y_3_c10 <= Y_3_c9;
               Y_4_c10 <= Y_4_c9;
               Y_5_c10 <= Y_5_c9;
               Y_6_c10 <= Y_6_c9;
               Y_7_c10 <= Y_7_c9;
               Y_8_c10 <= Y_8_c9;
               Y_9_c10 <= Y_9_c9;
               Y_10_c10 <= Y_10_c9;
               Y_11_c10 <= Y_11_c9;
               Y_12_c10 <= Y_12_c9;
            end if;
            if ce_11 = '1' then
               Y_1_c11 <= Y_1_c10;
               Y_2_c11 <= Y_2_c10;
               Y_3_c11 <= Y_3_c10;
               Y_4_c11 <= Y_4_c10;
               Y_5_c11 <= Y_5_c10;
               Y_6_c11 <= Y_6_c10;
               Y_7_c11 <= Y_7_c10;
               Y_8_c11 <= Y_8_c10;
               Y_9_c11 <= Y_9_c10;
               Y_10_c11 <= Y_10_c10;
               Y_11_c11 <= Y_11_c10;
               Y_12_c11 <= Y_12_c10;
            end if;
            if ce_12 = '1' then
               Y_1_c12 <= Y_1_c11;
               Y_2_c12 <= Y_2_c11;
               Y_3_c12 <= Y_3_c11;
               Y_4_c12 <= Y_4_c11;
               Y_5_c12 <= Y_5_c11;
               Y_6_c12 <= Y_6_c11;
               Y_7_c12 <= Y_7_c11;
               Y_8_c12 <= Y_8_c11;
               Y_9_c12 <= Y_9_c11;
               Y_10_c12 <= Y_10_c11;
               Y_11_c12 <= Y_11_c11;
               Y_12_c12 <= Y_12_c11;
            end if;
            if ce_13 = '1' then
               Y_1_c13 <= Y_1_c12;
               Y_2_c13 <= Y_2_c12;
               Y_3_c13 <= Y_3_c12;
               Y_4_c13 <= Y_4_c12;
               Y_5_c13 <= Y_5_c12;
               Y_6_c13 <= Y_6_c12;
               Y_7_c13 <= Y_7_c12;
               Y_8_c13 <= Y_8_c12;
               Y_9_c13 <= Y_9_c12;
               Y_10_c13 <= Y_10_c12;
               Y_11_c13 <= Y_11_c12;
               Y_12_c13 <= Y_12_c12;
            end if;
            if ce_14 = '1' then
               Y_1_c14 <= Y_1_c13;
               Y_2_c14 <= Y_2_c13;
               Y_3_c14 <= Y_3_c13;
               Y_4_c14 <= Y_4_c13;
               Y_5_c14 <= Y_5_c13;
               Y_6_c14 <= Y_6_c13;
               Y_7_c14 <= Y_7_c13;
               Y_8_c14 <= Y_8_c13;
               Y_9_c14 <= Y_9_c13;
               Y_10_c14 <= Y_10_c13;
               Y_11_c14 <= Y_11_c13;
               Y_12_c14 <= Y_12_c13;
            end if;
            if ce_15 = '1' then
               Y_1_c15 <= Y_1_c14;
               Y_2_c15 <= Y_2_c14;
               Y_3_c15 <= Y_3_c14;
               Y_4_c15 <= Y_4_c14;
               Y_5_c15 <= Y_5_c14;
               Y_6_c15 <= Y_6_c14;
               Y_7_c15 <= Y_7_c14;
               Y_8_c15 <= Y_8_c14;
               Y_9_c15 <= Y_9_c14;
               Y_10_c15 <= Y_10_c14;
               Y_11_c15 <= Y_11_c14;
               Y_12_c15 <= Y_12_c14;
            end if;
            if ce_16 = '1' then
               Y_1_c16 <= Y_1_c15;
               Y_2_c16 <= Y_2_c15;
               Y_3_c16 <= Y_3_c15;
               Y_4_c16 <= Y_4_c15;
               Y_5_c16 <= Y_5_c15;
               Y_6_c16 <= Y_6_c15;
               Y_7_c16 <= Y_7_c15;
               Y_8_c16 <= Y_8_c15;
               Y_9_c16 <= Y_9_c15;
               Y_10_c16 <= Y_10_c15;
               Y_11_c16 <= Y_11_c15;
               Y_12_c16 <= Y_12_c15;
            end if;
            if ce_17 = '1' then
               Y_1_c17 <= Y_1_c16;
               Y_2_c17 <= Y_2_c16;
               Y_3_c17 <= Y_3_c16;
               Y_4_c17 <= Y_4_c16;
               Y_5_c17 <= Y_5_c16;
               Y_6_c17 <= Y_6_c16;
               Y_7_c17 <= Y_7_c16;
               Y_8_c17 <= Y_8_c16;
               Y_9_c17 <= Y_9_c16;
               Y_10_c17 <= Y_10_c16;
               Y_11_c17 <= Y_11_c16;
               Y_12_c17 <= Y_12_c16;
            end if;
            if ce_18 = '1' then
               Y_1_c18 <= Y_1_c17;
               Y_2_c18 <= Y_2_c17;
               Y_3_c18 <= Y_3_c17;
               Y_4_c18 <= Y_4_c17;
               Y_5_c18 <= Y_5_c17;
               Y_6_c18 <= Y_6_c17;
               Y_7_c18 <= Y_7_c17;
               Y_8_c18 <= Y_8_c17;
               Y_9_c18 <= Y_9_c17;
               Y_10_c18 <= Y_10_c17;
               Y_11_c18 <= Y_11_c17;
               Y_12_c18 <= Y_12_c17;
            end if;
            if ce_19 = '1' then
               Y_1_c19 <= Y_1_c18;
               Y_2_c19 <= Y_2_c18;
               Y_3_c19 <= Y_3_c18;
               Y_4_c19 <= Y_4_c18;
               Y_5_c19 <= Y_5_c18;
               Y_6_c19 <= Y_6_c18;
               Y_7_c19 <= Y_7_c18;
               Y_8_c19 <= Y_8_c18;
               Y_9_c19 <= Y_9_c18;
               Y_10_c19 <= Y_10_c18;
               Y_11_c19 <= Y_11_c18;
               Y_12_c19 <= Y_12_c18;
            end if;
            if ce_20 = '1' then
               Y_1_c20 <= Y_1_c19;
               Y_2_c20 <= Y_2_c19;
               Y_3_c20 <= Y_3_c19;
               Y_4_c20 <= Y_4_c19;
               Y_5_c20 <= Y_5_c19;
               Y_6_c20 <= Y_6_c19;
               Y_7_c20 <= Y_7_c19;
               Y_8_c20 <= Y_8_c19;
               Y_9_c20 <= Y_9_c19;
               Y_10_c20 <= Y_10_c19;
               Y_11_c20 <= Y_11_c19;
               Y_12_c20 <= Y_12_c19;
            end if;
            if ce_21 = '1' then
               Y_1_c21 <= Y_1_c20;
               Y_2_c21 <= Y_2_c20;
               Y_3_c21 <= Y_3_c20;
               Y_4_c21 <= Y_4_c20;
               Y_5_c21 <= Y_5_c20;
               Y_6_c21 <= Y_6_c20;
               Y_7_c21 <= Y_7_c20;
               Y_8_c21 <= Y_8_c20;
               Y_9_c21 <= Y_9_c20;
               Y_10_c21 <= Y_10_c20;
               Y_11_c21 <= Y_11_c20;
               Y_12_c21 <= Y_12_c20;
            end if;
            if ce_22 = '1' then
               Y_1_c22 <= Y_1_c21;
               Y_2_c22 <= Y_2_c21;
               Y_3_c22 <= Y_3_c21;
               Y_4_c22 <= Y_4_c21;
               Y_5_c22 <= Y_5_c21;
               Y_6_c22 <= Y_6_c21;
               Y_7_c22 <= Y_7_c21;
               Y_8_c22 <= Y_8_c21;
               Y_9_c22 <= Y_9_c21;
               Y_10_c22 <= Y_10_c21;
               Y_11_c22 <= Y_11_c21;
               Y_12_c22 <= Y_12_c21;
            end if;
            if ce_23 = '1' then
               Y_1_c23 <= Y_1_c22;
               Y_2_c23 <= Y_2_c22;
               Y_3_c23 <= Y_3_c22;
               Y_4_c23 <= Y_4_c22;
               Y_5_c23 <= Y_5_c22;
               Y_6_c23 <= Y_6_c22;
               Y_7_c23 <= Y_7_c22;
               Y_8_c23 <= Y_8_c22;
               Y_9_c23 <= Y_9_c22;
               Y_10_c23 <= Y_10_c22;
               Y_11_c23 <= Y_11_c22;
               Y_12_c23 <= Y_12_c22;
            end if;
            if ce_24 = '1' then
               Cin_1_c24 <= Cin_1_c23;
               X_1_c24 <= X_1_c23;
               Y_1_c24 <= Y_1_c23;
               X_2_c24 <= X_2_c23;
               Y_2_c24 <= Y_2_c23;
               X_3_c24 <= X_3_c23;
               Y_3_c24 <= Y_3_c23;
               X_4_c24 <= X_4_c23;
               Y_4_c24 <= Y_4_c23;
               X_5_c24 <= X_5_c23;
               Y_5_c24 <= Y_5_c23;
               X_6_c24 <= X_6_c23;
               Y_6_c24 <= Y_6_c23;
               X_7_c24 <= X_7_c23;
               Y_7_c24 <= Y_7_c23;
               X_8_c24 <= X_8_c23;
               Y_8_c24 <= Y_8_c23;
               X_9_c24 <= X_9_c23;
               Y_9_c24 <= Y_9_c23;
               X_10_c24 <= X_10_c23;
               Y_10_c24 <= Y_10_c23;
               X_11_c24 <= X_11_c23;
               Y_11_c24 <= Y_11_c23;
               X_12_c24 <= X_12_c23;
               Y_12_c24 <= Y_12_c23;
            end if;
            if ce_25 = '1' then
               R_1_c25 <= R_1_c24;
               Cin_2_c25 <= Cin_2_c24;
               X_2_c25 <= X_2_c24;
               Y_2_c25 <= Y_2_c24;
               X_3_c25 <= X_3_c24;
               Y_3_c25 <= Y_3_c24;
               X_4_c25 <= X_4_c24;
               Y_4_c25 <= Y_4_c24;
               X_5_c25 <= X_5_c24;
               Y_5_c25 <= Y_5_c24;
               X_6_c25 <= X_6_c24;
               Y_6_c25 <= Y_6_c24;
               X_7_c25 <= X_7_c24;
               Y_7_c25 <= Y_7_c24;
               X_8_c25 <= X_8_c24;
               Y_8_c25 <= Y_8_c24;
               X_9_c25 <= X_9_c24;
               Y_9_c25 <= Y_9_c24;
               X_10_c25 <= X_10_c24;
               Y_10_c25 <= Y_10_c24;
               X_11_c25 <= X_11_c24;
               Y_11_c25 <= Y_11_c24;
               X_12_c25 <= X_12_c24;
               Y_12_c25 <= Y_12_c24;
            end if;
            if ce_26 = '1' then
               R_1_c26 <= R_1_c25;
               R_2_c26 <= R_2_c25;
               Cin_3_c26 <= Cin_3_c25;
               X_3_c26 <= X_3_c25;
               Y_3_c26 <= Y_3_c25;
               X_4_c26 <= X_4_c25;
               Y_4_c26 <= Y_4_c25;
               X_5_c26 <= X_5_c25;
               Y_5_c26 <= Y_5_c25;
               X_6_c26 <= X_6_c25;
               Y_6_c26 <= Y_6_c25;
               X_7_c26 <= X_7_c25;
               Y_7_c26 <= Y_7_c25;
               X_8_c26 <= X_8_c25;
               Y_8_c26 <= Y_8_c25;
               X_9_c26 <= X_9_c25;
               Y_9_c26 <= Y_9_c25;
               X_10_c26 <= X_10_c25;
               Y_10_c26 <= Y_10_c25;
               X_11_c26 <= X_11_c25;
               Y_11_c26 <= Y_11_c25;
               X_12_c26 <= X_12_c25;
               Y_12_c26 <= Y_12_c25;
            end if;
            if ce_27 = '1' then
               R_1_c27 <= R_1_c26;
               R_2_c27 <= R_2_c26;
               R_3_c27 <= R_3_c26;
               Cin_4_c27 <= Cin_4_c26;
               X_4_c27 <= X_4_c26;
               Y_4_c27 <= Y_4_c26;
               X_5_c27 <= X_5_c26;
               Y_5_c27 <= Y_5_c26;
               X_6_c27 <= X_6_c26;
               Y_6_c27 <= Y_6_c26;
               X_7_c27 <= X_7_c26;
               Y_7_c27 <= Y_7_c26;
               X_8_c27 <= X_8_c26;
               Y_8_c27 <= Y_8_c26;
               X_9_c27 <= X_9_c26;
               Y_9_c27 <= Y_9_c26;
               X_10_c27 <= X_10_c26;
               Y_10_c27 <= Y_10_c26;
               X_11_c27 <= X_11_c26;
               Y_11_c27 <= Y_11_c26;
               X_12_c27 <= X_12_c26;
               Y_12_c27 <= Y_12_c26;
            end if;
            if ce_28 = '1' then
               R_1_c28 <= R_1_c27;
               R_2_c28 <= R_2_c27;
               R_3_c28 <= R_3_c27;
               R_4_c28 <= R_4_c27;
               Cin_5_c28 <= Cin_5_c27;
               X_5_c28 <= X_5_c27;
               Y_5_c28 <= Y_5_c27;
               X_6_c28 <= X_6_c27;
               Y_6_c28 <= Y_6_c27;
               X_7_c28 <= X_7_c27;
               Y_7_c28 <= Y_7_c27;
               X_8_c28 <= X_8_c27;
               Y_8_c28 <= Y_8_c27;
               X_9_c28 <= X_9_c27;
               Y_9_c28 <= Y_9_c27;
               X_10_c28 <= X_10_c27;
               Y_10_c28 <= Y_10_c27;
               X_11_c28 <= X_11_c27;
               Y_11_c28 <= Y_11_c27;
               X_12_c28 <= X_12_c27;
               Y_12_c28 <= Y_12_c27;
            end if;
            if ce_29 = '1' then
               R_1_c29 <= R_1_c28;
               R_2_c29 <= R_2_c28;
               R_3_c29 <= R_3_c28;
               R_4_c29 <= R_4_c28;
               R_5_c29 <= R_5_c28;
               Cin_6_c29 <= Cin_6_c28;
               X_6_c29 <= X_6_c28;
               Y_6_c29 <= Y_6_c28;
               X_7_c29 <= X_7_c28;
               Y_7_c29 <= Y_7_c28;
               X_8_c29 <= X_8_c28;
               Y_8_c29 <= Y_8_c28;
               X_9_c29 <= X_9_c28;
               Y_9_c29 <= Y_9_c28;
               X_10_c29 <= X_10_c28;
               Y_10_c29 <= Y_10_c28;
               X_11_c29 <= X_11_c28;
               Y_11_c29 <= Y_11_c28;
               X_12_c29 <= X_12_c28;
               Y_12_c29 <= Y_12_c28;
            end if;
            if ce_30 = '1' then
               R_1_c30 <= R_1_c29;
               R_2_c30 <= R_2_c29;
               R_3_c30 <= R_3_c29;
               R_4_c30 <= R_4_c29;
               R_5_c30 <= R_5_c29;
               R_6_c30 <= R_6_c29;
               Cin_7_c30 <= Cin_7_c29;
               X_7_c30 <= X_7_c29;
               Y_7_c30 <= Y_7_c29;
               X_8_c30 <= X_8_c29;
               Y_8_c30 <= Y_8_c29;
               X_9_c30 <= X_9_c29;
               Y_9_c30 <= Y_9_c29;
               X_10_c30 <= X_10_c29;
               Y_10_c30 <= Y_10_c29;
               X_11_c30 <= X_11_c29;
               Y_11_c30 <= Y_11_c29;
               X_12_c30 <= X_12_c29;
               Y_12_c30 <= Y_12_c29;
            end if;
            if ce_31 = '1' then
               R_1_c31 <= R_1_c30;
               R_2_c31 <= R_2_c30;
               R_3_c31 <= R_3_c30;
               R_4_c31 <= R_4_c30;
               R_5_c31 <= R_5_c30;
               R_6_c31 <= R_6_c30;
               R_7_c31 <= R_7_c30;
               Cin_8_c31 <= Cin_8_c30;
               X_8_c31 <= X_8_c30;
               Y_8_c31 <= Y_8_c30;
               X_9_c31 <= X_9_c30;
               Y_9_c31 <= Y_9_c30;
               X_10_c31 <= X_10_c30;
               Y_10_c31 <= Y_10_c30;
               X_11_c31 <= X_11_c30;
               Y_11_c31 <= Y_11_c30;
               X_12_c31 <= X_12_c30;
               Y_12_c31 <= Y_12_c30;
            end if;
            if ce_32 = '1' then
               R_1_c32 <= R_1_c31;
               R_2_c32 <= R_2_c31;
               R_3_c32 <= R_3_c31;
               R_4_c32 <= R_4_c31;
               R_5_c32 <= R_5_c31;
               R_6_c32 <= R_6_c31;
               R_7_c32 <= R_7_c31;
               R_8_c32 <= R_8_c31;
               Cin_9_c32 <= Cin_9_c31;
               X_9_c32 <= X_9_c31;
               Y_9_c32 <= Y_9_c31;
               X_10_c32 <= X_10_c31;
               Y_10_c32 <= Y_10_c31;
               X_11_c32 <= X_11_c31;
               Y_11_c32 <= Y_11_c31;
               X_12_c32 <= X_12_c31;
               Y_12_c32 <= Y_12_c31;
            end if;
            if ce_33 = '1' then
               R_1_c33 <= R_1_c32;
               R_2_c33 <= R_2_c32;
               R_3_c33 <= R_3_c32;
               R_4_c33 <= R_4_c32;
               R_5_c33 <= R_5_c32;
               R_6_c33 <= R_6_c32;
               R_7_c33 <= R_7_c32;
               R_8_c33 <= R_8_c32;
               R_9_c33 <= R_9_c32;
               Cin_10_c33 <= Cin_10_c32;
               X_10_c33 <= X_10_c32;
               Y_10_c33 <= Y_10_c32;
               X_11_c33 <= X_11_c32;
               Y_11_c33 <= Y_11_c32;
               X_12_c33 <= X_12_c32;
               Y_12_c33 <= Y_12_c32;
            end if;
            if ce_34 = '1' then
               R_1_c34 <= R_1_c33;
               R_2_c34 <= R_2_c33;
               R_3_c34 <= R_3_c33;
               R_4_c34 <= R_4_c33;
               R_5_c34 <= R_5_c33;
               R_6_c34 <= R_6_c33;
               R_7_c34 <= R_7_c33;
               R_8_c34 <= R_8_c33;
               R_9_c34 <= R_9_c33;
               R_10_c34 <= R_10_c33;
               Cin_11_c34 <= Cin_11_c33;
               X_11_c34 <= X_11_c33;
               Y_11_c34 <= Y_11_c33;
               X_12_c34 <= X_12_c33;
               Y_12_c34 <= Y_12_c33;
            end if;
            if ce_35 = '1' then
               R_1_c35 <= R_1_c34;
               R_2_c35 <= R_2_c34;
               R_3_c35 <= R_3_c34;
               R_4_c35 <= R_4_c34;
               R_5_c35 <= R_5_c34;
               R_6_c35 <= R_6_c34;
               R_7_c35 <= R_7_c34;
               R_8_c35 <= R_8_c34;
               R_9_c35 <= R_9_c34;
               R_10_c35 <= R_10_c34;
               R_11_c35 <= R_11_c34;
               Cin_12_c35 <= Cin_12_c34;
               X_12_c35 <= X_12_c34;
               Y_12_c35 <= Y_12_c34;
            end if;
         end if;
      end process;
   Cin_1_c23 <= Cin;
   X_1_c23 <= '0' & X(2 downto 0);
   Y_1_c0 <= '0' & Y(2 downto 0);
   S_1_c24 <= X_1_c24 + Y_1_c24 + Cin_1_c24;
   R_1_c24 <= S_1_c24(2 downto 0);
   Cin_2_c24 <= S_1_c24(3);
   X_2_c23 <= '0' & X(5 downto 3);
   Y_2_c0 <= '0' & Y(5 downto 3);
   S_2_c25 <= X_2_c25 + Y_2_c25 + Cin_2_c25;
   R_2_c25 <= S_2_c25(2 downto 0);
   Cin_3_c25 <= S_2_c25(3);
   X_3_c23 <= '0' & X(8 downto 6);
   Y_3_c0 <= '0' & Y(8 downto 6);
   S_3_c26 <= X_3_c26 + Y_3_c26 + Cin_3_c26;
   R_3_c26 <= S_3_c26(2 downto 0);
   Cin_4_c26 <= S_3_c26(3);
   X_4_c23 <= '0' & X(11 downto 9);
   Y_4_c0 <= '0' & Y(11 downto 9);
   S_4_c27 <= X_4_c27 + Y_4_c27 + Cin_4_c27;
   R_4_c27 <= S_4_c27(2 downto 0);
   Cin_5_c27 <= S_4_c27(3);
   X_5_c23 <= '0' & X(14 downto 12);
   Y_5_c0 <= '0' & Y(14 downto 12);
   S_5_c28 <= X_5_c28 + Y_5_c28 + Cin_5_c28;
   R_5_c28 <= S_5_c28(2 downto 0);
   Cin_6_c28 <= S_5_c28(3);
   X_6_c23 <= '0' & X(17 downto 15);
   Y_6_c0 <= '0' & Y(17 downto 15);
   S_6_c29 <= X_6_c29 + Y_6_c29 + Cin_6_c29;
   R_6_c29 <= S_6_c29(2 downto 0);
   Cin_7_c29 <= S_6_c29(3);
   X_7_c23 <= '0' & X(20 downto 18);
   Y_7_c0 <= '0' & Y(20 downto 18);
   S_7_c30 <= X_7_c30 + Y_7_c30 + Cin_7_c30;
   R_7_c30 <= S_7_c30(2 downto 0);
   Cin_8_c30 <= S_7_c30(3);
   X_8_c23 <= '0' & X(23 downto 21);
   Y_8_c0 <= '0' & Y(23 downto 21);
   S_8_c31 <= X_8_c31 + Y_8_c31 + Cin_8_c31;
   R_8_c31 <= S_8_c31(2 downto 0);
   Cin_9_c31 <= S_8_c31(3);
   X_9_c23 <= '0' & X(26 downto 24);
   Y_9_c0 <= '0' & Y(26 downto 24);
   S_9_c32 <= X_9_c32 + Y_9_c32 + Cin_9_c32;
   R_9_c32 <= S_9_c32(2 downto 0);
   Cin_10_c32 <= S_9_c32(3);
   X_10_c23 <= '0' & X(29 downto 27);
   Y_10_c0 <= '0' & Y(29 downto 27);
   S_10_c33 <= X_10_c33 + Y_10_c33 + Cin_10_c33;
   R_10_c33 <= S_10_c33(2 downto 0);
   Cin_11_c33 <= S_10_c33(3);
   X_11_c23 <= '0' & X(32 downto 30);
   Y_11_c0 <= '0' & Y(32 downto 30);
   S_11_c34 <= X_11_c34 + Y_11_c34 + Cin_11_c34;
   R_11_c34 <= S_11_c34(2 downto 0);
   Cin_12_c34 <= S_11_c34(3);
   X_12_c23 <= '0' & X(33 downto 33);
   Y_12_c0 <= '0' & Y(33 downto 33);
   S_12_c35 <= X_12_c35 + Y_12_c35 + Cin_12_c35;
   R_12_c35 <= S_12_c35(0 downto 0);
   R <= R_12_c35 & R_11_c35 & R_10_c35 & R_9_c35 & R_8_c35 & R_7_c35 & R_6_c35 & R_5_c35 & R_4_c35 & R_3_c35 & R_2_c35 & R_1_c35 ;
end architecture;

--------------------------------------------------------------------------------
--                             FloatingPointAdder
--                         (FPAdd_8_23_Freq800_uid2)
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2010-2017)
--------------------------------------------------------------------------------
-- Pipeline depth: 36 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointAdder_32_2_798000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointAdder_32_2_798000 is
   component RightShifterSticky24_by_max_26_Freq800_uid4 is
      port ( clk, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8 : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(25 downto 0);
             Sticky : out  std_logic   );
   end component;

   component IntAdder_27_Freq800_uid6 is
      port ( clk, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17 : in std_logic;
             X : in  std_logic_vector(26 downto 0);
             Y : in  std_logic_vector(26 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(26 downto 0)   );
   end component;

   component Normalizer_Z_28_28_28_Freq800_uid8 is
      port ( clk, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23 : in std_logic;
             X : in  std_logic_vector(27 downto 0);
             Count : out  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_Freq800_uid11 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35 : in std_logic;
             X : in  std_logic_vector(33 downto 0);
             Y : in  std_logic_vector(33 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX_c0, excExpFracX_c1 :  std_logic_vector(32 downto 0);
signal excExpFracY_c0, excExpFracY_c1 :  std_logic_vector(32 downto 0);
signal swap_c1 :  std_logic;
signal eXmeY_c1 :  std_logic_vector(7 downto 0);
signal eYmeX_c1 :  std_logic_vector(7 downto 0);
signal expDiff_c1, expDiff_c2 :  std_logic_vector(7 downto 0);
signal newX_c1 :  std_logic_vector(33 downto 0);
signal newY_c1, newY_c2 :  std_logic_vector(33 downto 0);
signal expX_c1, expX_c2 :  std_logic_vector(7 downto 0);
signal excX_c1 :  std_logic_vector(1 downto 0);
signal excY_c1, excY_c2 :  std_logic_vector(1 downto 0);
signal signX_c1, signX_c2 :  std_logic;
signal signY_c1, signY_c2 :  std_logic;
signal EffSub_c2, EffSub_c3, EffSub_c4, EffSub_c5, EffSub_c6, EffSub_c7, EffSub_c8, EffSub_c9, EffSub_c10, EffSub_c11, EffSub_c12, EffSub_c13, EffSub_c14, EffSub_c15, EffSub_c16, EffSub_c17, EffSub_c18, EffSub_c19, EffSub_c20, EffSub_c21, EffSub_c22, EffSub_c23, EffSub_c24, EffSub_c25, EffSub_c26, EffSub_c27, EffSub_c28, EffSub_c29, EffSub_c30, EffSub_c31, EffSub_c32, EffSub_c33, EffSub_c34, EffSub_c35, EffSub_c36 :  std_logic;
signal sXsYExnXY_c1, sXsYExnXY_c2 :  std_logic_vector(5 downto 0);
signal sdExnXY_c1 :  std_logic_vector(3 downto 0);
signal fracY_c2 :  std_logic_vector(23 downto 0);
signal excRt_c2, excRt_c3, excRt_c4, excRt_c5, excRt_c6, excRt_c7, excRt_c8, excRt_c9, excRt_c10, excRt_c11, excRt_c12, excRt_c13, excRt_c14, excRt_c15, excRt_c16, excRt_c17, excRt_c18, excRt_c19, excRt_c20, excRt_c21, excRt_c22, excRt_c23, excRt_c24, excRt_c25, excRt_c26, excRt_c27, excRt_c28, excRt_c29, excRt_c30, excRt_c31, excRt_c32, excRt_c33, excRt_c34, excRt_c35, excRt_c36 :  std_logic_vector(1 downto 0);
signal signR_c2, signR_c3, signR_c4, signR_c5, signR_c6, signR_c7, signR_c8, signR_c9, signR_c10, signR_c11, signR_c12, signR_c13, signR_c14, signR_c15, signR_c16, signR_c17, signR_c18, signR_c19, signR_c20, signR_c21, signR_c22, signR_c23 :  std_logic;
signal shiftedOut_c2 :  std_logic;
signal shiftVal_c2 :  std_logic_vector(4 downto 0);
signal shiftedFracY_c3 :  std_logic_vector(25 downto 0);
signal sticky_c8, sticky_c9, sticky_c10, sticky_c11, sticky_c12, sticky_c13, sticky_c14, sticky_c15, sticky_c16, sticky_c17 :  std_logic;
signal fracYpad_c3, fracYpad_c4 :  std_logic_vector(26 downto 0);
signal EffSubVector_c2, EffSubVector_c3, EffSubVector_c4 :  std_logic_vector(26 downto 0);
signal fracYpadXorOp_c4 :  std_logic_vector(26 downto 0);
signal fracXpad_c1 :  std_logic_vector(26 downto 0);
signal cInSigAdd_c8 :  std_logic;
signal fracAddResult_c17 :  std_logic_vector(26 downto 0);
signal fracSticky_c17 :  std_logic_vector(27 downto 0);
signal nZerosNew_c22, nZerosNew_c23 :  std_logic_vector(4 downto 0);
signal shiftedFrac_c23 :  std_logic_vector(27 downto 0);
signal extendedExpInc_c2, extendedExpInc_c3, extendedExpInc_c4, extendedExpInc_c5, extendedExpInc_c6, extendedExpInc_c7, extendedExpInc_c8, extendedExpInc_c9, extendedExpInc_c10, extendedExpInc_c11, extendedExpInc_c12, extendedExpInc_c13, extendedExpInc_c14, extendedExpInc_c15, extendedExpInc_c16, extendedExpInc_c17, extendedExpInc_c18, extendedExpInc_c19, extendedExpInc_c20, extendedExpInc_c21, extendedExpInc_c22, extendedExpInc_c23 :  std_logic_vector(8 downto 0);
signal updatedExp_c23 :  std_logic_vector(9 downto 0);
signal eqdiffsign_c22, eqdiffsign_c23, eqdiffsign_c24, eqdiffsign_c25, eqdiffsign_c26, eqdiffsign_c27, eqdiffsign_c28, eqdiffsign_c29, eqdiffsign_c30, eqdiffsign_c31, eqdiffsign_c32, eqdiffsign_c33, eqdiffsign_c34, eqdiffsign_c35, eqdiffsign_c36 :  std_logic;
signal expFrac_c23 :  std_logic_vector(33 downto 0);
signal stk_c23 :  std_logic;
signal rnd_c23 :  std_logic;
signal lsb_c23 :  std_logic;
signal needToRound_c23 :  std_logic;
signal RoundedExpFrac_c35 :  std_logic_vector(33 downto 0);
signal upExc_c35 :  std_logic_vector(1 downto 0);
signal fracR_c35, fracR_c36 :  std_logic_vector(22 downto 0);
signal expR_c35, expR_c36 :  std_logic_vector(7 downto 0);
signal exExpExc_c35, exExpExc_c36 :  std_logic_vector(3 downto 0);
signal excRt2_c36 :  std_logic_vector(1 downto 0);
signal excR_c36 :  std_logic_vector(1 downto 0);
signal signR2_c23, signR2_c24, signR2_c25, signR2_c26, signR2_c27, signR2_c28, signR2_c29, signR2_c30, signR2_c31, signR2_c32, signR2_c33, signR2_c34, signR2_c35, signR2_c36 :  std_logic;
signal computedR_c36 :  std_logic_vector(33 downto 0);
signal X_c1 :  std_logic_vector(8+23+2 downto 0);
signal Y_c1 :  std_logic_vector(8+23+2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               excExpFracX_c1 <= excExpFracX_c0;
               excExpFracY_c1 <= excExpFracY_c0;
               X_c1 <= X;
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               expDiff_c2 <= expDiff_c1;
               newY_c2 <= newY_c1;
               expX_c2 <= expX_c1;
               excY_c2 <= excY_c1;
               signX_c2 <= signX_c1;
               signY_c2 <= signY_c1;
               sXsYExnXY_c2 <= sXsYExnXY_c1;
            end if;
            if ce_3 = '1' then
               EffSub_c3 <= EffSub_c2;
               excRt_c3 <= excRt_c2;
               signR_c3 <= signR_c2;
               EffSubVector_c3 <= EffSubVector_c2;
               extendedExpInc_c3 <= extendedExpInc_c2;
            end if;
            if ce_4 = '1' then
               EffSub_c4 <= EffSub_c3;
               excRt_c4 <= excRt_c3;
               signR_c4 <= signR_c3;
               fracYpad_c4 <= fracYpad_c3;
               EffSubVector_c4 <= EffSubVector_c3;
               extendedExpInc_c4 <= extendedExpInc_c3;
            end if;
            if ce_5 = '1' then
               EffSub_c5 <= EffSub_c4;
               excRt_c5 <= excRt_c4;
               signR_c5 <= signR_c4;
               extendedExpInc_c5 <= extendedExpInc_c4;
            end if;
            if ce_6 = '1' then
               EffSub_c6 <= EffSub_c5;
               excRt_c6 <= excRt_c5;
               signR_c6 <= signR_c5;
               extendedExpInc_c6 <= extendedExpInc_c5;
            end if;
            if ce_7 = '1' then
               EffSub_c7 <= EffSub_c6;
               excRt_c7 <= excRt_c6;
               signR_c7 <= signR_c6;
               extendedExpInc_c7 <= extendedExpInc_c6;
            end if;
            if ce_8 = '1' then
               EffSub_c8 <= EffSub_c7;
               excRt_c8 <= excRt_c7;
               signR_c8 <= signR_c7;
               extendedExpInc_c8 <= extendedExpInc_c7;
            end if;
            if ce_9 = '1' then
               EffSub_c9 <= EffSub_c8;
               excRt_c9 <= excRt_c8;
               signR_c9 <= signR_c8;
               sticky_c9 <= sticky_c8;
               extendedExpInc_c9 <= extendedExpInc_c8;
            end if;
            if ce_10 = '1' then
               EffSub_c10 <= EffSub_c9;
               excRt_c10 <= excRt_c9;
               signR_c10 <= signR_c9;
               sticky_c10 <= sticky_c9;
               extendedExpInc_c10 <= extendedExpInc_c9;
            end if;
            if ce_11 = '1' then
               EffSub_c11 <= EffSub_c10;
               excRt_c11 <= excRt_c10;
               signR_c11 <= signR_c10;
               sticky_c11 <= sticky_c10;
               extendedExpInc_c11 <= extendedExpInc_c10;
            end if;
            if ce_12 = '1' then
               EffSub_c12 <= EffSub_c11;
               excRt_c12 <= excRt_c11;
               signR_c12 <= signR_c11;
               sticky_c12 <= sticky_c11;
               extendedExpInc_c12 <= extendedExpInc_c11;
            end if;
            if ce_13 = '1' then
               EffSub_c13 <= EffSub_c12;
               excRt_c13 <= excRt_c12;
               signR_c13 <= signR_c12;
               sticky_c13 <= sticky_c12;
               extendedExpInc_c13 <= extendedExpInc_c12;
            end if;
            if ce_14 = '1' then
               EffSub_c14 <= EffSub_c13;
               excRt_c14 <= excRt_c13;
               signR_c14 <= signR_c13;
               sticky_c14 <= sticky_c13;
               extendedExpInc_c14 <= extendedExpInc_c13;
            end if;
            if ce_15 = '1' then
               EffSub_c15 <= EffSub_c14;
               excRt_c15 <= excRt_c14;
               signR_c15 <= signR_c14;
               sticky_c15 <= sticky_c14;
               extendedExpInc_c15 <= extendedExpInc_c14;
            end if;
            if ce_16 = '1' then
               EffSub_c16 <= EffSub_c15;
               excRt_c16 <= excRt_c15;
               signR_c16 <= signR_c15;
               sticky_c16 <= sticky_c15;
               extendedExpInc_c16 <= extendedExpInc_c15;
            end if;
            if ce_17 = '1' then
               EffSub_c17 <= EffSub_c16;
               excRt_c17 <= excRt_c16;
               signR_c17 <= signR_c16;
               sticky_c17 <= sticky_c16;
               extendedExpInc_c17 <= extendedExpInc_c16;
            end if;
            if ce_18 = '1' then
               EffSub_c18 <= EffSub_c17;
               excRt_c18 <= excRt_c17;
               signR_c18 <= signR_c17;
               extendedExpInc_c18 <= extendedExpInc_c17;
            end if;
            if ce_19 = '1' then
               EffSub_c19 <= EffSub_c18;
               excRt_c19 <= excRt_c18;
               signR_c19 <= signR_c18;
               extendedExpInc_c19 <= extendedExpInc_c18;
            end if;
            if ce_20 = '1' then
               EffSub_c20 <= EffSub_c19;
               excRt_c20 <= excRt_c19;
               signR_c20 <= signR_c19;
               extendedExpInc_c20 <= extendedExpInc_c19;
            end if;
            if ce_21 = '1' then
               EffSub_c21 <= EffSub_c20;
               excRt_c21 <= excRt_c20;
               signR_c21 <= signR_c20;
               extendedExpInc_c21 <= extendedExpInc_c20;
            end if;
            if ce_22 = '1' then
               EffSub_c22 <= EffSub_c21;
               excRt_c22 <= excRt_c21;
               signR_c22 <= signR_c21;
               extendedExpInc_c22 <= extendedExpInc_c21;
            end if;
            if ce_23 = '1' then
               EffSub_c23 <= EffSub_c22;
               excRt_c23 <= excRt_c22;
               signR_c23 <= signR_c22;
               nZerosNew_c23 <= nZerosNew_c22;
               extendedExpInc_c23 <= extendedExpInc_c22;
               eqdiffsign_c23 <= eqdiffsign_c22;
            end if;
            if ce_24 = '1' then
               EffSub_c24 <= EffSub_c23;
               excRt_c24 <= excRt_c23;
               eqdiffsign_c24 <= eqdiffsign_c23;
               signR2_c24 <= signR2_c23;
            end if;
            if ce_25 = '1' then
               EffSub_c25 <= EffSub_c24;
               excRt_c25 <= excRt_c24;
               eqdiffsign_c25 <= eqdiffsign_c24;
               signR2_c25 <= signR2_c24;
            end if;
            if ce_26 = '1' then
               EffSub_c26 <= EffSub_c25;
               excRt_c26 <= excRt_c25;
               eqdiffsign_c26 <= eqdiffsign_c25;
               signR2_c26 <= signR2_c25;
            end if;
            if ce_27 = '1' then
               EffSub_c27 <= EffSub_c26;
               excRt_c27 <= excRt_c26;
               eqdiffsign_c27 <= eqdiffsign_c26;
               signR2_c27 <= signR2_c26;
            end if;
            if ce_28 = '1' then
               EffSub_c28 <= EffSub_c27;
               excRt_c28 <= excRt_c27;
               eqdiffsign_c28 <= eqdiffsign_c27;
               signR2_c28 <= signR2_c27;
            end if;
            if ce_29 = '1' then
               EffSub_c29 <= EffSub_c28;
               excRt_c29 <= excRt_c28;
               eqdiffsign_c29 <= eqdiffsign_c28;
               signR2_c29 <= signR2_c28;
            end if;
            if ce_30 = '1' then
               EffSub_c30 <= EffSub_c29;
               excRt_c30 <= excRt_c29;
               eqdiffsign_c30 <= eqdiffsign_c29;
               signR2_c30 <= signR2_c29;
            end if;
            if ce_31 = '1' then
               EffSub_c31 <= EffSub_c30;
               excRt_c31 <= excRt_c30;
               eqdiffsign_c31 <= eqdiffsign_c30;
               signR2_c31 <= signR2_c30;
            end if;
            if ce_32 = '1' then
               EffSub_c32 <= EffSub_c31;
               excRt_c32 <= excRt_c31;
               eqdiffsign_c32 <= eqdiffsign_c31;
               signR2_c32 <= signR2_c31;
            end if;
            if ce_33 = '1' then
               EffSub_c33 <= EffSub_c32;
               excRt_c33 <= excRt_c32;
               eqdiffsign_c33 <= eqdiffsign_c32;
               signR2_c33 <= signR2_c32;
            end if;
            if ce_34 = '1' then
               EffSub_c34 <= EffSub_c33;
               excRt_c34 <= excRt_c33;
               eqdiffsign_c34 <= eqdiffsign_c33;
               signR2_c34 <= signR2_c33;
            end if;
            if ce_35 = '1' then
               EffSub_c35 <= EffSub_c34;
               excRt_c35 <= excRt_c34;
               eqdiffsign_c35 <= eqdiffsign_c34;
               signR2_c35 <= signR2_c34;
            end if;
            if ce_36 = '1' then
               EffSub_c36 <= EffSub_c35;
               excRt_c36 <= excRt_c35;
               eqdiffsign_c36 <= eqdiffsign_c35;
               fracR_c36 <= fracR_c35;
               expR_c36 <= expR_c35;
               exExpExc_c36 <= exExpExc_c35;
               signR2_c36 <= signR2_c35;
            end if;
         end if;
      end process;
   excExpFracX_c0 <= X(33 downto 32) & X(30 downto 0);
   excExpFracY_c0 <= Y(33 downto 32) & Y(30 downto 0);
   swap_c1 <= '1' when excExpFracX_c1 < excExpFracY_c1 else '0';
   -- exponent difference
   eXmeY_c1 <= (X_c1(30 downto 23)) - (Y_c1(30 downto 23));
   eYmeX_c1 <= (Y_c1(30 downto 23)) - (X_c1(30 downto 23));
   expDiff_c1 <= eXmeY_c1 when swap_c1 = '0' else eYmeX_c1;
   -- input swap so that |X|>|Y|
   newX_c1 <= X_c1 when swap_c1 = '0' else Y_c1;
   newY_c1 <= Y_c1 when swap_c1 = '0' else X_c1;
   -- now we decompose the inputs into their sign, exponent, fraction
   expX_c1<= newX_c1(30 downto 23);
   excX_c1<= newX_c1(33 downto 32);
   excY_c1<= newY_c1(33 downto 32);
   signX_c1<= newX_c1(31);
   signY_c1<= newY_c1(31);
   EffSub_c2 <= signX_c2 xor signY_c2;
   sXsYExnXY_c1 <= signX_c1 & signY_c1 & excX_c1 & excY_c1;
   sdExnXY_c1 <= excX_c1 & excY_c1;
   fracY_c2 <= "000000000000000000000000" when excY_c2="00" else ('1' & newY_c2(22 downto 0));
   -- Exception management logic
   with sXsYExnXY_c2  select  
   excRt_c2 <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR_c2<= '0' when (sXsYExnXY_c2="100000" or sXsYExnXY_c2="010000") else signX_c2;
   shiftedOut_c2 <= '1' when (expDiff_c2 > 25) else '0';
   shiftVal_c2 <= expDiff_c2(4 downto 0) when shiftedOut_c2='0' else CONV_STD_LOGIC_VECTOR(26,5);
   RightShifterComponent: RightShifterSticky24_by_max_26_Freq800_uid4
      port map ( clk  => clk,
                 ce_3 => ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 S => shiftVal_c2,
                 X => fracY_c2,
                 R => shiftedFracY_c3,
                 Sticky => sticky_c8);
   fracYpad_c3 <= "0" & shiftedFracY_c3;
   EffSubVector_c2 <= (26 downto 0 => EffSub_c2);
   fracYpadXorOp_c4 <= fracYpad_c4 xor EffSubVector_c4;
   fracXpad_c1 <= "01" & (newX_c1(22 downto 0)) & "00";
   cInSigAdd_c8 <= EffSub_c8 and not sticky_c8; -- if we subtract and the sticky was one, some of the negated sticky bits would have absorbed this carry 
   fracAdder: IntAdder_27_Freq800_uid6
      port map ( clk  => clk,
                 ce_2 => ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 Cin => cInSigAdd_c8,
                 X => fracXpad_c1,
                 Y => fracYpadXorOp_c4,
                 R => fracAddResult_c17);
   fracSticky_c17<= fracAddResult_c17 & sticky_c17; 
   LZCAndShifter: Normalizer_Z_28_28_28_Freq800_uid8
      port map ( clk  => clk,
                 ce_18 => ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 X => fracSticky_c17,
                 Count => nZerosNew_c22,
                 R => shiftedFrac_c23);
   extendedExpInc_c2<= ("0" & expX_c2) + '1';
   updatedExp_c23 <= ("0" &extendedExpInc_c23) - ("00000" & nZerosNew_c23);
   eqdiffsign_c22 <= '1' when nZerosNew_c22="11111" else '0';
   expFrac_c23<= updatedExp_c23 & shiftedFrac_c23(26 downto 3);
   stk_c23<= shiftedFrac_c23(2) or shiftedFrac_c23(1) or shiftedFrac_c23(0);
   rnd_c23<= shiftedFrac_c23(3);
   lsb_c23<= shiftedFrac_c23(4);
   needToRound_c23<= '1' when (rnd_c23='1' and stk_c23='1') or (rnd_c23='1' and stk_c23='0' and lsb_c23='1')
  else '0';
   roundingAdder: IntAdder_34_Freq800_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 Cin => needToRound_c23,
                 X => expFrac_c23,
                 Y => "0000000000000000000000000000000000",
                 R => RoundedExpFrac_c35);
   -- possible update to exception bits
   upExc_c35 <= RoundedExpFrac_c35(33 downto 32);
   fracR_c35 <= RoundedExpFrac_c35(23 downto 1);
   expR_c35 <= RoundedExpFrac_c35(31 downto 24);
   exExpExc_c35 <= upExc_c35 & excRt_c35;
   with exExpExc_c36  select  
   excRt2_c36<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR_c36 <= "00" when (eqdiffsign_c36='1' and EffSub_c36='1'  and not(excRt_c36="11")) else excRt2_c36;
   signR2_c23 <= '0' when (eqdiffsign_c23='1' and EffSub_c23='1') else signR_c23;
   computedR_c36 <= excR_c36 & signR2_c36 & expR_c36 & fracR_c36;
   R <= computedR_c36;
end architecture;




--------------------------------------------------------------------------------
--                RightShifterSticky24_by_max_26_Freq500_uid4
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X S
-- Output signals: R Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifterSticky24_by_max_26_Freq500_uid4 is
    port (clk, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(25 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of RightShifterSticky24_by_max_26_Freq500_uid4 is
signal ps_c1, ps_c2, ps_c3, ps_c4 :  std_logic_vector(4 downto 0);
signal Xpadded_c1 :  std_logic_vector(25 downto 0);
signal level5_c1, level5_c2 :  std_logic_vector(25 downto 0);
signal stk4_c2 :  std_logic;
signal level4_c1, level4_c2 :  std_logic_vector(25 downto 0);
signal stk3_c2, stk3_c3 :  std_logic;
signal level3_c1, level3_c2, level3_c3 :  std_logic_vector(25 downto 0);
signal stk2_c3, stk2_c4 :  std_logic;
signal level2_c1, level2_c2, level2_c3, level2_c4 :  std_logic_vector(25 downto 0);
signal stk1_c4 :  std_logic;
signal level1_c2, level1_c3, level1_c4 :  std_logic_vector(25 downto 0);
signal stk0_c4 :  std_logic;
signal level0_c2 :  std_logic_vector(25 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_2 = '1' then
               ps_c2 <= ps_c1;
               level5_c2 <= level5_c1;
               level4_c2 <= level4_c1;
               level3_c2 <= level3_c1;
               level2_c2 <= level2_c1;
            end if;
            if ce_3 = '1' then
               ps_c3 <= ps_c2;
               stk3_c3 <= stk3_c2;
               level3_c3 <= level3_c2;
               level2_c3 <= level2_c2;
               level1_c3 <= level1_c2;
            end if;
            if ce_4 = '1' then
               ps_c4 <= ps_c3;
               stk2_c4 <= stk2_c3;
               level2_c4 <= level2_c3;
               level1_c4 <= level1_c3;
            end if;
         end if;
      end process;
   ps_c1<= S;
   Xpadded_c1 <= X&(1 downto 0 => '0');
   level5_c1<= Xpadded_c1;
   stk4_c2 <= '1' when (level5_c2(15 downto 0)/="0000000000000000" and ps_c2(4)='1')   else '0';
   level4_c1 <=  level5_c1 when  ps_c1(4)='0'    else (15 downto 0 => '0') & level5_c1(25 downto 16);
   stk3_c2 <= '1' when (level4_c2(7 downto 0)/="00000000" and ps_c2(3)='1') or stk4_c2 ='1'   else '0';
   level3_c1 <=  level4_c1 when  ps_c1(3)='0'    else (7 downto 0 => '0') & level4_c1(25 downto 8);
   stk2_c3 <= '1' when (level3_c3(3 downto 0)/="0000" and ps_c3(2)='1') or stk3_c3 ='1'   else '0';
   level2_c1 <=  level3_c1 when  ps_c1(2)='0'    else (3 downto 0 => '0') & level3_c1(25 downto 4);
   stk1_c4 <= '1' when (level2_c4(1 downto 0)/="00" and ps_c4(1)='1') or stk2_c4 ='1'   else '0';
   level1_c2 <=  level2_c2 when  ps_c2(1)='0'    else (1 downto 0 => '0') & level2_c2(25 downto 2);
   stk0_c4 <= '1' when (level1_c4(0 downto 0)/="0" and ps_c4(0)='1') or stk1_c4 ='1'   else '0';
   level0_c2 <=  level1_c2 when  ps_c2(0)='0'    else (0 downto 0 => '0') & level1_c2(25 downto 1);
   R <= level0_c2;
   Sticky <= stk0_c4;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_27_Freq500_uid6
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_Freq500_uid6 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5 : in std_logic;
          X : in  std_logic_vector(26 downto 0);
          Y : in  std_logic_vector(26 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_Freq500_uid6 is
signal Rtmp_c5 :  std_logic_vector(26 downto 0);
signal X_c1, X_c2, X_c3, X_c4, X_c5 :  std_logic_vector(26 downto 0);
signal Y_c3, Y_c4, Y_c5 :  std_logic_vector(26 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               X_c1 <= X;
            end if;
            if ce_2 = '1' then
               X_c2 <= X_c1;
            end if;
            if ce_3 = '1' then
               X_c3 <= X_c2;
               Y_c3 <= Y;
            end if;
            if ce_4 = '1' then
               X_c4 <= X_c3;
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               X_c5 <= X_c4;
               Y_c5 <= Y_c4;
            end if;
         end if;
      end process;
   Rtmp_c5 <= X_c5 + Y_c5 + Cin;
   R <= Rtmp_c5;
end architecture;

--------------------------------------------------------------------------------
--                     Normalizer_Z_28_28_28_Freq500_uid8
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_28_28_28_Freq500_uid8 is
    port (clk, ce_6, ce_7, ce_8 : in std_logic;
          X : in  std_logic_vector(27 downto 0);
          Count : out  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of Normalizer_Z_28_28_28_Freq500_uid8 is
signal level5_c5, level5_c6 :  std_logic_vector(27 downto 0);
signal count4_c6, count4_c7, count4_c8 :  std_logic;
signal level4_c6 :  std_logic_vector(27 downto 0);
signal count3_c6, count3_c7, count3_c8 :  std_logic;
signal level3_c6, level3_c7 :  std_logic_vector(27 downto 0);
signal count2_c7, count2_c8 :  std_logic;
signal level2_c7, level2_c8 :  std_logic_vector(27 downto 0);
signal count1_c7, count1_c8 :  std_logic;
signal level1_c8 :  std_logic_vector(27 downto 0);
signal count0_c8 :  std_logic;
signal level0_c8 :  std_logic_vector(27 downto 0);
signal sCount_c8 :  std_logic_vector(4 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_6 = '1' then
               level5_c6 <= level5_c5;
            end if;
            if ce_7 = '1' then
               count4_c7 <= count4_c6;
               count3_c7 <= count3_c6;
               level3_c7 <= level3_c6;
            end if;
            if ce_8 = '1' then
               count4_c8 <= count4_c7;
               count3_c8 <= count3_c7;
               count2_c8 <= count2_c7;
               level2_c8 <= level2_c7;
               count1_c8 <= count1_c7;
            end if;
         end if;
      end process;
   level5_c5 <= X ;
   count4_c6<= '1' when level5_c6(27 downto 12) = (27 downto 12=>'0') else '0';
   level4_c6<= level5_c6(27 downto 0) when count4_c6='0' else level5_c6(11 downto 0) & (15 downto 0 => '0');

   count3_c6<= '1' when level4_c6(27 downto 20) = (27 downto 20=>'0') else '0';
   level3_c6<= level4_c6(27 downto 0) when count3_c6='0' else level4_c6(19 downto 0) & (7 downto 0 => '0');

   count2_c7<= '1' when level3_c7(27 downto 24) = (27 downto 24=>'0') else '0';
   level2_c7<= level3_c7(27 downto 0) when count2_c7='0' else level3_c7(23 downto 0) & (3 downto 0 => '0');

   count1_c7<= '1' when level2_c7(27 downto 26) = (27 downto 26=>'0') else '0';
   level1_c8<= level2_c8(27 downto 0) when count1_c8='0' else level2_c8(25 downto 0) & (1 downto 0 => '0');

   count0_c8<= '1' when level1_c8(27 downto 27) = (27 downto 27=>'0') else '0';
   level0_c8<= level1_c8(27 downto 0) when count0_c8='0' else level1_c8(26 downto 0) & (0 downto 0 => '0');

   R <= level0_c8;
   sCount_c8 <= count4_c8 & count3_c8 & count2_c8 & count1_c8 & count0_c8;
   Count <= sCount_c8;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_Freq500_uid11
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_Freq500_uid11 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(33 downto 0);
          Y : in  std_logic_vector(33 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_Freq500_uid11 is
signal Rtmp_c9 :  std_logic_vector(33 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5, Y_c6, Y_c7, Y_c8, Y_c9 :  std_logic_vector(33 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
            if ce_6 = '1' then
               Y_c6 <= Y_c5;
            end if;
            if ce_7 = '1' then
               Y_c7 <= Y_c6;
            end if;
            if ce_8 = '1' then
               Y_c8 <= Y_c7;
            end if;
            if ce_9 = '1' then
               Y_c9 <= Y_c8;
            end if;
         end if;
      end process;
   Rtmp_c9 <= X + Y_c9 + Cin;
   R <= Rtmp_c9;
end architecture;

--------------------------------------------------------------------------------
--                             FloatingPointAdder
--                         (FPAdd_8_23_Freq500_uid2)
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2010-2017)
--------------------------------------------------------------------------------
-- Pipeline depth: 10 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointAdder_32_2_922000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointAdder_32_2_922000 is
   component RightShifterSticky24_by_max_26_Freq500_uid4 is
      port ( clk, ce_2, ce_3, ce_4 : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(25 downto 0);
             Sticky : out  std_logic   );
   end component;

   component IntAdder_27_Freq500_uid6 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5 : in std_logic;
             X : in  std_logic_vector(26 downto 0);
             Y : in  std_logic_vector(26 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(26 downto 0)   );
   end component;

   component Normalizer_Z_28_28_28_Freq500_uid8 is
      port ( clk, ce_6, ce_7, ce_8 : in std_logic;
             X : in  std_logic_vector(27 downto 0);
             Count : out  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_Freq500_uid11 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9 : in std_logic;
             X : in  std_logic_vector(33 downto 0);
             Y : in  std_logic_vector(33 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX_c0 :  std_logic_vector(32 downto 0);
signal excExpFracY_c0 :  std_logic_vector(32 downto 0);
signal swap_c0 :  std_logic;
signal eXmeY_c0 :  std_logic_vector(7 downto 0);
signal eYmeX_c0 :  std_logic_vector(7 downto 0);
signal expDiff_c0, expDiff_c1 :  std_logic_vector(7 downto 0);
signal newX_c0 :  std_logic_vector(33 downto 0);
signal newY_c0, newY_c1 :  std_logic_vector(33 downto 0);
signal expX_c0, expX_c1 :  std_logic_vector(7 downto 0);
signal excX_c0 :  std_logic_vector(1 downto 0);
signal excY_c0, excY_c1 :  std_logic_vector(1 downto 0);
signal signX_c0, signX_c1 :  std_logic;
signal signY_c0, signY_c1 :  std_logic;
signal EffSub_c1, EffSub_c2, EffSub_c3, EffSub_c4, EffSub_c5, EffSub_c6, EffSub_c7, EffSub_c8, EffSub_c9, EffSub_c10 :  std_logic;
signal sXsYExnXY_c0, sXsYExnXY_c1 :  std_logic_vector(5 downto 0);
signal sdExnXY_c0 :  std_logic_vector(3 downto 0);
signal fracY_c1 :  std_logic_vector(23 downto 0);
signal excRt_c1, excRt_c2, excRt_c3, excRt_c4, excRt_c5, excRt_c6, excRt_c7, excRt_c8, excRt_c9, excRt_c10 :  std_logic_vector(1 downto 0);
signal signR_c1, signR_c2, signR_c3, signR_c4, signR_c5, signR_c6, signR_c7, signR_c8 :  std_logic;
signal shiftedOut_c1 :  std_logic;
signal shiftVal_c1 :  std_logic_vector(4 downto 0);
signal shiftedFracY_c2 :  std_logic_vector(25 downto 0);
signal sticky_c4, sticky_c5 :  std_logic;
signal fracYpad_c2 :  std_logic_vector(26 downto 0);
signal EffSubVector_c1, EffSubVector_c2 :  std_logic_vector(26 downto 0);
signal fracYpadXorOp_c2 :  std_logic_vector(26 downto 0);
signal fracXpad_c0 :  std_logic_vector(26 downto 0);
signal cInSigAdd_c5 :  std_logic;
signal fracAddResult_c5 :  std_logic_vector(26 downto 0);
signal fracSticky_c5 :  std_logic_vector(27 downto 0);
signal nZerosNew_c8, nZerosNew_c9 :  std_logic_vector(4 downto 0);
signal shiftedFrac_c8, shiftedFrac_c9 :  std_logic_vector(27 downto 0);
signal extendedExpInc_c1, extendedExpInc_c2, extendedExpInc_c3, extendedExpInc_c4, extendedExpInc_c5, extendedExpInc_c6, extendedExpInc_c7, extendedExpInc_c8, extendedExpInc_c9 :  std_logic_vector(8 downto 0);
signal updatedExp_c9 :  std_logic_vector(9 downto 0);
signal eqdiffsign_c8, eqdiffsign_c9, eqdiffsign_c10 :  std_logic;
signal expFrac_c9 :  std_logic_vector(33 downto 0);
signal stk_c8, stk_c9 :  std_logic;
signal rnd_c8, rnd_c9 :  std_logic;
signal lsb_c8, lsb_c9 :  std_logic;
signal needToRound_c9 :  std_logic;
signal RoundedExpFrac_c9 :  std_logic_vector(33 downto 0);
signal upExc_c9 :  std_logic_vector(1 downto 0);
signal fracR_c9, fracR_c10 :  std_logic_vector(22 downto 0);
signal expR_c9, expR_c10 :  std_logic_vector(7 downto 0);
signal exExpExc_c9, exExpExc_c10 :  std_logic_vector(3 downto 0);
signal excRt2_c10 :  std_logic_vector(1 downto 0);
signal excR_c10 :  std_logic_vector(1 downto 0);
signal signR2_c8, signR2_c9, signR2_c10 :  std_logic;
signal computedR_c10 :  std_logic_vector(33 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               expDiff_c1 <= expDiff_c0;
               newY_c1 <= newY_c0;
               expX_c1 <= expX_c0;
               excY_c1 <= excY_c0;
               signX_c1 <= signX_c0;
               signY_c1 <= signY_c0;
               sXsYExnXY_c1 <= sXsYExnXY_c0;
            end if;
            if ce_2 = '1' then
               EffSub_c2 <= EffSub_c1;
               excRt_c2 <= excRt_c1;
               signR_c2 <= signR_c1;
               EffSubVector_c2 <= EffSubVector_c1;
               extendedExpInc_c2 <= extendedExpInc_c1;
            end if;
            if ce_3 = '1' then
               EffSub_c3 <= EffSub_c2;
               excRt_c3 <= excRt_c2;
               signR_c3 <= signR_c2;
               extendedExpInc_c3 <= extendedExpInc_c2;
            end if;
            if ce_4 = '1' then
               EffSub_c4 <= EffSub_c3;
               excRt_c4 <= excRt_c3;
               signR_c4 <= signR_c3;
               extendedExpInc_c4 <= extendedExpInc_c3;
            end if;
            if ce_5 = '1' then
               EffSub_c5 <= EffSub_c4;
               excRt_c5 <= excRt_c4;
               signR_c5 <= signR_c4;
               sticky_c5 <= sticky_c4;
               extendedExpInc_c5 <= extendedExpInc_c4;
            end if;
            if ce_6 = '1' then
               EffSub_c6 <= EffSub_c5;
               excRt_c6 <= excRt_c5;
               signR_c6 <= signR_c5;
               extendedExpInc_c6 <= extendedExpInc_c5;
            end if;
            if ce_7 = '1' then
               EffSub_c7 <= EffSub_c6;
               excRt_c7 <= excRt_c6;
               signR_c7 <= signR_c6;
               extendedExpInc_c7 <= extendedExpInc_c6;
            end if;
            if ce_8 = '1' then
               EffSub_c8 <= EffSub_c7;
               excRt_c8 <= excRt_c7;
               signR_c8 <= signR_c7;
               extendedExpInc_c8 <= extendedExpInc_c7;
            end if;
            if ce_9 = '1' then
               EffSub_c9 <= EffSub_c8;
               excRt_c9 <= excRt_c8;
               nZerosNew_c9 <= nZerosNew_c8;
               shiftedFrac_c9 <= shiftedFrac_c8;
               extendedExpInc_c9 <= extendedExpInc_c8;
               eqdiffsign_c9 <= eqdiffsign_c8;
               stk_c9 <= stk_c8;
               rnd_c9 <= rnd_c8;
               lsb_c9 <= lsb_c8;
               signR2_c9 <= signR2_c8;
            end if;
            if ce_10 = '1' then
               EffSub_c10 <= EffSub_c9;
               excRt_c10 <= excRt_c9;
               eqdiffsign_c10 <= eqdiffsign_c9;
               fracR_c10 <= fracR_c9;
               expR_c10 <= expR_c9;
               exExpExc_c10 <= exExpExc_c9;
               signR2_c10 <= signR2_c9;
            end if;
         end if;
      end process;
   excExpFracX_c0 <= X(33 downto 32) & X(30 downto 0);
   excExpFracY_c0 <= Y(33 downto 32) & Y(30 downto 0);
   swap_c0 <= '1' when excExpFracX_c0 < excExpFracY_c0 else '0';
   -- exponent difference
   eXmeY_c0 <= (X(30 downto 23)) - (Y(30 downto 23));
   eYmeX_c0 <= (Y(30 downto 23)) - (X(30 downto 23));
   expDiff_c0 <= eXmeY_c0 when swap_c0 = '0' else eYmeX_c0;
   -- input swap so that |X|>|Y|
   newX_c0 <= X when swap_c0 = '0' else Y;
   newY_c0 <= Y when swap_c0 = '0' else X;
   -- now we decompose the inputs into their sign, exponent, fraction
   expX_c0<= newX_c0(30 downto 23);
   excX_c0<= newX_c0(33 downto 32);
   excY_c0<= newY_c0(33 downto 32);
   signX_c0<= newX_c0(31);
   signY_c0<= newY_c0(31);
   EffSub_c1 <= signX_c1 xor signY_c1;
   sXsYExnXY_c0 <= signX_c0 & signY_c0 & excX_c0 & excY_c0;
   sdExnXY_c0 <= excX_c0 & excY_c0;
   fracY_c1 <= "000000000000000000000000" when excY_c1="00" else ('1' & newY_c1(22 downto 0));
   -- Exception management logic
   with sXsYExnXY_c1  select  
   excRt_c1 <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR_c1<= '0' when (sXsYExnXY_c1="100000" or sXsYExnXY_c1="010000") else signX_c1;
   shiftedOut_c1 <= '1' when (expDiff_c1 > 25) else '0';
   shiftVal_c1 <= expDiff_c1(4 downto 0) when shiftedOut_c1='0' else CONV_STD_LOGIC_VECTOR(26,5);
   RightShifterComponent: RightShifterSticky24_by_max_26_Freq500_uid4
      port map ( clk  => clk,
                 ce_2 => ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 S => shiftVal_c1,
                 X => fracY_c1,
                 R => shiftedFracY_c2,
                 Sticky => sticky_c4);
   fracYpad_c2 <= "0" & shiftedFracY_c2;
   EffSubVector_c1 <= (26 downto 0 => EffSub_c1);
   fracYpadXorOp_c2 <= fracYpad_c2 xor EffSubVector_c2;
   fracXpad_c0 <= "01" & (newX_c0(22 downto 0)) & "00";
   cInSigAdd_c5 <= EffSub_c5 and not sticky_c5; -- if we subtract and the sticky was one, some of the negated sticky bits would have absorbed this carry 
   fracAdder: IntAdder_27_Freq500_uid6
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 Cin => cInSigAdd_c5,
                 X => fracXpad_c0,
                 Y => fracYpadXorOp_c2,
                 R => fracAddResult_c5);
   fracSticky_c5<= fracAddResult_c5 & sticky_c5; 
   LZCAndShifter: Normalizer_Z_28_28_28_Freq500_uid8
      port map ( clk  => clk,
                 ce_6 => ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 X => fracSticky_c5,
                 Count => nZerosNew_c8,
                 R => shiftedFrac_c8);
   extendedExpInc_c1<= ("0" & expX_c1) + '1';
   updatedExp_c9 <= ("0" &extendedExpInc_c9) - ("00000" & nZerosNew_c9);
   eqdiffsign_c8 <= '1' when nZerosNew_c8="11111" else '0';
   expFrac_c9<= updatedExp_c9 & shiftedFrac_c9(26 downto 3);
   stk_c8<= shiftedFrac_c8(2) or shiftedFrac_c8(1) or shiftedFrac_c8(0);
   rnd_c8<= shiftedFrac_c8(3);
   lsb_c8<= shiftedFrac_c8(4);
   needToRound_c9<= '1' when (rnd_c9='1' and stk_c9='1') or (rnd_c9='1' and stk_c9='0' and lsb_c9='1')
  else '0';
   roundingAdder: IntAdder_34_Freq500_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 Cin => needToRound_c9,
                 X => expFrac_c9,
                 Y => "0000000000000000000000000000000000",
                 R => RoundedExpFrac_c9);
   -- possible update to exception bits
   upExc_c9 <= RoundedExpFrac_c9(33 downto 32);
   fracR_c9 <= RoundedExpFrac_c9(23 downto 1);
   expR_c9 <= RoundedExpFrac_c9(31 downto 24);
   exExpExc_c9 <= upExc_c9 & excRt_c9;
   with exExpExc_c10  select  
   excRt2_c10<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR_c10 <= "00" when (eqdiffsign_c10='1' and EffSub_c10='1'  and not(excRt_c10="11")) else excRt2_c10;
   signR2_c8 <= '0' when (eqdiffsign_c8='1' and EffSub_c8='1') else signR_c8;
   computedR_c10 <= excR_c10 & signR2_c10 & expR_c10 & fracR_c10;
   R <= computedR_c10;
end architecture;




--------------------------------------------------------------------------------
--                RightShifterSticky24_by_max_26_Freq300_uid4
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X S
-- Output signals: R Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifterSticky24_by_max_26_Freq300_uid4 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(25 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of RightShifterSticky24_by_max_26_Freq300_uid4 is
signal ps_c0, ps_c1, ps_c2 :  std_logic_vector(4 downto 0);
signal Xpadded_c0 :  std_logic_vector(25 downto 0);
signal level5_c0, level5_c1 :  std_logic_vector(25 downto 0);
signal stk4_c1 :  std_logic;
signal level4_c0, level4_c1 :  std_logic_vector(25 downto 0);
signal stk3_c1 :  std_logic;
signal level3_c1 :  std_logic_vector(25 downto 0);
signal stk2_c1, stk2_c2 :  std_logic;
signal level2_c1, level2_c2 :  std_logic_vector(25 downto 0);
signal stk1_c2 :  std_logic;
signal level1_c1, level1_c2 :  std_logic_vector(25 downto 0);
signal stk0_c2 :  std_logic;
signal level0_c1 :  std_logic_vector(25 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               ps_c1 <= ps_c0;
               level5_c1 <= level5_c0;
               level4_c1 <= level4_c0;
            end if;
            if ce_2 = '1' then
               ps_c2 <= ps_c1;
               stk2_c2 <= stk2_c1;
               level2_c2 <= level2_c1;
               level1_c2 <= level1_c1;
            end if;
         end if;
      end process;
   ps_c0<= S;
   Xpadded_c0 <= X&(1 downto 0 => '0');
   level5_c0<= Xpadded_c0;
   stk4_c1 <= '1' when (level5_c1(15 downto 0)/="0000000000000000" and ps_c1(4)='1')   else '0';
   level4_c0 <=  level5_c0 when  ps_c0(4)='0'    else (15 downto 0 => '0') & level5_c0(25 downto 16);
   stk3_c1 <= '1' when (level4_c1(7 downto 0)/="00000000" and ps_c1(3)='1') or stk4_c1 ='1'   else '0';
   level3_c1 <=  level4_c1 when  ps_c1(3)='0'    else (7 downto 0 => '0') & level4_c1(25 downto 8);
   stk2_c1 <= '1' when (level3_c1(3 downto 0)/="0000" and ps_c1(2)='1') or stk3_c1 ='1'   else '0';
   level2_c1 <=  level3_c1 when  ps_c1(2)='0'    else (3 downto 0 => '0') & level3_c1(25 downto 4);
   stk1_c2 <= '1' when (level2_c2(1 downto 0)/="00" and ps_c2(1)='1') or stk2_c2 ='1'   else '0';
   level1_c1 <=  level2_c1 when  ps_c1(1)='0'    else (1 downto 0 => '0') & level2_c1(25 downto 2);
   stk0_c2 <= '1' when (level1_c2(0 downto 0)/="0" and ps_c2(0)='1') or stk1_c2 ='1'   else '0';
   level0_c1 <=  level1_c1 when  ps_c1(0)='0'    else (0 downto 0 => '0') & level1_c1(25 downto 1);
   R <= level0_c1;
   Sticky <= stk0_c2;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_27_Freq300_uid6
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_Freq300_uid6 is
    port (clk, ce_1, ce_2, ce_3 : in std_logic;
          X : in  std_logic_vector(26 downto 0);
          Y : in  std_logic_vector(26 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_Freq300_uid6 is
signal Cin_1_c2, Cin_1_c3 :  std_logic;
signal X_1_c0, X_1_c1, X_1_c2, X_1_c3 :  std_logic_vector(27 downto 0);
signal Y_1_c1, Y_1_c2, Y_1_c3 :  std_logic_vector(27 downto 0);
signal S_1_c3 :  std_logic_vector(27 downto 0);
signal R_1_c3 :  std_logic_vector(26 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               X_1_c1 <= X_1_c0;
            end if;
            if ce_2 = '1' then
               X_1_c2 <= X_1_c1;
               Y_1_c2 <= Y_1_c1;
            end if;
            if ce_3 = '1' then
               Cin_1_c3 <= Cin_1_c2;
               X_1_c3 <= X_1_c2;
               Y_1_c3 <= Y_1_c2;
            end if;
         end if;
      end process;
   Cin_1_c2 <= Cin;
   X_1_c0 <= '0' & X(26 downto 0);
   Y_1_c1 <= '0' & Y(26 downto 0);
   S_1_c3 <= X_1_c3 + Y_1_c3 + Cin_1_c3;
   R_1_c3 <= S_1_c3(26 downto 0);
   R <= R_1_c3 ;
end architecture;

--------------------------------------------------------------------------------
--                     Normalizer_Z_28_28_28_Freq300_uid8
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_28_28_28_Freq300_uid8 is
    port (clk, ce_4, ce_5 : in std_logic;
          X : in  std_logic_vector(27 downto 0);
          Count : out  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of Normalizer_Z_28_28_28_Freq300_uid8 is
signal level5_c3 :  std_logic_vector(27 downto 0);
signal count4_c3, count4_c4 :  std_logic;
signal level4_c3, level4_c4 :  std_logic_vector(27 downto 0);
signal count3_c3, count3_c4 :  std_logic;
signal level3_c4 :  std_logic_vector(27 downto 0);
signal count2_c4 :  std_logic;
signal level2_c4 :  std_logic_vector(27 downto 0);
signal count1_c4 :  std_logic;
signal level1_c4, level1_c5 :  std_logic_vector(27 downto 0);
signal count0_c4, count0_c5 :  std_logic;
signal level0_c5 :  std_logic_vector(27 downto 0);
signal sCount_c4 :  std_logic_vector(4 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_4 = '1' then
               count4_c4 <= count4_c3;
               level4_c4 <= level4_c3;
               count3_c4 <= count3_c3;
            end if;
            if ce_5 = '1' then
               level1_c5 <= level1_c4;
               count0_c5 <= count0_c4;
            end if;
         end if;
      end process;
   level5_c3 <= X ;
   count4_c3<= '1' when level5_c3(27 downto 12) = (27 downto 12=>'0') else '0';
   level4_c3<= level5_c3(27 downto 0) when count4_c3='0' else level5_c3(11 downto 0) & (15 downto 0 => '0');

   count3_c3<= '1' when level4_c3(27 downto 20) = (27 downto 20=>'0') else '0';
   level3_c4<= level4_c4(27 downto 0) when count3_c4='0' else level4_c4(19 downto 0) & (7 downto 0 => '0');

   count2_c4<= '1' when level3_c4(27 downto 24) = (27 downto 24=>'0') else '0';
   level2_c4<= level3_c4(27 downto 0) when count2_c4='0' else level3_c4(23 downto 0) & (3 downto 0 => '0');

   count1_c4<= '1' when level2_c4(27 downto 26) = (27 downto 26=>'0') else '0';
   level1_c4<= level2_c4(27 downto 0) when count1_c4='0' else level2_c4(25 downto 0) & (1 downto 0 => '0');

   count0_c4<= '1' when level1_c4(27 downto 27) = (27 downto 27=>'0') else '0';
   level0_c5<= level1_c5(27 downto 0) when count0_c5='0' else level1_c5(26 downto 0) & (0 downto 0 => '0');

   R <= level0_c5;
   sCount_c4 <= count4_c4 & count3_c4 & count2_c4 & count1_c4 & count0_c4;
   Count <= sCount_c4;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_Freq300_uid11
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_Freq300_uid11 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5 : in std_logic;
          X : in  std_logic_vector(33 downto 0);
          Y : in  std_logic_vector(33 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_Freq300_uid11 is
signal Rtmp_c5 :  std_logic_vector(33 downto 0);
signal Y_c1, Y_c2, Y_c3, Y_c4, Y_c5 :  std_logic_vector(33 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               Y_c2 <= Y_c1;
            end if;
            if ce_3 = '1' then
               Y_c3 <= Y_c2;
            end if;
            if ce_4 = '1' then
               Y_c4 <= Y_c3;
            end if;
            if ce_5 = '1' then
               Y_c5 <= Y_c4;
            end if;
         end if;
      end process;
   Rtmp_c5 <= X + Y_c5 + Cin;
   R <= Rtmp_c5;
end architecture;

--------------------------------------------------------------------------------
--                             FloatingPointAdder
--                         (FPAdd_8_23_Freq300_uid2)
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2010-2017)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointAdder_32_3_649333 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointAdder_32_3_649333 is
   component RightShifterSticky24_by_max_26_Freq300_uid4 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(25 downto 0);
             Sticky : out  std_logic   );
   end component;

   component IntAdder_27_Freq300_uid6 is
      port ( clk, ce_1, ce_2, ce_3 : in std_logic;
             X : in  std_logic_vector(26 downto 0);
             Y : in  std_logic_vector(26 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(26 downto 0)   );
   end component;

   component Normalizer_Z_28_28_28_Freq300_uid8 is
      port ( clk, ce_4, ce_5 : in std_logic;
             X : in  std_logic_vector(27 downto 0);
             Count : out  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_Freq300_uid11 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5 : in std_logic;
             X : in  std_logic_vector(33 downto 0);
             Y : in  std_logic_vector(33 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX_c0 :  std_logic_vector(32 downto 0);
signal excExpFracY_c0 :  std_logic_vector(32 downto 0);
signal swap_c0 :  std_logic;
signal eXmeY_c0 :  std_logic_vector(7 downto 0);
signal eYmeX_c0 :  std_logic_vector(7 downto 0);
signal expDiff_c0 :  std_logic_vector(7 downto 0);
signal newX_c0 :  std_logic_vector(33 downto 0);
signal newY_c0 :  std_logic_vector(33 downto 0);
signal expX_c0 :  std_logic_vector(7 downto 0);
signal excX_c0 :  std_logic_vector(1 downto 0);
signal excY_c0 :  std_logic_vector(1 downto 0);
signal signX_c0 :  std_logic;
signal signY_c0 :  std_logic;
signal EffSub_c0, EffSub_c1, EffSub_c2, EffSub_c3, EffSub_c4, EffSub_c5, EffSub_c6 :  std_logic;
signal sXsYExnXY_c0 :  std_logic_vector(5 downto 0);
signal sdExnXY_c0 :  std_logic_vector(3 downto 0);
signal fracY_c0 :  std_logic_vector(23 downto 0);
signal excRt_c0, excRt_c1, excRt_c2, excRt_c3, excRt_c4, excRt_c5, excRt_c6 :  std_logic_vector(1 downto 0);
signal signR_c0, signR_c1, signR_c2, signR_c3, signR_c4, signR_c5 :  std_logic;
signal shiftedOut_c0 :  std_logic;
signal shiftVal_c0 :  std_logic_vector(4 downto 0);
signal shiftedFracY_c1 :  std_logic_vector(25 downto 0);
signal sticky_c2, sticky_c3 :  std_logic;
signal fracYpad_c1 :  std_logic_vector(26 downto 0);
signal EffSubVector_c0, EffSubVector_c1 :  std_logic_vector(26 downto 0);
signal fracYpadXorOp_c1 :  std_logic_vector(26 downto 0);
signal fracXpad_c0 :  std_logic_vector(26 downto 0);
signal cInSigAdd_c2 :  std_logic;
signal fracAddResult_c3 :  std_logic_vector(26 downto 0);
signal fracSticky_c3 :  std_logic_vector(27 downto 0);
signal nZerosNew_c4, nZerosNew_c5 :  std_logic_vector(4 downto 0);
signal shiftedFrac_c5 :  std_logic_vector(27 downto 0);
signal extendedExpInc_c0, extendedExpInc_c1, extendedExpInc_c2, extendedExpInc_c3, extendedExpInc_c4, extendedExpInc_c5 :  std_logic_vector(8 downto 0);
signal updatedExp_c5 :  std_logic_vector(9 downto 0);
signal eqdiffsign_c4, eqdiffsign_c5, eqdiffsign_c6 :  std_logic;
signal expFrac_c5 :  std_logic_vector(33 downto 0);
signal stk_c5 :  std_logic;
signal rnd_c5 :  std_logic;
signal lsb_c5 :  std_logic;
signal needToRound_c5 :  std_logic;
signal RoundedExpFrac_c5 :  std_logic_vector(33 downto 0);
signal upExc_c5 :  std_logic_vector(1 downto 0);
signal fracR_c5, fracR_c6 :  std_logic_vector(22 downto 0);
signal expR_c5, expR_c6 :  std_logic_vector(7 downto 0);
signal exExpExc_c5 :  std_logic_vector(3 downto 0);
signal excRt2_c5, excRt2_c6 :  std_logic_vector(1 downto 0);
signal excR_c6 :  std_logic_vector(1 downto 0);
signal signR2_c5, signR2_c6 :  std_logic;
signal computedR_c6 :  std_logic_vector(33 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               EffSub_c1 <= EffSub_c0;
               excRt_c1 <= excRt_c0;
               signR_c1 <= signR_c0;
               EffSubVector_c1 <= EffSubVector_c0;
               extendedExpInc_c1 <= extendedExpInc_c0;
            end if;
            if ce_2 = '1' then
               EffSub_c2 <= EffSub_c1;
               excRt_c2 <= excRt_c1;
               signR_c2 <= signR_c1;
               extendedExpInc_c2 <= extendedExpInc_c1;
            end if;
            if ce_3 = '1' then
               EffSub_c3 <= EffSub_c2;
               excRt_c3 <= excRt_c2;
               signR_c3 <= signR_c2;
               sticky_c3 <= sticky_c2;
               extendedExpInc_c3 <= extendedExpInc_c2;
            end if;
            if ce_4 = '1' then
               EffSub_c4 <= EffSub_c3;
               excRt_c4 <= excRt_c3;
               signR_c4 <= signR_c3;
               extendedExpInc_c4 <= extendedExpInc_c3;
            end if;
            if ce_5 = '1' then
               EffSub_c5 <= EffSub_c4;
               excRt_c5 <= excRt_c4;
               signR_c5 <= signR_c4;
               nZerosNew_c5 <= nZerosNew_c4;
               extendedExpInc_c5 <= extendedExpInc_c4;
               eqdiffsign_c5 <= eqdiffsign_c4;
            end if;
            if ce_6 = '1' then
               EffSub_c6 <= EffSub_c5;
               excRt_c6 <= excRt_c5;
               eqdiffsign_c6 <= eqdiffsign_c5;
               fracR_c6 <= fracR_c5;
               expR_c6 <= expR_c5;
               excRt2_c6 <= excRt2_c5;
               signR2_c6 <= signR2_c5;
            end if;
         end if;
      end process;
   excExpFracX_c0 <= X(33 downto 32) & X(30 downto 0);
   excExpFracY_c0 <= Y(33 downto 32) & Y(30 downto 0);
   swap_c0 <= '1' when excExpFracX_c0 < excExpFracY_c0 else '0';
   -- exponent difference
   eXmeY_c0 <= (X(30 downto 23)) - (Y(30 downto 23));
   eYmeX_c0 <= (Y(30 downto 23)) - (X(30 downto 23));
   expDiff_c0 <= eXmeY_c0 when swap_c0 = '0' else eYmeX_c0;
   -- input swap so that |X|>|Y|
   newX_c0 <= X when swap_c0 = '0' else Y;
   newY_c0 <= Y when swap_c0 = '0' else X;
   -- now we decompose the inputs into their sign, exponent, fraction
   expX_c0<= newX_c0(30 downto 23);
   excX_c0<= newX_c0(33 downto 32);
   excY_c0<= newY_c0(33 downto 32);
   signX_c0<= newX_c0(31);
   signY_c0<= newY_c0(31);
   EffSub_c0 <= signX_c0 xor signY_c0;
   sXsYExnXY_c0 <= signX_c0 & signY_c0 & excX_c0 & excY_c0;
   sdExnXY_c0 <= excX_c0 & excY_c0;
   fracY_c0 <= "000000000000000000000000" when excY_c0="00" else ('1' & newY_c0(22 downto 0));
   -- Exception management logic
   with sXsYExnXY_c0  select  
   excRt_c0 <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR_c0<= '0' when (sXsYExnXY_c0="100000" or sXsYExnXY_c0="010000") else signX_c0;
   shiftedOut_c0 <= '1' when (expDiff_c0 > 25) else '0';
   shiftVal_c0 <= expDiff_c0(4 downto 0) when shiftedOut_c0='0' else CONV_STD_LOGIC_VECTOR(26,5);
   RightShifterComponent: RightShifterSticky24_by_max_26_Freq300_uid4
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 S => shiftVal_c0,
                 X => fracY_c0,
                 R => shiftedFracY_c1,
                 Sticky => sticky_c2);
   fracYpad_c1 <= "0" & shiftedFracY_c1;
   EffSubVector_c0 <= (26 downto 0 => EffSub_c0);
   fracYpadXorOp_c1 <= fracYpad_c1 xor EffSubVector_c1;
   fracXpad_c0 <= "01" & (newX_c0(22 downto 0)) & "00";
   cInSigAdd_c2 <= EffSub_c2 and not sticky_c2; -- if we subtract and the sticky was one, some of the negated sticky bits would have absorbed this carry 
   fracAdder: IntAdder_27_Freq300_uid6
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 Cin => cInSigAdd_c2,
                 X => fracXpad_c0,
                 Y => fracYpadXorOp_c1,
                 R => fracAddResult_c3);
   fracSticky_c3<= fracAddResult_c3 & sticky_c3; 
   LZCAndShifter: Normalizer_Z_28_28_28_Freq300_uid8
      port map ( clk  => clk,
                 ce_4 => ce_4,
                 ce_5=> ce_5,
                 X => fracSticky_c3,
                 Count => nZerosNew_c4,
                 R => shiftedFrac_c5);
   extendedExpInc_c0<= ("0" & expX_c0) + '1';
   updatedExp_c5 <= ("0" &extendedExpInc_c5) - ("00000" & nZerosNew_c5);
   eqdiffsign_c4 <= '1' when nZerosNew_c4="11111" else '0';
   expFrac_c5<= updatedExp_c5 & shiftedFrac_c5(26 downto 3);
   stk_c5<= shiftedFrac_c5(2) or shiftedFrac_c5(1) or shiftedFrac_c5(0);
   rnd_c5<= shiftedFrac_c5(3);
   lsb_c5<= shiftedFrac_c5(4);
   needToRound_c5<= '1' when (rnd_c5='1' and stk_c5='1') or (rnd_c5='1' and stk_c5='0' and lsb_c5='1')
  else '0';
   roundingAdder: IntAdder_34_Freq300_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 Cin => needToRound_c5,
                 X => expFrac_c5,
                 Y => "0000000000000000000000000000000000",
                 R => RoundedExpFrac_c5);
   -- possible update to exception bits
   upExc_c5 <= RoundedExpFrac_c5(33 downto 32);
   fracR_c5 <= RoundedExpFrac_c5(23 downto 1);
   expR_c5 <= RoundedExpFrac_c5(31 downto 24);
   exExpExc_c5 <= upExc_c5 & excRt_c5;
   with exExpExc_c5  select  
   excRt2_c5<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR_c6 <= "00" when (eqdiffsign_c6='1' and EffSub_c6='1'  and not(excRt_c6="11")) else excRt2_c6;
   signR2_c5 <= '0' when (eqdiffsign_c5='1' and EffSub_c5='1') else signR_c5;
   computedR_c6 <= excR_c6 & signR2_c6 & expR_c6 & fracR_c6;
   R <= computedR_c6;
end architecture;




--------------------------------------------------------------------------------
--                RightShifterSticky24_by_max_26_Freq100_uid4
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X S
-- Output signals: R Sticky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifterSticky24_by_max_26_Freq100_uid4 is
    port (clk : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(25 downto 0);
          Sticky : out  std_logic   );
end entity;

architecture arch of RightShifterSticky24_by_max_26_Freq100_uid4 is
signal ps_c0 :  std_logic_vector(4 downto 0);
signal Xpadded_c0 :  std_logic_vector(25 downto 0);
signal level5_c0 :  std_logic_vector(25 downto 0);
signal stk4_c0 :  std_logic;
signal level4_c0 :  std_logic_vector(25 downto 0);
signal stk3_c0 :  std_logic;
signal level3_c0 :  std_logic_vector(25 downto 0);
signal stk2_c0 :  std_logic;
signal level2_c0 :  std_logic_vector(25 downto 0);
signal stk1_c0 :  std_logic;
signal level1_c0 :  std_logic_vector(25 downto 0);
signal stk0_c0 :  std_logic;
signal level0_c0 :  std_logic_vector(25 downto 0);
begin
   ps_c0<= S;
   Xpadded_c0 <= X&(1 downto 0 => '0');
   level5_c0<= Xpadded_c0;
   stk4_c0 <= '1' when (level5_c0(15 downto 0)/="0000000000000000" and ps_c0(4)='1')   else '0';
   level4_c0 <=  level5_c0 when  ps_c0(4)='0'    else (15 downto 0 => '0') & level5_c0(25 downto 16);
   stk3_c0 <= '1' when (level4_c0(7 downto 0)/="00000000" and ps_c0(3)='1') or stk4_c0 ='1'   else '0';
   level3_c0 <=  level4_c0 when  ps_c0(3)='0'    else (7 downto 0 => '0') & level4_c0(25 downto 8);
   stk2_c0 <= '1' when (level3_c0(3 downto 0)/="0000" and ps_c0(2)='1') or stk3_c0 ='1'   else '0';
   level2_c0 <=  level3_c0 when  ps_c0(2)='0'    else (3 downto 0 => '0') & level3_c0(25 downto 4);
   stk1_c0 <= '1' when (level2_c0(1 downto 0)/="00" and ps_c0(1)='1') or stk2_c0 ='1'   else '0';
   level1_c0 <=  level2_c0 when  ps_c0(1)='0'    else (1 downto 0 => '0') & level2_c0(25 downto 2);
   stk0_c0 <= '1' when (level1_c0(0 downto 0)/="0" and ps_c0(0)='1') or stk1_c0 ='1'   else '0';
   level0_c0 <=  level1_c0 when  ps_c0(0)='0'    else (0 downto 0 => '0') & level1_c0(25 downto 1);
   R <= level0_c0;
   Sticky <= stk0_c0;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_27_Freq100_uid6
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_27_Freq100_uid6 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(26 downto 0);
          Y : in  std_logic_vector(26 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(26 downto 0)   );
end entity;

architecture arch of IntAdder_27_Freq100_uid6 is
signal Cin_1_c0, Cin_1_c1 :  std_logic;
signal X_1_c0, X_1_c1 :  std_logic_vector(27 downto 0);
signal Y_1_c0, Y_1_c1 :  std_logic_vector(27 downto 0);
signal S_1_c1 :  std_logic_vector(27 downto 0);
signal R_1_c1 :  std_logic_vector(26 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_1_c1 <= Cin_1_c0;
               X_1_c1 <= X_1_c0;
               Y_1_c1 <= Y_1_c0;
            end if;
         end if;
      end process;
   Cin_1_c0 <= Cin;
   X_1_c0 <= '0' & X(26 downto 0);
   Y_1_c0 <= '0' & Y(26 downto 0);
   S_1_c1 <= X_1_c1 + Y_1_c1 + Cin_1_c1;
   R_1_c1 <= S_1_c1(26 downto 0);
   R <= R_1_c1 ;
end architecture;

--------------------------------------------------------------------------------
--                     Normalizer_Z_28_28_28_Freq100_uid8
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_Z_28_28_28_Freq100_uid8 is
    port (clk : in std_logic;
          X : in  std_logic_vector(27 downto 0);
          Count : out  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(27 downto 0)   );
end entity;

architecture arch of Normalizer_Z_28_28_28_Freq100_uid8 is
signal level5_c1 :  std_logic_vector(27 downto 0);
signal count4_c1 :  std_logic;
signal level4_c1 :  std_logic_vector(27 downto 0);
signal count3_c1 :  std_logic;
signal level3_c1 :  std_logic_vector(27 downto 0);
signal count2_c1 :  std_logic;
signal level2_c1 :  std_logic_vector(27 downto 0);
signal count1_c1 :  std_logic;
signal level1_c1 :  std_logic_vector(27 downto 0);
signal count0_c1 :  std_logic;
signal level0_c1 :  std_logic_vector(27 downto 0);
signal sCount_c1 :  std_logic_vector(4 downto 0);
begin
   level5_c1 <= X ;
   count4_c1<= '1' when level5_c1(27 downto 12) = (27 downto 12=>'0') else '0';
   level4_c1<= level5_c1(27 downto 0) when count4_c1='0' else level5_c1(11 downto 0) & (15 downto 0 => '0');

   count3_c1<= '1' when level4_c1(27 downto 20) = (27 downto 20=>'0') else '0';
   level3_c1<= level4_c1(27 downto 0) when count3_c1='0' else level4_c1(19 downto 0) & (7 downto 0 => '0');

   count2_c1<= '1' when level3_c1(27 downto 24) = (27 downto 24=>'0') else '0';
   level2_c1<= level3_c1(27 downto 0) when count2_c1='0' else level3_c1(23 downto 0) & (3 downto 0 => '0');

   count1_c1<= '1' when level2_c1(27 downto 26) = (27 downto 26=>'0') else '0';
   level1_c1<= level2_c1(27 downto 0) when count1_c1='0' else level2_c1(25 downto 0) & (1 downto 0 => '0');

   count0_c1<= '1' when level1_c1(27 downto 27) = (27 downto 27=>'0') else '0';
   level0_c1<= level1_c1(27 downto 0) when count0_c1='0' else level1_c1(26 downto 0) & (0 downto 0 => '0');

   R <= level0_c1;
   sCount_c1 <= count4_c1 & count3_c1 & count2_c1 & count1_c1 & count0_c1;
   Count <= sCount_c1;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_34_Freq100_uid11
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_34_Freq100_uid11 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(33 downto 0);
          Y : in  std_logic_vector(33 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(33 downto 0)   );
end entity;

architecture arch of IntAdder_34_Freq100_uid11 is
signal Rtmp_c1 :  std_logic_vector(33 downto 0);
signal Y_c1 :  std_logic_vector(33 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
         end if;
      end process;
   Rtmp_c1 <= X + Y_c1 + Cin;
   R <= Rtmp_c1;
end architecture;

--------------------------------------------------------------------------------
--                             FloatingPointAdder
--                         (FPAdd_8_23_Freq100_uid2)
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2010-2017)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointAdder_32_9_068000 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointAdder_32_9_068000 is
   component RightShifterSticky24_by_max_26_Freq100_uid4 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(25 downto 0);
             Sticky : out  std_logic   );
   end component;

   component IntAdder_27_Freq100_uid6 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(26 downto 0);
             Y : in  std_logic_vector(26 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(26 downto 0)   );
   end component;

   component Normalizer_Z_28_28_28_Freq100_uid8 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(27 downto 0);
             Count : out  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(27 downto 0)   );
   end component;

   component IntAdder_34_Freq100_uid11 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(33 downto 0);
             Y : in  std_logic_vector(33 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(33 downto 0)   );
   end component;

signal excExpFracX_c0 :  std_logic_vector(32 downto 0);
signal excExpFracY_c0 :  std_logic_vector(32 downto 0);
signal swap_c0 :  std_logic;
signal eXmeY_c0 :  std_logic_vector(7 downto 0);
signal eYmeX_c0 :  std_logic_vector(7 downto 0);
signal expDiff_c0 :  std_logic_vector(7 downto 0);
signal newX_c0 :  std_logic_vector(33 downto 0);
signal newY_c0 :  std_logic_vector(33 downto 0);
signal expX_c0 :  std_logic_vector(7 downto 0);
signal excX_c0 :  std_logic_vector(1 downto 0);
signal excY_c0 :  std_logic_vector(1 downto 0);
signal signX_c0 :  std_logic;
signal signY_c0 :  std_logic;
signal EffSub_c0, EffSub_c1 :  std_logic;
signal sXsYExnXY_c0 :  std_logic_vector(5 downto 0);
signal sdExnXY_c0 :  std_logic_vector(3 downto 0);
signal fracY_c0 :  std_logic_vector(23 downto 0);
signal excRt_c0, excRt_c1 :  std_logic_vector(1 downto 0);
signal signR_c0, signR_c1 :  std_logic;
signal shiftedOut_c0 :  std_logic;
signal shiftVal_c0 :  std_logic_vector(4 downto 0);
signal shiftedFracY_c0 :  std_logic_vector(25 downto 0);
signal sticky_c0, sticky_c1 :  std_logic;
signal fracYpad_c0 :  std_logic_vector(26 downto 0);
signal EffSubVector_c0 :  std_logic_vector(26 downto 0);
signal fracYpadXorOp_c0 :  std_logic_vector(26 downto 0);
signal fracXpad_c0 :  std_logic_vector(26 downto 0);
signal cInSigAdd_c0 :  std_logic;
signal fracAddResult_c1 :  std_logic_vector(26 downto 0);
signal fracSticky_c1 :  std_logic_vector(27 downto 0);
signal nZerosNew_c1 :  std_logic_vector(4 downto 0);
signal shiftedFrac_c1 :  std_logic_vector(27 downto 0);
signal extendedExpInc_c0, extendedExpInc_c1 :  std_logic_vector(8 downto 0);
signal updatedExp_c1 :  std_logic_vector(9 downto 0);
signal eqdiffsign_c1 :  std_logic;
signal expFrac_c1 :  std_logic_vector(33 downto 0);
signal stk_c1 :  std_logic;
signal rnd_c1 :  std_logic;
signal lsb_c1 :  std_logic;
signal needToRound_c1 :  std_logic;
signal RoundedExpFrac_c1 :  std_logic_vector(33 downto 0);
signal upExc_c1 :  std_logic_vector(1 downto 0);
signal fracR_c1 :  std_logic_vector(22 downto 0);
signal expR_c1 :  std_logic_vector(7 downto 0);
signal exExpExc_c1 :  std_logic_vector(3 downto 0);
signal excRt2_c1 :  std_logic_vector(1 downto 0);
signal excR_c1 :  std_logic_vector(1 downto 0);
signal signR2_c1 :  std_logic;
signal computedR_c1 :  std_logic_vector(33 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               EffSub_c1 <= EffSub_c0;
               excRt_c1 <= excRt_c0;
               signR_c1 <= signR_c0;
               sticky_c1 <= sticky_c0;
               extendedExpInc_c1 <= extendedExpInc_c0;
            end if;
         end if;
      end process;
   excExpFracX_c0 <= X(33 downto 32) & X(30 downto 0);
   excExpFracY_c0 <= Y(33 downto 32) & Y(30 downto 0);
   swap_c0 <= '1' when excExpFracX_c0 < excExpFracY_c0 else '0';
   -- exponent difference
   eXmeY_c0 <= (X(30 downto 23)) - (Y(30 downto 23));
   eYmeX_c0 <= (Y(30 downto 23)) - (X(30 downto 23));
   expDiff_c0 <= eXmeY_c0 when swap_c0 = '0' else eYmeX_c0;
   -- input swap so that |X|>|Y|
   newX_c0 <= X when swap_c0 = '0' else Y;
   newY_c0 <= Y when swap_c0 = '0' else X;
   -- now we decompose the inputs into their sign, exponent, fraction
   expX_c0<= newX_c0(30 downto 23);
   excX_c0<= newX_c0(33 downto 32);
   excY_c0<= newY_c0(33 downto 32);
   signX_c0<= newX_c0(31);
   signY_c0<= newY_c0(31);
   EffSub_c0 <= signX_c0 xor signY_c0;
   sXsYExnXY_c0 <= signX_c0 & signY_c0 & excX_c0 & excY_c0;
   sdExnXY_c0 <= excX_c0 & excY_c0;
   fracY_c0 <= "000000000000000000000000" when excY_c0="00" else ('1' & newY_c0(22 downto 0));
   -- Exception management logic
   with sXsYExnXY_c0  select  
   excRt_c0 <= "00" when "000000"|"010000"|"100000"|"110000",
      "01" when "000101"|"010101"|"100101"|"110101"|"000100"|"010100"|"100100"|"110100"|"000001"|"010001"|"100001"|"110001",
      "10" when "111010"|"001010"|"001000"|"011000"|"101000"|"111000"|"000010"|"010010"|"100010"|"110010"|"001001"|"011001"|"101001"|"111001"|"000110"|"010110"|"100110"|"110110", 
      "11" when others;
   signR_c0<= '0' when (sXsYExnXY_c0="100000" or sXsYExnXY_c0="010000") else signX_c0;
   shiftedOut_c0 <= '1' when (expDiff_c0 > 25) else '0';
   shiftVal_c0 <= expDiff_c0(4 downto 0) when shiftedOut_c0='0' else CONV_STD_LOGIC_VECTOR(26,5);
   RightShifterComponent: RightShifterSticky24_by_max_26_Freq100_uid4
      port map ( clk  => clk,
                 S => shiftVal_c0,
                 X => fracY_c0,
                 R => shiftedFracY_c0,
                 Sticky => sticky_c0);
   fracYpad_c0 <= "0" & shiftedFracY_c0;
   EffSubVector_c0 <= (26 downto 0 => EffSub_c0);
   fracYpadXorOp_c0 <= fracYpad_c0 xor EffSubVector_c0;
   fracXpad_c0 <= "01" & (newX_c0(22 downto 0)) & "00";
   cInSigAdd_c0 <= EffSub_c0 and not sticky_c0; -- if we subtract and the sticky was one, some of the negated sticky bits would have absorbed this carry 
   fracAdder: IntAdder_27_Freq100_uid6
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 Cin => cInSigAdd_c0,
                 X => fracXpad_c0,
                 Y => fracYpadXorOp_c0,
                 R => fracAddResult_c1);
   fracSticky_c1<= fracAddResult_c1 & sticky_c1; 
   LZCAndShifter: Normalizer_Z_28_28_28_Freq100_uid8
      port map ( clk  => clk,
                 X => fracSticky_c1,
                 Count => nZerosNew_c1,
                 R => shiftedFrac_c1);
   extendedExpInc_c0<= ("0" & expX_c0) + '1';
   updatedExp_c1 <= ("0" &extendedExpInc_c1) - ("00000" & nZerosNew_c1);
   eqdiffsign_c1 <= '1' when nZerosNew_c1="11111" else '0';
   expFrac_c1<= updatedExp_c1 & shiftedFrac_c1(26 downto 3);
   stk_c1<= shiftedFrac_c1(2) or shiftedFrac_c1(1) or shiftedFrac_c1(0);
   rnd_c1<= shiftedFrac_c1(3);
   lsb_c1<= shiftedFrac_c1(4);
   needToRound_c1<= '1' when (rnd_c1='1' and stk_c1='1') or (rnd_c1='1' and stk_c1='0' and lsb_c1='1')
  else '0';
   roundingAdder: IntAdder_34_Freq100_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 Cin => needToRound_c1,
                 X => expFrac_c1,
                 Y => "0000000000000000000000000000000000",
                 R => RoundedExpFrac_c1);
   -- possible update to exception bits
   upExc_c1 <= RoundedExpFrac_c1(33 downto 32);
   fracR_c1 <= RoundedExpFrac_c1(23 downto 1);
   expR_c1 <= RoundedExpFrac_c1(31 downto 24);
   exExpExc_c1 <= upExc_c1 & excRt_c1;
   with exExpExc_c1  select  
   excRt2_c1<= "00" when "0000"|"0100"|"1000"|"1100"|"1001"|"1101",
      "01" when "0001",
      "10" when "0010"|"0110"|"1010"|"1110"|"0101",
      "11" when others;
   excR_c1 <= "00" when (eqdiffsign_c1='1' and EffSub_c1='1'  and not(excRt_c1="11")) else excRt2_c1;
   signR2_c1 <= '0' when (eqdiffsign_c1='1' and EffSub_c1='1') else signR_c1;
   computedR_c1 <= excR_c1 & signR2_c1 & expR_c1 & fracR_c1;
   R <= computedR_c1;
end architecture;




--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid15
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid15 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid15 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid20
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid20 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid20 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid27
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid27 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid27 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid32
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid32 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid32 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid39
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid39 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid39 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid44
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid44 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid44 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid51
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid51 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid51 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid56
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid56 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid56 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid63
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid63 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid63 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid68
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid68 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid68 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid75
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid75 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid75 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid80
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid80 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid80 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid87
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid87 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid87 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid92
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid92 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid92 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid99
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid99 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid99 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid104
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid104 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid104 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid111
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid111 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid111 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid116
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid116 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid116 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid123
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid128
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid128 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid128 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid135
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid135 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid135 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid140
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid140 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid140 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid147
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid147 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid147 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid152
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid152 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid152 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq800_uid156
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq800_uid156 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq800_uid156 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq800_uid160
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq800_uid160 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq800_uid160 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq800_uid164
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq800_uid164 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq800_uid164 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq800_uid170
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq800_uid170 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq800_uid170 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid9
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid9 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid9 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq800_uid11
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid11 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid11 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid13
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid13 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid13 is
   component MultTable_Freq800_uid15 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy16_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid15
      port map ( X => Xtable_c0,
                 Y => Y1_copy16_c0);
   Y1_c0 <= Y1_copy16_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid18
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid18 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid18 is
   component MultTable_Freq800_uid20 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy21_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid20
      port map ( X => Xtable_c0,
                 Y => Y1_copy21_c0);
   Y1_c0 <= Y1_copy21_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq800_uid23
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid23 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid23 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid25
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid25 is
   component MultTable_Freq800_uid27 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy28_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid27
      port map ( X => Xtable_c0,
                 Y => Y1_copy28_c0);
   Y1_c0 <= Y1_copy28_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid30
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid30 is
   component MultTable_Freq800_uid32 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy33_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid32
      port map ( X => Xtable_c0,
                 Y => Y1_copy33_c0);
   Y1_c0 <= Y1_copy33_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq800_uid35
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid35 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid35 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid37
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid37 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid37 is
   component MultTable_Freq800_uid39 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy40_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid39
      port map ( X => Xtable_c0,
                 Y => Y1_copy40_c0);
   Y1_c0 <= Y1_copy40_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid42
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid42 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid42 is
   component MultTable_Freq800_uid44 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy45_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid44
      port map ( X => Xtable_c0,
                 Y => Y1_copy45_c0);
   Y1_c0 <= Y1_copy45_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq800_uid47
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid47 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid47 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid49
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid49 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid49 is
   component MultTable_Freq800_uid51 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy52_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid51
      port map ( X => Xtable_c0,
                 Y => Y1_copy52_c0);
   Y1_c0 <= Y1_copy52_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid54
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid54 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid54 is
   component MultTable_Freq800_uid56 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy57_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid56
      port map ( X => Xtable_c0,
                 Y => Y1_copy57_c0);
   Y1_c0 <= Y1_copy57_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq800_uid59
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid59 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid59 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid61
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid61 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid61 is
   component MultTable_Freq800_uid63 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy64_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid63
      port map ( X => Xtable_c0,
                 Y => Y1_copy64_c0);
   Y1_c0 <= Y1_copy64_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid66
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid66 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid66 is
   component MultTable_Freq800_uid68 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy69_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid68
      port map ( X => Xtable_c0,
                 Y => Y1_copy69_c0);
   Y1_c0 <= Y1_copy69_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq800_uid71
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid71 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid73
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid73 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid73 is
   component MultTable_Freq800_uid75 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy76_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid75
      port map ( X => Xtable_c0,
                 Y => Y1_copy76_c0);
   Y1_c0 <= Y1_copy76_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid78
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid78 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid78 is
   component MultTable_Freq800_uid80 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy81_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid80
      port map ( X => Xtable_c0,
                 Y => Y1_copy81_c0);
   Y1_c0 <= Y1_copy81_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq800_uid83
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid83 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid83 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid85
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid85 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid85 is
   component MultTable_Freq800_uid87 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy88_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid87
      port map ( X => Xtable_c0,
                 Y => Y1_copy88_c0);
   Y1_c0 <= Y1_copy88_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid90
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid90 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid90 is
   component MultTable_Freq800_uid92 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy93_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid92
      port map ( X => Xtable_c0,
                 Y => Y1_copy93_c0);
   Y1_c0 <= Y1_copy93_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq800_uid95
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid95 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid95 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq800_uid97
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid97 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid97 is
   component MultTable_Freq800_uid99 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy100_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid99
      port map ( X => Xtable_c0,
                 Y => Y1_copy100_c0);
   Y1_c0 <= Y1_copy100_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid102
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid102 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid102 is
   component MultTable_Freq800_uid104 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy105_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid104
      port map ( X => Xtable_c0,
                 Y => Y1_copy105_c0);
   Y1_c0 <= Y1_copy105_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq800_uid107
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid107 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid107 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid109
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid109 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid109 is
   component MultTable_Freq800_uid111 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy112_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid111
      port map ( X => Xtable_c0,
                 Y => Y1_copy112_c0);
   Y1_c0 <= Y1_copy112_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid114
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid114 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid114 is
   component MultTable_Freq800_uid116 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy117_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid116
      port map ( X => Xtable_c0,
                 Y => Y1_copy117_c0);
   Y1_c0 <= Y1_copy117_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq800_uid119
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid119 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid119 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid121
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid121 is
   component MultTable_Freq800_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy124_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid123
      port map ( X => Xtable_c0,
                 Y => Y1_copy124_c0);
   Y1_c0 <= Y1_copy124_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid126
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid126 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid126 is
   component MultTable_Freq800_uid128 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy129_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid128
      port map ( X => Xtable_c0,
                 Y => Y1_copy129_c0);
   Y1_c0 <= Y1_copy129_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq800_uid131
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid131 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid131 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid133
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid133 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid133 is
   component MultTable_Freq800_uid135 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy136_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid135
      port map ( X => Xtable_c0,
                 Y => Y1_copy136_c0);
   Y1_c0 <= Y1_copy136_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid138
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid138 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid138 is
   component MultTable_Freq800_uid140 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy141_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid140
      port map ( X => Xtable_c0,
                 Y => Y1_copy141_c0);
   Y1_c0 <= Y1_copy141_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq800_uid143
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq800_uid143 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq800_uid143 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid145
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid145 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid145 is
   component MultTable_Freq800_uid147 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy148_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid147
      port map ( X => Xtable_c0,
                 Y => Y1_copy148_c0);
   Y1_c0 <= Y1_copy148_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid150
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid150 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid150 is
   component MultTable_Freq800_uid152 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy153_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid152
      port map ( X => Xtable_c0,
                 Y => Y1_copy153_c0);
   Y1_c0 <= Y1_copy153_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_30_Freq800_uid352
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_30_Freq800_uid352 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13 : in std_logic;
          X : in  std_logic_vector(29 downto 0);
          Y : in  std_logic_vector(29 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of IntAdder_30_Freq800_uid352 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3, Cin_0_c4 :  std_logic;
signal X_0_c3, X_0_c4 :  std_logic_vector(3 downto 0);
signal Y_0_c3, Y_0_c4 :  std_logic_vector(3 downto 0);
signal S_0_c4 :  std_logic_vector(3 downto 0);
signal R_0_c4, R_0_c5, R_0_c6, R_0_c7, R_0_c8, R_0_c9, R_0_c10, R_0_c11, R_0_c12, R_0_c13 :  std_logic_vector(2 downto 0);
signal Cin_1_c4, Cin_1_c5 :  std_logic;
signal X_1_c3, X_1_c4, X_1_c5 :  std_logic_vector(3 downto 0);
signal Y_1_c3, Y_1_c4, Y_1_c5 :  std_logic_vector(3 downto 0);
signal S_1_c5 :  std_logic_vector(3 downto 0);
signal R_1_c5, R_1_c6, R_1_c7, R_1_c8, R_1_c9, R_1_c10, R_1_c11, R_1_c12, R_1_c13 :  std_logic_vector(2 downto 0);
signal Cin_2_c5, Cin_2_c6 :  std_logic;
signal X_2_c3, X_2_c4, X_2_c5, X_2_c6 :  std_logic_vector(3 downto 0);
signal Y_2_c3, Y_2_c4, Y_2_c5, Y_2_c6 :  std_logic_vector(3 downto 0);
signal S_2_c6 :  std_logic_vector(3 downto 0);
signal R_2_c6, R_2_c7, R_2_c8, R_2_c9, R_2_c10, R_2_c11, R_2_c12, R_2_c13 :  std_logic_vector(2 downto 0);
signal Cin_3_c6, Cin_3_c7 :  std_logic;
signal X_3_c3, X_3_c4, X_3_c5, X_3_c6, X_3_c7 :  std_logic_vector(3 downto 0);
signal Y_3_c3, Y_3_c4, Y_3_c5, Y_3_c6, Y_3_c7 :  std_logic_vector(3 downto 0);
signal S_3_c7 :  std_logic_vector(3 downto 0);
signal R_3_c7, R_3_c8, R_3_c9, R_3_c10, R_3_c11, R_3_c12, R_3_c13 :  std_logic_vector(2 downto 0);
signal Cin_4_c7, Cin_4_c8 :  std_logic;
signal X_4_c3, X_4_c4, X_4_c5, X_4_c6, X_4_c7, X_4_c8 :  std_logic_vector(3 downto 0);
signal Y_4_c3, Y_4_c4, Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8 :  std_logic_vector(3 downto 0);
signal S_4_c8 :  std_logic_vector(3 downto 0);
signal R_4_c8, R_4_c9, R_4_c10, R_4_c11, R_4_c12, R_4_c13 :  std_logic_vector(2 downto 0);
signal Cin_5_c8, Cin_5_c9 :  std_logic;
signal X_5_c3, X_5_c4, X_5_c5, X_5_c6, X_5_c7, X_5_c8, X_5_c9 :  std_logic_vector(3 downto 0);
signal Y_5_c3, Y_5_c4, Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9 :  std_logic_vector(3 downto 0);
signal S_5_c9 :  std_logic_vector(3 downto 0);
signal R_5_c9, R_5_c10, R_5_c11, R_5_c12, R_5_c13 :  std_logic_vector(2 downto 0);
signal Cin_6_c9, Cin_6_c10 :  std_logic;
signal X_6_c3, X_6_c4, X_6_c5, X_6_c6, X_6_c7, X_6_c8, X_6_c9, X_6_c10 :  std_logic_vector(3 downto 0);
signal Y_6_c3, Y_6_c4, Y_6_c5, Y_6_c6, Y_6_c7, Y_6_c8, Y_6_c9, Y_6_c10 :  std_logic_vector(3 downto 0);
signal S_6_c10 :  std_logic_vector(3 downto 0);
signal R_6_c10, R_6_c11, R_6_c12, R_6_c13 :  std_logic_vector(2 downto 0);
signal Cin_7_c10, Cin_7_c11 :  std_logic;
signal X_7_c3, X_7_c4, X_7_c5, X_7_c6, X_7_c7, X_7_c8, X_7_c9, X_7_c10, X_7_c11 :  std_logic_vector(3 downto 0);
signal Y_7_c3, Y_7_c4, Y_7_c5, Y_7_c6, Y_7_c7, Y_7_c8, Y_7_c9, Y_7_c10, Y_7_c11 :  std_logic_vector(3 downto 0);
signal S_7_c11 :  std_logic_vector(3 downto 0);
signal R_7_c11, R_7_c12, R_7_c13 :  std_logic_vector(2 downto 0);
signal Cin_8_c11, Cin_8_c12 :  std_logic;
signal X_8_c3, X_8_c4, X_8_c5, X_8_c6, X_8_c7, X_8_c8, X_8_c9, X_8_c10, X_8_c11, X_8_c12 :  std_logic_vector(3 downto 0);
signal Y_8_c3, Y_8_c4, Y_8_c5, Y_8_c6, Y_8_c7, Y_8_c8, Y_8_c9, Y_8_c10, Y_8_c11, Y_8_c12 :  std_logic_vector(3 downto 0);
signal S_8_c12 :  std_logic_vector(3 downto 0);
signal R_8_c12, R_8_c13 :  std_logic_vector(2 downto 0);
signal Cin_9_c12, Cin_9_c13 :  std_logic;
signal X_9_c3, X_9_c4, X_9_c5, X_9_c6, X_9_c7, X_9_c8, X_9_c9, X_9_c10, X_9_c11, X_9_c12, X_9_c13 :  std_logic_vector(3 downto 0);
signal Y_9_c3, Y_9_c4, Y_9_c5, Y_9_c6, Y_9_c7, Y_9_c8, Y_9_c9, Y_9_c10, Y_9_c11, Y_9_c12, Y_9_c13 :  std_logic_vector(3 downto 0);
signal S_9_c13 :  std_logic_vector(3 downto 0);
signal R_9_c13 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
            end if;
            if ce_4 = '1' then
               Cin_0_c4 <= Cin_0_c3;
               X_0_c4 <= X_0_c3;
               Y_0_c4 <= Y_0_c3;
               X_1_c4 <= X_1_c3;
               Y_1_c4 <= Y_1_c3;
               X_2_c4 <= X_2_c3;
               Y_2_c4 <= Y_2_c3;
               X_3_c4 <= X_3_c3;
               Y_3_c4 <= Y_3_c3;
               X_4_c4 <= X_4_c3;
               Y_4_c4 <= Y_4_c3;
               X_5_c4 <= X_5_c3;
               Y_5_c4 <= Y_5_c3;
               X_6_c4 <= X_6_c3;
               Y_6_c4 <= Y_6_c3;
               X_7_c4 <= X_7_c3;
               Y_7_c4 <= Y_7_c3;
               X_8_c4 <= X_8_c3;
               Y_8_c4 <= Y_8_c3;
               X_9_c4 <= X_9_c3;
               Y_9_c4 <= Y_9_c3;
            end if;
            if ce_5 = '1' then
               R_0_c5 <= R_0_c4;
               Cin_1_c5 <= Cin_1_c4;
               X_1_c5 <= X_1_c4;
               Y_1_c5 <= Y_1_c4;
               X_2_c5 <= X_2_c4;
               Y_2_c5 <= Y_2_c4;
               X_3_c5 <= X_3_c4;
               Y_3_c5 <= Y_3_c4;
               X_4_c5 <= X_4_c4;
               Y_4_c5 <= Y_4_c4;
               X_5_c5 <= X_5_c4;
               Y_5_c5 <= Y_5_c4;
               X_6_c5 <= X_6_c4;
               Y_6_c5 <= Y_6_c4;
               X_7_c5 <= X_7_c4;
               Y_7_c5 <= Y_7_c4;
               X_8_c5 <= X_8_c4;
               Y_8_c5 <= Y_8_c4;
               X_9_c5 <= X_9_c4;
               Y_9_c5 <= Y_9_c4;
            end if;
            if ce_6 = '1' then
               R_0_c6 <= R_0_c5;
               R_1_c6 <= R_1_c5;
               Cin_2_c6 <= Cin_2_c5;
               X_2_c6 <= X_2_c5;
               Y_2_c6 <= Y_2_c5;
               X_3_c6 <= X_3_c5;
               Y_3_c6 <= Y_3_c5;
               X_4_c6 <= X_4_c5;
               Y_4_c6 <= Y_4_c5;
               X_5_c6 <= X_5_c5;
               Y_5_c6 <= Y_5_c5;
               X_6_c6 <= X_6_c5;
               Y_6_c6 <= Y_6_c5;
               X_7_c6 <= X_7_c5;
               Y_7_c6 <= Y_7_c5;
               X_8_c6 <= X_8_c5;
               Y_8_c6 <= Y_8_c5;
               X_9_c6 <= X_9_c5;
               Y_9_c6 <= Y_9_c5;
            end if;
            if ce_7 = '1' then
               R_0_c7 <= R_0_c6;
               R_1_c7 <= R_1_c6;
               R_2_c7 <= R_2_c6;
               Cin_3_c7 <= Cin_3_c6;
               X_3_c7 <= X_3_c6;
               Y_3_c7 <= Y_3_c6;
               X_4_c7 <= X_4_c6;
               Y_4_c7 <= Y_4_c6;
               X_5_c7 <= X_5_c6;
               Y_5_c7 <= Y_5_c6;
               X_6_c7 <= X_6_c6;
               Y_6_c7 <= Y_6_c6;
               X_7_c7 <= X_7_c6;
               Y_7_c7 <= Y_7_c6;
               X_8_c7 <= X_8_c6;
               Y_8_c7 <= Y_8_c6;
               X_9_c7 <= X_9_c6;
               Y_9_c7 <= Y_9_c6;
            end if;
            if ce_8 = '1' then
               R_0_c8 <= R_0_c7;
               R_1_c8 <= R_1_c7;
               R_2_c8 <= R_2_c7;
               R_3_c8 <= R_3_c7;
               Cin_4_c8 <= Cin_4_c7;
               X_4_c8 <= X_4_c7;
               Y_4_c8 <= Y_4_c7;
               X_5_c8 <= X_5_c7;
               Y_5_c8 <= Y_5_c7;
               X_6_c8 <= X_6_c7;
               Y_6_c8 <= Y_6_c7;
               X_7_c8 <= X_7_c7;
               Y_7_c8 <= Y_7_c7;
               X_8_c8 <= X_8_c7;
               Y_8_c8 <= Y_8_c7;
               X_9_c8 <= X_9_c7;
               Y_9_c8 <= Y_9_c7;
            end if;
            if ce_9 = '1' then
               R_0_c9 <= R_0_c8;
               R_1_c9 <= R_1_c8;
               R_2_c9 <= R_2_c8;
               R_3_c9 <= R_3_c8;
               R_4_c9 <= R_4_c8;
               Cin_5_c9 <= Cin_5_c8;
               X_5_c9 <= X_5_c8;
               Y_5_c9 <= Y_5_c8;
               X_6_c9 <= X_6_c8;
               Y_6_c9 <= Y_6_c8;
               X_7_c9 <= X_7_c8;
               Y_7_c9 <= Y_7_c8;
               X_8_c9 <= X_8_c8;
               Y_8_c9 <= Y_8_c8;
               X_9_c9 <= X_9_c8;
               Y_9_c9 <= Y_9_c8;
            end if;
            if ce_10 = '1' then
               R_0_c10 <= R_0_c9;
               R_1_c10 <= R_1_c9;
               R_2_c10 <= R_2_c9;
               R_3_c10 <= R_3_c9;
               R_4_c10 <= R_4_c9;
               R_5_c10 <= R_5_c9;
               Cin_6_c10 <= Cin_6_c9;
               X_6_c10 <= X_6_c9;
               Y_6_c10 <= Y_6_c9;
               X_7_c10 <= X_7_c9;
               Y_7_c10 <= Y_7_c9;
               X_8_c10 <= X_8_c9;
               Y_8_c10 <= Y_8_c9;
               X_9_c10 <= X_9_c9;
               Y_9_c10 <= Y_9_c9;
            end if;
            if ce_11 = '1' then
               R_0_c11 <= R_0_c10;
               R_1_c11 <= R_1_c10;
               R_2_c11 <= R_2_c10;
               R_3_c11 <= R_3_c10;
               R_4_c11 <= R_4_c10;
               R_5_c11 <= R_5_c10;
               R_6_c11 <= R_6_c10;
               Cin_7_c11 <= Cin_7_c10;
               X_7_c11 <= X_7_c10;
               Y_7_c11 <= Y_7_c10;
               X_8_c11 <= X_8_c10;
               Y_8_c11 <= Y_8_c10;
               X_9_c11 <= X_9_c10;
               Y_9_c11 <= Y_9_c10;
            end if;
            if ce_12 = '1' then
               R_0_c12 <= R_0_c11;
               R_1_c12 <= R_1_c11;
               R_2_c12 <= R_2_c11;
               R_3_c12 <= R_3_c11;
               R_4_c12 <= R_4_c11;
               R_5_c12 <= R_5_c11;
               R_6_c12 <= R_6_c11;
               R_7_c12 <= R_7_c11;
               Cin_8_c12 <= Cin_8_c11;
               X_8_c12 <= X_8_c11;
               Y_8_c12 <= Y_8_c11;
               X_9_c12 <= X_9_c11;
               Y_9_c12 <= Y_9_c11;
            end if;
            if ce_13 = '1' then
               R_0_c13 <= R_0_c12;
               R_1_c13 <= R_1_c12;
               R_2_c13 <= R_2_c12;
               R_3_c13 <= R_3_c12;
               R_4_c13 <= R_4_c12;
               R_5_c13 <= R_5_c12;
               R_6_c13 <= R_6_c12;
               R_7_c13 <= R_7_c12;
               R_8_c13 <= R_8_c12;
               Cin_9_c13 <= Cin_9_c12;
               X_9_c13 <= X_9_c12;
               Y_9_c13 <= Y_9_c12;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c3 <= '0' & X(2 downto 0);
   Y_0_c3 <= '0' & Y(2 downto 0);
   S_0_c4 <= X_0_c4 + Y_0_c4 + Cin_0_c4;
   R_0_c4 <= S_0_c4(2 downto 0);
   Cin_1_c4 <= S_0_c4(3);
   X_1_c3 <= '0' & X(5 downto 3);
   Y_1_c3 <= '0' & Y(5 downto 3);
   S_1_c5 <= X_1_c5 + Y_1_c5 + Cin_1_c5;
   R_1_c5 <= S_1_c5(2 downto 0);
   Cin_2_c5 <= S_1_c5(3);
   X_2_c3 <= '0' & X(8 downto 6);
   Y_2_c3 <= '0' & Y(8 downto 6);
   S_2_c6 <= X_2_c6 + Y_2_c6 + Cin_2_c6;
   R_2_c6 <= S_2_c6(2 downto 0);
   Cin_3_c6 <= S_2_c6(3);
   X_3_c3 <= '0' & X(11 downto 9);
   Y_3_c3 <= '0' & Y(11 downto 9);
   S_3_c7 <= X_3_c7 + Y_3_c7 + Cin_3_c7;
   R_3_c7 <= S_3_c7(2 downto 0);
   Cin_4_c7 <= S_3_c7(3);
   X_4_c3 <= '0' & X(14 downto 12);
   Y_4_c3 <= '0' & Y(14 downto 12);
   S_4_c8 <= X_4_c8 + Y_4_c8 + Cin_4_c8;
   R_4_c8 <= S_4_c8(2 downto 0);
   Cin_5_c8 <= S_4_c8(3);
   X_5_c3 <= '0' & X(17 downto 15);
   Y_5_c3 <= '0' & Y(17 downto 15);
   S_5_c9 <= X_5_c9 + Y_5_c9 + Cin_5_c9;
   R_5_c9 <= S_5_c9(2 downto 0);
   Cin_6_c9 <= S_5_c9(3);
   X_6_c3 <= '0' & X(20 downto 18);
   Y_6_c3 <= '0' & Y(20 downto 18);
   S_6_c10 <= X_6_c10 + Y_6_c10 + Cin_6_c10;
   R_6_c10 <= S_6_c10(2 downto 0);
   Cin_7_c10 <= S_6_c10(3);
   X_7_c3 <= '0' & X(23 downto 21);
   Y_7_c3 <= '0' & Y(23 downto 21);
   S_7_c11 <= X_7_c11 + Y_7_c11 + Cin_7_c11;
   R_7_c11 <= S_7_c11(2 downto 0);
   Cin_8_c11 <= S_7_c11(3);
   X_8_c3 <= '0' & X(26 downto 24);
   Y_8_c3 <= '0' & Y(26 downto 24);
   S_8_c12 <= X_8_c12 + Y_8_c12 + Cin_8_c12;
   R_8_c12 <= S_8_c12(2 downto 0);
   Cin_9_c12 <= S_8_c12(3);
   X_9_c3 <= '0' & X(29 downto 27);
   Y_9_c3 <= '0' & Y(29 downto 27);
   S_9_c13 <= X_9_c13 + Y_9_c13 + Cin_9_c13;
   R_9_c13 <= S_9_c13(2 downto 0);
   R <= R_9_c13 & R_8_c13 & R_7_c13 & R_6_c13 & R_5_c13 & R_4_c13 & R_3_c13 & R_2_c13 & R_1_c13 & R_0_c13 ;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_24x24_48_Freq800_uid5
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 13 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_24x24_48_Freq800_uid5 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13 : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_24x24_48_Freq800_uid5 is
   component DSPBlock_17x24_Freq800_uid9 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid11 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid13 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid18 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid23 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid35 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid37 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid42 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid47 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid49 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid54 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid59 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid61 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid66 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid73 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid78 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid83 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid85 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid90 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid95 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid97 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid102 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid107 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid109 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid114 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid119 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid126 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid131 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid133 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid138 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq800_uid143 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid145 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid150 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq800_uid156 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq800_uid160 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_14_3_Freq800_uid164 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq800_uid170 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_30_Freq800_uid352 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13 : in std_logic;
             X : in  std_logic_vector(29 downto 0);
             Y : in  std_logic_vector(29 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(29 downto 0)   );
   end component;

signal XX_m6_c0 :  std_logic_vector(23 downto 0);
signal YY_m6_c0 :  std_logic_vector(23 downto 0);
signal tile_0_X_c0 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_0_output_c2 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w0_0_c2, bh7_w0_0_c3 :  std_logic;
signal bh7_w1_0_c2, bh7_w1_0_c3 :  std_logic;
signal bh7_w2_0_c2, bh7_w2_0_c3 :  std_logic;
signal bh7_w3_0_c2, bh7_w3_0_c3 :  std_logic;
signal bh7_w4_0_c2, bh7_w4_0_c3 :  std_logic;
signal bh7_w5_0_c2, bh7_w5_0_c3 :  std_logic;
signal bh7_w6_0_c2, bh7_w6_0_c3 :  std_logic;
signal bh7_w7_0_c2, bh7_w7_0_c3 :  std_logic;
signal bh7_w8_0_c2, bh7_w8_0_c3 :  std_logic;
signal bh7_w9_0_c2, bh7_w9_0_c3 :  std_logic;
signal bh7_w10_0_c2, bh7_w10_0_c3 :  std_logic;
signal bh7_w11_0_c2, bh7_w11_0_c3 :  std_logic;
signal bh7_w12_0_c2, bh7_w12_0_c3 :  std_logic;
signal bh7_w13_0_c2, bh7_w13_0_c3 :  std_logic;
signal bh7_w14_0_c2, bh7_w14_0_c3 :  std_logic;
signal bh7_w15_0_c2, bh7_w15_0_c3 :  std_logic;
signal bh7_w16_0_c2, bh7_w16_0_c3 :  std_logic;
signal bh7_w17_0_c2 :  std_logic;
signal bh7_w18_0_c2 :  std_logic;
signal bh7_w19_0_c2 :  std_logic;
signal bh7_w20_0_c2 :  std_logic;
signal bh7_w21_0_c2 :  std_logic;
signal bh7_w22_0_c2 :  std_logic;
signal bh7_w23_0_c2 :  std_logic;
signal bh7_w24_0_c2 :  std_logic;
signal bh7_w25_0_c2 :  std_logic;
signal bh7_w26_0_c2, bh7_w26_0_c3 :  std_logic;
signal bh7_w27_0_c2, bh7_w27_0_c3 :  std_logic;
signal bh7_w28_0_c2, bh7_w28_0_c3 :  std_logic;
signal bh7_w29_0_c2, bh7_w29_0_c3 :  std_logic;
signal bh7_w30_0_c2, bh7_w30_0_c3 :  std_logic;
signal bh7_w31_0_c2, bh7_w31_0_c3 :  std_logic;
signal bh7_w32_0_c2, bh7_w32_0_c3 :  std_logic;
signal bh7_w33_0_c2, bh7_w33_0_c3 :  std_logic;
signal bh7_w34_0_c2, bh7_w34_0_c3 :  std_logic;
signal bh7_w35_0_c2, bh7_w35_0_c3 :  std_logic;
signal bh7_w36_0_c2, bh7_w36_0_c3 :  std_logic;
signal bh7_w37_0_c2, bh7_w37_0_c3 :  std_logic;
signal bh7_w38_0_c2, bh7_w38_0_c3 :  std_logic;
signal bh7_w39_0_c2, bh7_w39_0_c3 :  std_logic;
signal bh7_w40_0_c2, bh7_w40_0_c3 :  std_logic;
signal tile_1_X_c0 :  std_logic_vector(0 downto 0);
signal tile_1_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_1_output_c0 :  std_logic_vector(1 downto 0);
signal tile_1_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w45_0_c0 :  std_logic;
signal bh7_w46_0_c0 :  std_logic;
signal tile_2_X_c0 :  std_logic_vector(2 downto 0);
signal tile_2_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_2_output_c0 :  std_logic_vector(4 downto 0);
signal tile_2_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w42_0_c0 :  std_logic;
signal bh7_w43_0_c0 :  std_logic;
signal bh7_w44_0_c0 :  std_logic;
signal bh7_w45_1_c0 :  std_logic;
signal bh7_w46_1_c0 :  std_logic;
signal tile_3_X_c0 :  std_logic_vector(2 downto 0);
signal tile_3_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_3_output_c0 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w39_1_c0 :  std_logic;
signal bh7_w40_1_c0 :  std_logic;
signal bh7_w41_0_c0 :  std_logic;
signal bh7_w42_1_c0 :  std_logic;
signal bh7_w43_1_c0 :  std_logic;
signal tile_4_X_c0 :  std_logic_vector(0 downto 0);
signal tile_4_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_4_output_c0 :  std_logic_vector(1 downto 0);
signal tile_4_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w43_2_c0 :  std_logic;
signal bh7_w44_1_c0 :  std_logic;
signal tile_5_X_c0 :  std_logic_vector(2 downto 0);
signal tile_5_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_5_output_c0 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w40_2_c0 :  std_logic;
signal bh7_w41_1_c0 :  std_logic;
signal bh7_w42_2_c0 :  std_logic;
signal bh7_w43_3_c0 :  std_logic;
signal bh7_w44_2_c0, bh7_w44_2_c1 :  std_logic;
signal tile_6_X_c0 :  std_logic_vector(2 downto 0);
signal tile_6_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_6_output_c0 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w37_1_c0 :  std_logic;
signal bh7_w38_1_c0 :  std_logic;
signal bh7_w39_2_c0 :  std_logic;
signal bh7_w40_3_c0 :  std_logic;
signal bh7_w41_2_c0 :  std_logic;
signal tile_7_X_c0 :  std_logic_vector(0 downto 0);
signal tile_7_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_7_output_c0 :  std_logic_vector(1 downto 0);
signal tile_7_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w41_3_c0 :  std_logic;
signal bh7_w42_3_c0 :  std_logic;
signal tile_8_X_c0 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_8_output_c0 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w38_2_c0 :  std_logic;
signal bh7_w39_3_c0 :  std_logic;
signal bh7_w40_4_c0 :  std_logic;
signal bh7_w41_4_c0, bh7_w41_4_c1 :  std_logic;
signal bh7_w42_4_c0 :  std_logic;
signal tile_9_X_c0 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_9_output_c0 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w35_1_c0 :  std_logic;
signal bh7_w36_1_c0 :  std_logic;
signal bh7_w37_2_c0 :  std_logic;
signal bh7_w38_3_c0 :  std_logic;
signal bh7_w39_4_c0 :  std_logic;
signal tile_10_X_c0 :  std_logic_vector(0 downto 0);
signal tile_10_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_10_output_c0 :  std_logic_vector(1 downto 0);
signal tile_10_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w39_5_c0 :  std_logic;
signal bh7_w40_5_c0 :  std_logic;
signal tile_11_X_c0 :  std_logic_vector(2 downto 0);
signal tile_11_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_11_output_c0 :  std_logic_vector(4 downto 0);
signal tile_11_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w36_2_c0 :  std_logic;
signal bh7_w37_3_c0 :  std_logic;
signal bh7_w38_4_c0 :  std_logic;
signal bh7_w39_6_c0 :  std_logic;
signal bh7_w40_6_c0 :  std_logic;
signal tile_12_X_c0 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_12_output_c0 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w33_1_c0 :  std_logic;
signal bh7_w34_1_c0 :  std_logic;
signal bh7_w35_2_c0 :  std_logic;
signal bh7_w36_3_c0 :  std_logic;
signal bh7_w37_4_c0 :  std_logic;
signal tile_13_X_c0 :  std_logic_vector(0 downto 0);
signal tile_13_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_13_output_c0 :  std_logic_vector(1 downto 0);
signal tile_13_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w37_5_c0 :  std_logic;
signal bh7_w38_5_c0 :  std_logic;
signal tile_14_X_c0 :  std_logic_vector(2 downto 0);
signal tile_14_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_14_output_c0 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w34_2_c0 :  std_logic;
signal bh7_w35_3_c0 :  std_logic;
signal bh7_w36_4_c0 :  std_logic;
signal bh7_w37_6_c0 :  std_logic;
signal bh7_w38_6_c0 :  std_logic;
signal tile_15_X_c0 :  std_logic_vector(2 downto 0);
signal tile_15_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_15_output_c0 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w31_1_c0 :  std_logic;
signal bh7_w32_1_c0 :  std_logic;
signal bh7_w33_2_c0 :  std_logic;
signal bh7_w34_3_c0 :  std_logic;
signal bh7_w35_4_c0 :  std_logic;
signal tile_16_X_c0 :  std_logic_vector(0 downto 0);
signal tile_16_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_16_output_c0 :  std_logic_vector(1 downto 0);
signal tile_16_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w35_5_c0 :  std_logic;
signal bh7_w36_5_c0 :  std_logic;
signal tile_17_X_c0 :  std_logic_vector(2 downto 0);
signal tile_17_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_17_output_c0 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w32_2_c0 :  std_logic;
signal bh7_w33_3_c0 :  std_logic;
signal bh7_w34_4_c0 :  std_logic;
signal bh7_w35_6_c0 :  std_logic;
signal bh7_w36_6_c0 :  std_logic;
signal tile_18_X_c0 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_18_output_c0 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w29_1_c0 :  std_logic;
signal bh7_w30_1_c0 :  std_logic;
signal bh7_w31_2_c0 :  std_logic;
signal bh7_w32_3_c0 :  std_logic;
signal bh7_w33_4_c0 :  std_logic;
signal tile_19_X_c0 :  std_logic_vector(0 downto 0);
signal tile_19_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_19_output_c0 :  std_logic_vector(1 downto 0);
signal tile_19_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w33_5_c0 :  std_logic;
signal bh7_w34_5_c0 :  std_logic;
signal tile_20_X_c0 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_20_output_c0 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w30_2_c0 :  std_logic;
signal bh7_w31_3_c0 :  std_logic;
signal bh7_w32_4_c0 :  std_logic;
signal bh7_w33_6_c0 :  std_logic;
signal bh7_w34_6_c0 :  std_logic;
signal tile_21_X_c0 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_21_output_c0 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w27_1_c0 :  std_logic;
signal bh7_w28_1_c0 :  std_logic;
signal bh7_w29_2_c0 :  std_logic;
signal bh7_w30_3_c0 :  std_logic;
signal bh7_w31_4_c0 :  std_logic;
signal tile_22_X_c0 :  std_logic_vector(0 downto 0);
signal tile_22_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_22_output_c0 :  std_logic_vector(1 downto 0);
signal tile_22_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w31_5_c0 :  std_logic;
signal bh7_w32_5_c0 :  std_logic;
signal tile_23_X_c0 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_23_output_c0 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w28_2_c0 :  std_logic;
signal bh7_w29_3_c0 :  std_logic;
signal bh7_w30_4_c0 :  std_logic;
signal bh7_w31_6_c0 :  std_logic;
signal bh7_w32_6_c0 :  std_logic;
signal tile_24_X_c0 :  std_logic_vector(2 downto 0);
signal tile_24_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_24_output_c0 :  std_logic_vector(4 downto 0);
signal tile_24_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w25_1_c0 :  std_logic;
signal bh7_w26_1_c0 :  std_logic;
signal bh7_w27_2_c0 :  std_logic;
signal bh7_w28_3_c0 :  std_logic;
signal bh7_w29_4_c0 :  std_logic;
signal tile_25_X_c0 :  std_logic_vector(0 downto 0);
signal tile_25_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_25_output_c0 :  std_logic_vector(1 downto 0);
signal tile_25_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w29_5_c0 :  std_logic;
signal bh7_w30_5_c0 :  std_logic;
signal tile_26_X_c0 :  std_logic_vector(2 downto 0);
signal tile_26_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_26_output_c0 :  std_logic_vector(4 downto 0);
signal tile_26_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w26_2_c0 :  std_logic;
signal bh7_w27_3_c0 :  std_logic;
signal bh7_w28_4_c0 :  std_logic;
signal bh7_w29_6_c0 :  std_logic;
signal bh7_w30_6_c0 :  std_logic;
signal tile_27_X_c0 :  std_logic_vector(2 downto 0);
signal tile_27_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_27_output_c0 :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w23_1_c0 :  std_logic;
signal bh7_w24_1_c0 :  std_logic;
signal bh7_w25_2_c0 :  std_logic;
signal bh7_w26_3_c0 :  std_logic;
signal bh7_w27_4_c0 :  std_logic;
signal tile_28_X_c0 :  std_logic_vector(0 downto 0);
signal tile_28_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_28_output_c0 :  std_logic_vector(1 downto 0);
signal tile_28_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w27_5_c0 :  std_logic;
signal bh7_w28_5_c0 :  std_logic;
signal tile_29_X_c0 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_29_output_c0 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w24_2_c0 :  std_logic;
signal bh7_w25_3_c0 :  std_logic;
signal bh7_w26_4_c0 :  std_logic;
signal bh7_w27_6_c0 :  std_logic;
signal bh7_w28_6_c0 :  std_logic;
signal tile_30_X_c0 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_30_output_c0 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w21_1_c0 :  std_logic;
signal bh7_w22_1_c0 :  std_logic;
signal bh7_w23_2_c0 :  std_logic;
signal bh7_w24_3_c0 :  std_logic;
signal bh7_w25_4_c0 :  std_logic;
signal tile_31_X_c0 :  std_logic_vector(0 downto 0);
signal tile_31_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_31_output_c0 :  std_logic_vector(1 downto 0);
signal tile_31_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w25_5_c0 :  std_logic;
signal bh7_w26_5_c0 :  std_logic;
signal tile_32_X_c0 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_32_output_c0 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w22_2_c0 :  std_logic;
signal bh7_w23_3_c0 :  std_logic;
signal bh7_w24_4_c0 :  std_logic;
signal bh7_w25_6_c0 :  std_logic;
signal bh7_w26_6_c0 :  std_logic;
signal tile_33_X_c0 :  std_logic_vector(2 downto 0);
signal tile_33_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_33_output_c0 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w19_1_c0 :  std_logic;
signal bh7_w20_1_c0 :  std_logic;
signal bh7_w21_2_c0 :  std_logic;
signal bh7_w22_3_c0 :  std_logic;
signal bh7_w23_4_c0 :  std_logic;
signal tile_34_X_c0 :  std_logic_vector(0 downto 0);
signal tile_34_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_34_output_c0 :  std_logic_vector(1 downto 0);
signal tile_34_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w23_5_c0 :  std_logic;
signal bh7_w24_5_c0 :  std_logic;
signal tile_35_X_c0 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_35_output_c0 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w20_2_c0 :  std_logic;
signal bh7_w21_3_c0 :  std_logic;
signal bh7_w22_4_c0 :  std_logic;
signal bh7_w23_6_c0 :  std_logic;
signal bh7_w24_6_c0 :  std_logic;
signal tile_36_X_c0 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_36_output_c0 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w17_1_c0, bh7_w17_1_c1, bh7_w17_1_c2 :  std_logic;
signal bh7_w18_1_c0 :  std_logic;
signal bh7_w19_2_c0 :  std_logic;
signal bh7_w20_3_c0 :  std_logic;
signal bh7_w21_4_c0 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid157_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid157_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w18_2_c1, bh7_w18_2_c2 :  std_logic;
signal bh7_w19_3_c1, bh7_w19_3_c2 :  std_logic;
signal bh7_w20_4_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_copy158_c0, Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_copy158_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid161_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w20_5_c1 :  std_logic;
signal bh7_w21_5_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_copy162_c0, Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_copy162_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid165_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid165_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_6_c1 :  std_logic;
signal bh7_w22_5_c1 :  std_logic;
signal bh7_w23_7_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_copy166_c0, Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_copy166_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid167_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w22_6_c1 :  std_logic;
signal bh7_w23_8_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_copy168_c0, Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_copy168_c1 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid171_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w23_9_c1 :  std_logic;
signal bh7_w24_7_c1 :  std_logic;
signal bh7_w25_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_copy172_c0, Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_copy172_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid173_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w24_8_c1 :  std_logic;
signal bh7_w25_8_c1 :  std_logic;
signal bh7_w26_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_copy174_c0, Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_copy174_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid175_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w25_9_c1 :  std_logic;
signal bh7_w26_8_c1 :  std_logic;
signal bh7_w27_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_copy176_c0, Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_copy176_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid177_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w26_9_c1 :  std_logic;
signal bh7_w27_8_c1 :  std_logic;
signal bh7_w28_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_copy178_c0, Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_copy178_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid179_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w27_9_c1 :  std_logic;
signal bh7_w28_8_c1 :  std_logic;
signal bh7_w29_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_copy180_c0, Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_copy180_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid181_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w28_9_c1 :  std_logic;
signal bh7_w29_8_c1 :  std_logic;
signal bh7_w30_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_copy182_c0, Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_copy182_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid183_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_9_c1 :  std_logic;
signal bh7_w30_8_c1 :  std_logic;
signal bh7_w31_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_copy184_c0, Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_copy184_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid185_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w30_9_c1 :  std_logic;
signal bh7_w31_8_c1 :  std_logic;
signal bh7_w32_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_copy186_c0, Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_copy186_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid187_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_9_c1 :  std_logic;
signal bh7_w32_8_c1 :  std_logic;
signal bh7_w33_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_copy188_c0, Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_copy188_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid189_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w32_9_c1 :  std_logic;
signal bh7_w33_8_c1 :  std_logic;
signal bh7_w34_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_copy190_c0, Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_copy190_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid191_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_9_c1 :  std_logic;
signal bh7_w34_8_c1 :  std_logic;
signal bh7_w35_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_copy192_c0, Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_copy192_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid193_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w34_9_c1 :  std_logic;
signal bh7_w35_8_c1 :  std_logic;
signal bh7_w36_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_copy194_c0, Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_copy194_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid195_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w35_9_c1 :  std_logic;
signal bh7_w36_8_c1 :  std_logic;
signal bh7_w37_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_copy196_c0, Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_copy196_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid197_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w36_9_c1 :  std_logic;
signal bh7_w37_8_c1 :  std_logic;
signal bh7_w38_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_copy198_c0, Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_copy198_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid199_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w37_9_c1 :  std_logic;
signal bh7_w38_8_c1 :  std_logic;
signal bh7_w39_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_copy200_c0, Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_copy200_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid201_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w38_9_c1 :  std_logic;
signal bh7_w39_8_c1 :  std_logic;
signal bh7_w40_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_copy202_c0, Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_copy202_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid203_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w39_9_c1 :  std_logic;
signal bh7_w40_8_c1 :  std_logic;
signal bh7_w41_5_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_copy204_c0, Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_copy204_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid205_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w40_9_c1 :  std_logic;
signal bh7_w41_6_c1 :  std_logic;
signal bh7_w42_5_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_copy206_c0, Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_copy206_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid207_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid207_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w41_7_c1 :  std_logic;
signal bh7_w42_6_c1 :  std_logic;
signal bh7_w43_4_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_copy208_c0, Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_copy208_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid209_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid209_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w42_7_c1 :  std_logic;
signal bh7_w43_5_c1 :  std_logic;
signal bh7_w44_3_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_copy210_c0, Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_copy210_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid211_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid211_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w43_6_c1 :  std_logic;
signal bh7_w44_4_c1 :  std_logic;
signal bh7_w45_2_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_copy212_c0, Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_copy212_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid213_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid213_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w45_3_c1 :  std_logic;
signal bh7_w46_2_c1 :  std_logic;
signal bh7_w47_0_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_copy214_c0, Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_copy214_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid215_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid215_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid215_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w20_6_c1, bh7_w20_6_c2 :  std_logic;
signal bh7_w21_7_c1, bh7_w21_7_c2 :  std_logic;
signal bh7_w22_7_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid215_Out0_copy216_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid217_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid217_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w22_8_c1 :  std_logic;
signal bh7_w23_10_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid160_bh7_uid217_Out0_copy218_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid219_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid219_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid219_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w23_11_c1 :  std_logic;
signal bh7_w24_9_c1, bh7_w24_9_c2 :  std_logic;
signal bh7_w25_10_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid219_Out0_copy220_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid221_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid221_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid221_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w25_11_c1 :  std_logic;
signal bh7_w26_10_c1 :  std_logic;
signal bh7_w27_10_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid221_Out0_copy222_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid223_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid223_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid223_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w27_11_c1 :  std_logic;
signal bh7_w28_10_c1 :  std_logic;
signal bh7_w29_10_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid223_Out0_copy224_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid225_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid225_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid225_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_11_c1 :  std_logic;
signal bh7_w30_10_c1 :  std_logic;
signal bh7_w31_10_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid225_Out0_copy226_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid227_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid227_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid227_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_11_c1 :  std_logic;
signal bh7_w32_10_c1 :  std_logic;
signal bh7_w33_10_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid227_Out0_copy228_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid229_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid229_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid229_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_11_c1 :  std_logic;
signal bh7_w34_10_c1 :  std_logic;
signal bh7_w35_10_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid229_Out0_copy230_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid231_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid231_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid231_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w35_11_c1 :  std_logic;
signal bh7_w36_10_c1 :  std_logic;
signal bh7_w37_10_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid231_Out0_copy232_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid233_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid233_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid233_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w37_11_c1 :  std_logic;
signal bh7_w38_10_c1 :  std_logic;
signal bh7_w39_10_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid233_Out0_copy234_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid235_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid235_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid235_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w39_11_c1 :  std_logic;
signal bh7_w40_10_c1 :  std_logic;
signal bh7_w41_8_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid235_Out0_copy236_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid237_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid237_In1_c0, Compressor_14_3_Freq800_uid164_bh7_uid237_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid237_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w41_9_c1 :  std_logic;
signal bh7_w42_8_c1 :  std_logic;
signal bh7_w43_7_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid237_Out0_copy238_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid239_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid239_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w42_9_c1 :  std_logic;
signal bh7_w43_8_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid160_bh7_uid239_Out0_copy240_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid241_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid241_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid241_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w43_9_c1 :  std_logic;
signal bh7_w44_5_c1 :  std_logic;
signal bh7_w45_4_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid241_Out0_copy242_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid243_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid243_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid243_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w45_5_c1 :  std_logic;
signal bh7_w46_3_c1 :  std_logic;
signal bh7_w47_1_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid243_Out0_copy244_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid245_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid245_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w22_9_c2 :  std_logic;
signal bh7_w23_12_c2 :  std_logic;
signal bh7_w24_10_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_copy246_c1, Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_copy246_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid247_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid247_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w25_12_c2 :  std_logic;
signal bh7_w26_11_c2 :  std_logic;
signal bh7_w27_12_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_copy248_c1, Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_copy248_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid249_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid249_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w27_13_c2 :  std_logic;
signal bh7_w28_11_c2 :  std_logic;
signal bh7_w29_12_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_copy250_c1, Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_copy250_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid251_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid251_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w29_13_c2 :  std_logic;
signal bh7_w30_11_c2 :  std_logic;
signal bh7_w31_12_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_copy252_c1, Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_copy252_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid253_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid253_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w31_13_c2 :  std_logic;
signal bh7_w32_11_c2 :  std_logic;
signal bh7_w33_12_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_copy254_c1, Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_copy254_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid255_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid255_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w33_13_c2 :  std_logic;
signal bh7_w34_11_c2 :  std_logic;
signal bh7_w35_12_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_copy256_c1, Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_copy256_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid257_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid257_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w35_13_c2 :  std_logic;
signal bh7_w36_11_c2 :  std_logic;
signal bh7_w37_12_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_copy258_c1, Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_copy258_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid259_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid259_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w37_13_c2 :  std_logic;
signal bh7_w38_11_c2 :  std_logic;
signal bh7_w39_12_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_copy260_c1, Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_copy260_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid261_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid261_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w39_13_c2 :  std_logic;
signal bh7_w40_11_c2 :  std_logic;
signal bh7_w41_10_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_copy262_c1, Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_copy262_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid263_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid263_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w41_11_c2 :  std_logic;
signal bh7_w42_10_c2 :  std_logic;
signal bh7_w43_10_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_copy264_c1, Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_copy264_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid265_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid265_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w43_11_c2 :  std_logic;
signal bh7_w44_6_c2 :  std_logic;
signal bh7_w45_6_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_copy266_c1, Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_copy266_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid267_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid267_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w45_7_c2 :  std_logic;
signal bh7_w46_4_c2 :  std_logic;
signal bh7_w47_2_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_copy268_c1, Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_copy268_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid269_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid269_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w47_3_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid160_bh7_uid269_Out0_copy270_c1, Compressor_3_2_Freq800_uid160_bh7_uid269_Out0_copy270_c2 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid271_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid271_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid271_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w24_11_c2 :  std_logic;
signal bh7_w25_13_c2 :  std_logic;
signal bh7_w26_12_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid271_Out0_copy272_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid273_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid273_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid273_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w27_14_c2 :  std_logic;
signal bh7_w28_12_c2, bh7_w28_12_c3 :  std_logic;
signal bh7_w29_14_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid273_Out0_copy274_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid275_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid275_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid275_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w29_15_c2 :  std_logic;
signal bh7_w30_12_c2 :  std_logic;
signal bh7_w31_14_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid275_Out0_copy276_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid277_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid277_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid277_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w31_15_c2 :  std_logic;
signal bh7_w32_12_c2 :  std_logic;
signal bh7_w33_14_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid277_Out0_copy278_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid279_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid279_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid279_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w33_15_c2 :  std_logic;
signal bh7_w34_12_c2 :  std_logic;
signal bh7_w35_14_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid279_Out0_copy280_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid281_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid281_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid281_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w35_15_c2 :  std_logic;
signal bh7_w36_12_c2 :  std_logic;
signal bh7_w37_14_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid281_Out0_copy282_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid283_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid283_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid283_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w37_15_c2 :  std_logic;
signal bh7_w38_12_c2 :  std_logic;
signal bh7_w39_14_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid283_Out0_copy284_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid285_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid285_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid285_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w39_15_c2 :  std_logic;
signal bh7_w40_12_c2 :  std_logic;
signal bh7_w41_12_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid285_Out0_copy286_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid287_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid287_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid287_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w41_13_c2 :  std_logic;
signal bh7_w42_11_c2 :  std_logic;
signal bh7_w43_12_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid287_Out0_copy288_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid289_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid289_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid289_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w43_13_c2 :  std_logic;
signal bh7_w44_7_c2 :  std_logic;
signal bh7_w45_8_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid289_Out0_copy290_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid291_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid291_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid291_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w45_9_c2 :  std_logic;
signal bh7_w46_5_c2 :  std_logic;
signal bh7_w47_4_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid291_Out0_copy292_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid293_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid293_In1_c0, Compressor_14_3_Freq800_uid164_bh7_uid293_In1_c1, Compressor_14_3_Freq800_uid164_bh7_uid293_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid293_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w47_5_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid293_Out0_copy294_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid295_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid295_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w26_13_c3 :  std_logic;
signal bh7_w27_15_c3 :  std_logic;
signal bh7_w28_13_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_copy296_c2, Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_copy296_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid297_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid297_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w29_16_c3 :  std_logic;
signal bh7_w30_13_c3 :  std_logic;
signal bh7_w31_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_copy298_c2, Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_copy298_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid299_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid299_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w31_17_c3 :  std_logic;
signal bh7_w32_13_c3 :  std_logic;
signal bh7_w33_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_copy300_c2, Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_copy300_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid301_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid301_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w33_17_c3 :  std_logic;
signal bh7_w34_13_c3 :  std_logic;
signal bh7_w35_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_copy302_c2, Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_copy302_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid303_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid303_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w35_17_c3 :  std_logic;
signal bh7_w36_13_c3 :  std_logic;
signal bh7_w37_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_copy304_c2, Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_copy304_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid305_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid305_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w37_17_c3 :  std_logic;
signal bh7_w38_13_c3 :  std_logic;
signal bh7_w39_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_copy306_c2, Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_copy306_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid307_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid307_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w39_17_c3 :  std_logic;
signal bh7_w40_13_c3 :  std_logic;
signal bh7_w41_14_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_copy308_c2, Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_copy308_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid309_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid309_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w41_15_c3 :  std_logic;
signal bh7_w42_12_c3 :  std_logic;
signal bh7_w43_14_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_copy310_c2, Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_copy310_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid311_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid311_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w43_15_c3 :  std_logic;
signal bh7_w44_8_c3 :  std_logic;
signal bh7_w45_10_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_copy312_c2, Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_copy312_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid313_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid313_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w45_11_c3 :  std_logic;
signal bh7_w46_6_c3 :  std_logic;
signal bh7_w47_6_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_copy314_c2, Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_copy314_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid315_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid315_In1_c0, Compressor_14_3_Freq800_uid164_bh7_uid315_In1_c1, Compressor_14_3_Freq800_uid164_bh7_uid315_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid315_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w47_7_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid315_Out0_copy316_c2, Compressor_14_3_Freq800_uid164_bh7_uid315_Out0_copy316_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid317_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid317_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w17_2_c3 :  std_logic;
signal bh7_w18_3_c3 :  std_logic;
signal bh7_w19_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_copy318_c2, Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_copy318_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid319_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid319_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w19_5_c3 :  std_logic;
signal bh7_w20_7_c3 :  std_logic;
signal bh7_w21_8_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_copy320_c2, Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_copy320_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid321_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid321_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w21_9_c3 :  std_logic;
signal bh7_w22_10_c3 :  std_logic;
signal bh7_w23_13_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_copy322_c2, Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_copy322_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid323_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid323_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w23_14_c3 :  std_logic;
signal bh7_w24_12_c3 :  std_logic;
signal bh7_w25_14_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_copy324_c2, Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_copy324_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid325_In0_c2, Compressor_23_3_Freq800_uid156_bh7_uid325_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid325_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid325_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w25_15_c3 :  std_logic;
signal bh7_w26_14_c3 :  std_logic;
signal bh7_w27_16_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid325_Out0_copy326_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid327_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid327_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w27_17_c3 :  std_logic;
signal bh7_w28_14_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid160_bh7_uid327_Out0_copy328_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid329_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid329_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid329_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w28_15_c3 :  std_logic;
signal bh7_w29_17_c3 :  std_logic;
signal bh7_w30_14_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid329_Out0_copy330_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid331_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid160_bh7_uid331_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w30_15_c3 :  std_logic;
signal bh7_w31_18_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid160_bh7_uid331_Out0_copy332_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid333_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid333_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid333_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w31_19_c3 :  std_logic;
signal bh7_w32_14_c3 :  std_logic;
signal bh7_w33_18_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid333_Out0_copy334_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid335_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid335_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid335_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w33_19_c3 :  std_logic;
signal bh7_w34_14_c3 :  std_logic;
signal bh7_w35_18_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid335_Out0_copy336_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid337_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid337_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid337_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w35_19_c3 :  std_logic;
signal bh7_w36_14_c3 :  std_logic;
signal bh7_w37_18_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid337_Out0_copy338_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid339_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid339_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid339_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w37_19_c3 :  std_logic;
signal bh7_w38_14_c3 :  std_logic;
signal bh7_w39_18_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid339_Out0_copy340_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid341_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid341_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid156_bh7_uid341_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w39_19_c3 :  std_logic;
signal bh7_w40_14_c3 :  std_logic;
signal bh7_w41_16_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid156_bh7_uid341_Out0_copy342_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid343_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid343_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid343_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w41_17_c3 :  std_logic;
signal bh7_w42_13_c3 :  std_logic;
signal bh7_w43_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid343_Out0_copy344_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid345_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid345_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid345_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w43_17_c3 :  std_logic;
signal bh7_w44_9_c3 :  std_logic;
signal bh7_w45_12_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid345_Out0_copy346_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid347_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid347_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid347_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w45_13_c3 :  std_logic;
signal bh7_w46_7_c3 :  std_logic;
signal bh7_w47_8_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid347_Out0_copy348_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid349_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c0, Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c1, Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c2, Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid164_bh7_uid349_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w47_9_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid164_bh7_uid349_Out0_copy350_c3 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh7_18_c3, tmp_bitheapResult_bh7_18_c4, tmp_bitheapResult_bh7_18_c5, tmp_bitheapResult_bh7_18_c6, tmp_bitheapResult_bh7_18_c7, tmp_bitheapResult_bh7_18_c8, tmp_bitheapResult_bh7_18_c9, tmp_bitheapResult_bh7_18_c10, tmp_bitheapResult_bh7_18_c11, tmp_bitheapResult_bh7_18_c12, tmp_bitheapResult_bh7_18_c13 :  std_logic_vector(18 downto 0);
signal bitheapFinalAdd_bh7_In0_c3 :  std_logic_vector(29 downto 0);
signal bitheapFinalAdd_bh7_In1_c3 :  std_logic_vector(29 downto 0);
signal bitheapFinalAdd_bh7_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh7_Out_c13 :  std_logic_vector(29 downto 0);
signal bitheapResult_bh7_c13 :  std_logic_vector(47 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               bh7_w44_2_c1 <= bh7_w44_2_c0;
               bh7_w41_4_c1 <= bh7_w41_4_c0;
               bh7_w17_1_c1 <= bh7_w17_1_c0;
               Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_copy158_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_copy158_c0;
               Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_copy162_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_copy162_c0;
               Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_copy166_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_copy166_c0;
               Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_copy168_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_copy168_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_copy172_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_copy172_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_copy174_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_copy174_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_copy176_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_copy176_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_copy178_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_copy178_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_copy180_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_copy180_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_copy182_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_copy182_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_copy184_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_copy184_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_copy186_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_copy186_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_copy188_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_copy188_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_copy190_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_copy190_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_copy192_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_copy192_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_copy194_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_copy194_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_copy196_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_copy196_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_copy198_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_copy198_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_copy200_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_copy200_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_copy202_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_copy202_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_copy204_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_copy204_c0;
               Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_copy206_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_copy206_c0;
               Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_copy208_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_copy208_c0;
               Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_copy210_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_copy210_c0;
               Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_copy212_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_copy212_c0;
               Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_copy214_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_copy214_c0;
               Compressor_14_3_Freq800_uid164_bh7_uid237_In1_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid237_In1_c0;
               Compressor_14_3_Freq800_uid164_bh7_uid293_In1_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid293_In1_c0;
               Compressor_14_3_Freq800_uid164_bh7_uid315_In1_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid315_In1_c0;
               Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c0;
            end if;
            if ce_2 = '1' then
               bh7_w17_1_c2 <= bh7_w17_1_c1;
               bh7_w18_2_c2 <= bh7_w18_2_c1;
               bh7_w19_3_c2 <= bh7_w19_3_c1;
               bh7_w20_6_c2 <= bh7_w20_6_c1;
               bh7_w21_7_c2 <= bh7_w21_7_c1;
               bh7_w24_9_c2 <= bh7_w24_9_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_copy246_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_copy246_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_copy248_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_copy248_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_copy250_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_copy250_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_copy252_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_copy252_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_copy254_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_copy254_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_copy256_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_copy256_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_copy258_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_copy258_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_copy260_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_copy260_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_copy262_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_copy262_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_copy264_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_copy264_c1;
               Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_copy266_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_copy266_c1;
               Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_copy268_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_copy268_c1;
               Compressor_3_2_Freq800_uid160_bh7_uid269_Out0_copy270_c2 <= Compressor_3_2_Freq800_uid160_bh7_uid269_Out0_copy270_c1;
               Compressor_14_3_Freq800_uid164_bh7_uid293_In1_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid293_In1_c1;
               Compressor_14_3_Freq800_uid164_bh7_uid315_In1_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid315_In1_c1;
               Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c1;
            end if;
            if ce_3 = '1' then
               bh7_w0_0_c3 <= bh7_w0_0_c2;
               bh7_w1_0_c3 <= bh7_w1_0_c2;
               bh7_w2_0_c3 <= bh7_w2_0_c2;
               bh7_w3_0_c3 <= bh7_w3_0_c2;
               bh7_w4_0_c3 <= bh7_w4_0_c2;
               bh7_w5_0_c3 <= bh7_w5_0_c2;
               bh7_w6_0_c3 <= bh7_w6_0_c2;
               bh7_w7_0_c3 <= bh7_w7_0_c2;
               bh7_w8_0_c3 <= bh7_w8_0_c2;
               bh7_w9_0_c3 <= bh7_w9_0_c2;
               bh7_w10_0_c3 <= bh7_w10_0_c2;
               bh7_w11_0_c3 <= bh7_w11_0_c2;
               bh7_w12_0_c3 <= bh7_w12_0_c2;
               bh7_w13_0_c3 <= bh7_w13_0_c2;
               bh7_w14_0_c3 <= bh7_w14_0_c2;
               bh7_w15_0_c3 <= bh7_w15_0_c2;
               bh7_w16_0_c3 <= bh7_w16_0_c2;
               bh7_w26_0_c3 <= bh7_w26_0_c2;
               bh7_w27_0_c3 <= bh7_w27_0_c2;
               bh7_w28_0_c3 <= bh7_w28_0_c2;
               bh7_w29_0_c3 <= bh7_w29_0_c2;
               bh7_w30_0_c3 <= bh7_w30_0_c2;
               bh7_w31_0_c3 <= bh7_w31_0_c2;
               bh7_w32_0_c3 <= bh7_w32_0_c2;
               bh7_w33_0_c3 <= bh7_w33_0_c2;
               bh7_w34_0_c3 <= bh7_w34_0_c2;
               bh7_w35_0_c3 <= bh7_w35_0_c2;
               bh7_w36_0_c3 <= bh7_w36_0_c2;
               bh7_w37_0_c3 <= bh7_w37_0_c2;
               bh7_w38_0_c3 <= bh7_w38_0_c2;
               bh7_w39_0_c3 <= bh7_w39_0_c2;
               bh7_w40_0_c3 <= bh7_w40_0_c2;
               bh7_w28_12_c3 <= bh7_w28_12_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_copy296_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_copy296_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_copy298_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_copy298_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_copy300_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_copy300_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_copy302_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_copy302_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_copy304_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_copy304_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_copy306_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_copy306_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_copy308_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_copy308_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_copy310_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_copy310_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_copy312_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_copy312_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_copy314_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_copy314_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid315_Out0_copy316_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid315_Out0_copy316_c2;
               Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_copy318_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_copy318_c2;
               Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_copy320_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_copy320_c2;
               Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_copy322_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_copy322_c2;
               Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_copy324_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_copy324_c2;
               Compressor_23_3_Freq800_uid156_bh7_uid325_In0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid325_In0_c2;
               Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c2;
            end if;
            if ce_4 = '1' then
               tmp_bitheapResult_bh7_18_c4 <= tmp_bitheapResult_bh7_18_c3;
            end if;
            if ce_5 = '1' then
               tmp_bitheapResult_bh7_18_c5 <= tmp_bitheapResult_bh7_18_c4;
            end if;
            if ce_6 = '1' then
               tmp_bitheapResult_bh7_18_c6 <= tmp_bitheapResult_bh7_18_c5;
            end if;
            if ce_7 = '1' then
               tmp_bitheapResult_bh7_18_c7 <= tmp_bitheapResult_bh7_18_c6;
            end if;
            if ce_8 = '1' then
               tmp_bitheapResult_bh7_18_c8 <= tmp_bitheapResult_bh7_18_c7;
            end if;
            if ce_9 = '1' then
               tmp_bitheapResult_bh7_18_c9 <= tmp_bitheapResult_bh7_18_c8;
            end if;
            if ce_10 = '1' then
               tmp_bitheapResult_bh7_18_c10 <= tmp_bitheapResult_bh7_18_c9;
            end if;
            if ce_11 = '1' then
               tmp_bitheapResult_bh7_18_c11 <= tmp_bitheapResult_bh7_18_c10;
            end if;
            if ce_12 = '1' then
               tmp_bitheapResult_bh7_18_c12 <= tmp_bitheapResult_bh7_18_c11;
            end if;
            if ce_13 = '1' then
               tmp_bitheapResult_bh7_18_c13 <= tmp_bitheapResult_bh7_18_c12;
            end if;
         end if;
      end process;
   XX_m6_c0 <= X ;
   YY_m6_c0 <= Y ;
   tile_0_X_c0 <= X(16 downto 0);
   tile_0_Y_c0 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq800_uid9
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_0_X_c0,
                 Y => tile_0_Y_c0,
                 R => tile_0_output_c2);

   tile_0_filtered_output_c2 <= unsigned(tile_0_output_c2(40 downto 0));
   bh7_w0_0_c2 <= tile_0_filtered_output_c2(0);
   bh7_w1_0_c2 <= tile_0_filtered_output_c2(1);
   bh7_w2_0_c2 <= tile_0_filtered_output_c2(2);
   bh7_w3_0_c2 <= tile_0_filtered_output_c2(3);
   bh7_w4_0_c2 <= tile_0_filtered_output_c2(4);
   bh7_w5_0_c2 <= tile_0_filtered_output_c2(5);
   bh7_w6_0_c2 <= tile_0_filtered_output_c2(6);
   bh7_w7_0_c2 <= tile_0_filtered_output_c2(7);
   bh7_w8_0_c2 <= tile_0_filtered_output_c2(8);
   bh7_w9_0_c2 <= tile_0_filtered_output_c2(9);
   bh7_w10_0_c2 <= tile_0_filtered_output_c2(10);
   bh7_w11_0_c2 <= tile_0_filtered_output_c2(11);
   bh7_w12_0_c2 <= tile_0_filtered_output_c2(12);
   bh7_w13_0_c2 <= tile_0_filtered_output_c2(13);
   bh7_w14_0_c2 <= tile_0_filtered_output_c2(14);
   bh7_w15_0_c2 <= tile_0_filtered_output_c2(15);
   bh7_w16_0_c2 <= tile_0_filtered_output_c2(16);
   bh7_w17_0_c2 <= tile_0_filtered_output_c2(17);
   bh7_w18_0_c2 <= tile_0_filtered_output_c2(18);
   bh7_w19_0_c2 <= tile_0_filtered_output_c2(19);
   bh7_w20_0_c2 <= tile_0_filtered_output_c2(20);
   bh7_w21_0_c2 <= tile_0_filtered_output_c2(21);
   bh7_w22_0_c2 <= tile_0_filtered_output_c2(22);
   bh7_w23_0_c2 <= tile_0_filtered_output_c2(23);
   bh7_w24_0_c2 <= tile_0_filtered_output_c2(24);
   bh7_w25_0_c2 <= tile_0_filtered_output_c2(25);
   bh7_w26_0_c2 <= tile_0_filtered_output_c2(26);
   bh7_w27_0_c2 <= tile_0_filtered_output_c2(27);
   bh7_w28_0_c2 <= tile_0_filtered_output_c2(28);
   bh7_w29_0_c2 <= tile_0_filtered_output_c2(29);
   bh7_w30_0_c2 <= tile_0_filtered_output_c2(30);
   bh7_w31_0_c2 <= tile_0_filtered_output_c2(31);
   bh7_w32_0_c2 <= tile_0_filtered_output_c2(32);
   bh7_w33_0_c2 <= tile_0_filtered_output_c2(33);
   bh7_w34_0_c2 <= tile_0_filtered_output_c2(34);
   bh7_w35_0_c2 <= tile_0_filtered_output_c2(35);
   bh7_w36_0_c2 <= tile_0_filtered_output_c2(36);
   bh7_w37_0_c2 <= tile_0_filtered_output_c2(37);
   bh7_w38_0_c2 <= tile_0_filtered_output_c2(38);
   bh7_w39_0_c2 <= tile_0_filtered_output_c2(39);
   bh7_w40_0_c2 <= tile_0_filtered_output_c2(40);
   tile_1_X_c0 <= X(23 downto 23);
   tile_1_Y_c0 <= Y(23 downto 22);
   tile_1_mult: IntMultiplierLUT_1x2_Freq800_uid11
      port map ( clk  => clk,
                 X => tile_1_X_c0,
                 Y => tile_1_Y_c0,
                 R => tile_1_output_c0);

   tile_1_filtered_output_c0 <= unsigned(tile_1_output_c0(1 downto 0));
   bh7_w45_0_c0 <= tile_1_filtered_output_c0(0);
   bh7_w46_0_c0 <= tile_1_filtered_output_c0(1);
   tile_2_X_c0 <= X(22 downto 20);
   tile_2_Y_c0 <= Y(23 downto 22);
   tile_2_mult: IntMultiplierLUT_3x2_Freq800_uid13
      port map ( clk  => clk,
                 X => tile_2_X_c0,
                 Y => tile_2_Y_c0,
                 R => tile_2_output_c0);

   tile_2_filtered_output_c0 <= unsigned(tile_2_output_c0(4 downto 0));
   bh7_w42_0_c0 <= tile_2_filtered_output_c0(0);
   bh7_w43_0_c0 <= tile_2_filtered_output_c0(1);
   bh7_w44_0_c0 <= tile_2_filtered_output_c0(2);
   bh7_w45_1_c0 <= tile_2_filtered_output_c0(3);
   bh7_w46_1_c0 <= tile_2_filtered_output_c0(4);
   tile_3_X_c0 <= X(19 downto 17);
   tile_3_Y_c0 <= Y(23 downto 22);
   tile_3_mult: IntMultiplierLUT_3x2_Freq800_uid18
      port map ( clk  => clk,
                 X => tile_3_X_c0,
                 Y => tile_3_Y_c0,
                 R => tile_3_output_c0);

   tile_3_filtered_output_c0 <= unsigned(tile_3_output_c0(4 downto 0));
   bh7_w39_1_c0 <= tile_3_filtered_output_c0(0);
   bh7_w40_1_c0 <= tile_3_filtered_output_c0(1);
   bh7_w41_0_c0 <= tile_3_filtered_output_c0(2);
   bh7_w42_1_c0 <= tile_3_filtered_output_c0(3);
   bh7_w43_1_c0 <= tile_3_filtered_output_c0(4);
   tile_4_X_c0 <= X(23 downto 23);
   tile_4_Y_c0 <= Y(21 downto 20);
   tile_4_mult: IntMultiplierLUT_1x2_Freq800_uid23
      port map ( clk  => clk,
                 X => tile_4_X_c0,
                 Y => tile_4_Y_c0,
                 R => tile_4_output_c0);

   tile_4_filtered_output_c0 <= unsigned(tile_4_output_c0(1 downto 0));
   bh7_w43_2_c0 <= tile_4_filtered_output_c0(0);
   bh7_w44_1_c0 <= tile_4_filtered_output_c0(1);
   tile_5_X_c0 <= X(22 downto 20);
   tile_5_Y_c0 <= Y(21 downto 20);
   tile_5_mult: IntMultiplierLUT_3x2_Freq800_uid25
      port map ( clk  => clk,
                 X => tile_5_X_c0,
                 Y => tile_5_Y_c0,
                 R => tile_5_output_c0);

   tile_5_filtered_output_c0 <= unsigned(tile_5_output_c0(4 downto 0));
   bh7_w40_2_c0 <= tile_5_filtered_output_c0(0);
   bh7_w41_1_c0 <= tile_5_filtered_output_c0(1);
   bh7_w42_2_c0 <= tile_5_filtered_output_c0(2);
   bh7_w43_3_c0 <= tile_5_filtered_output_c0(3);
   bh7_w44_2_c0 <= tile_5_filtered_output_c0(4);
   tile_6_X_c0 <= X(19 downto 17);
   tile_6_Y_c0 <= Y(21 downto 20);
   tile_6_mult: IntMultiplierLUT_3x2_Freq800_uid30
      port map ( clk  => clk,
                 X => tile_6_X_c0,
                 Y => tile_6_Y_c0,
                 R => tile_6_output_c0);

   tile_6_filtered_output_c0 <= unsigned(tile_6_output_c0(4 downto 0));
   bh7_w37_1_c0 <= tile_6_filtered_output_c0(0);
   bh7_w38_1_c0 <= tile_6_filtered_output_c0(1);
   bh7_w39_2_c0 <= tile_6_filtered_output_c0(2);
   bh7_w40_3_c0 <= tile_6_filtered_output_c0(3);
   bh7_w41_2_c0 <= tile_6_filtered_output_c0(4);
   tile_7_X_c0 <= X(23 downto 23);
   tile_7_Y_c0 <= Y(19 downto 18);
   tile_7_mult: IntMultiplierLUT_1x2_Freq800_uid35
      port map ( clk  => clk,
                 X => tile_7_X_c0,
                 Y => tile_7_Y_c0,
                 R => tile_7_output_c0);

   tile_7_filtered_output_c0 <= unsigned(tile_7_output_c0(1 downto 0));
   bh7_w41_3_c0 <= tile_7_filtered_output_c0(0);
   bh7_w42_3_c0 <= tile_7_filtered_output_c0(1);
   tile_8_X_c0 <= X(22 downto 20);
   tile_8_Y_c0 <= Y(19 downto 18);
   tile_8_mult: IntMultiplierLUT_3x2_Freq800_uid37
      port map ( clk  => clk,
                 X => tile_8_X_c0,
                 Y => tile_8_Y_c0,
                 R => tile_8_output_c0);

   tile_8_filtered_output_c0 <= unsigned(tile_8_output_c0(4 downto 0));
   bh7_w38_2_c0 <= tile_8_filtered_output_c0(0);
   bh7_w39_3_c0 <= tile_8_filtered_output_c0(1);
   bh7_w40_4_c0 <= tile_8_filtered_output_c0(2);
   bh7_w41_4_c0 <= tile_8_filtered_output_c0(3);
   bh7_w42_4_c0 <= tile_8_filtered_output_c0(4);
   tile_9_X_c0 <= X(19 downto 17);
   tile_9_Y_c0 <= Y(19 downto 18);
   tile_9_mult: IntMultiplierLUT_3x2_Freq800_uid42
      port map ( clk  => clk,
                 X => tile_9_X_c0,
                 Y => tile_9_Y_c0,
                 R => tile_9_output_c0);

   tile_9_filtered_output_c0 <= unsigned(tile_9_output_c0(4 downto 0));
   bh7_w35_1_c0 <= tile_9_filtered_output_c0(0);
   bh7_w36_1_c0 <= tile_9_filtered_output_c0(1);
   bh7_w37_2_c0 <= tile_9_filtered_output_c0(2);
   bh7_w38_3_c0 <= tile_9_filtered_output_c0(3);
   bh7_w39_4_c0 <= tile_9_filtered_output_c0(4);
   tile_10_X_c0 <= X(23 downto 23);
   tile_10_Y_c0 <= Y(17 downto 16);
   tile_10_mult: IntMultiplierLUT_1x2_Freq800_uid47
      port map ( clk  => clk,
                 X => tile_10_X_c0,
                 Y => tile_10_Y_c0,
                 R => tile_10_output_c0);

   tile_10_filtered_output_c0 <= unsigned(tile_10_output_c0(1 downto 0));
   bh7_w39_5_c0 <= tile_10_filtered_output_c0(0);
   bh7_w40_5_c0 <= tile_10_filtered_output_c0(1);
   tile_11_X_c0 <= X(22 downto 20);
   tile_11_Y_c0 <= Y(17 downto 16);
   tile_11_mult: IntMultiplierLUT_3x2_Freq800_uid49
      port map ( clk  => clk,
                 X => tile_11_X_c0,
                 Y => tile_11_Y_c0,
                 R => tile_11_output_c0);

   tile_11_filtered_output_c0 <= unsigned(tile_11_output_c0(4 downto 0));
   bh7_w36_2_c0 <= tile_11_filtered_output_c0(0);
   bh7_w37_3_c0 <= tile_11_filtered_output_c0(1);
   bh7_w38_4_c0 <= tile_11_filtered_output_c0(2);
   bh7_w39_6_c0 <= tile_11_filtered_output_c0(3);
   bh7_w40_6_c0 <= tile_11_filtered_output_c0(4);
   tile_12_X_c0 <= X(19 downto 17);
   tile_12_Y_c0 <= Y(17 downto 16);
   tile_12_mult: IntMultiplierLUT_3x2_Freq800_uid54
      port map ( clk  => clk,
                 X => tile_12_X_c0,
                 Y => tile_12_Y_c0,
                 R => tile_12_output_c0);

   tile_12_filtered_output_c0 <= unsigned(tile_12_output_c0(4 downto 0));
   bh7_w33_1_c0 <= tile_12_filtered_output_c0(0);
   bh7_w34_1_c0 <= tile_12_filtered_output_c0(1);
   bh7_w35_2_c0 <= tile_12_filtered_output_c0(2);
   bh7_w36_3_c0 <= tile_12_filtered_output_c0(3);
   bh7_w37_4_c0 <= tile_12_filtered_output_c0(4);
   tile_13_X_c0 <= X(23 downto 23);
   tile_13_Y_c0 <= Y(15 downto 14);
   tile_13_mult: IntMultiplierLUT_1x2_Freq800_uid59
      port map ( clk  => clk,
                 X => tile_13_X_c0,
                 Y => tile_13_Y_c0,
                 R => tile_13_output_c0);

   tile_13_filtered_output_c0 <= unsigned(tile_13_output_c0(1 downto 0));
   bh7_w37_5_c0 <= tile_13_filtered_output_c0(0);
   bh7_w38_5_c0 <= tile_13_filtered_output_c0(1);
   tile_14_X_c0 <= X(22 downto 20);
   tile_14_Y_c0 <= Y(15 downto 14);
   tile_14_mult: IntMultiplierLUT_3x2_Freq800_uid61
      port map ( clk  => clk,
                 X => tile_14_X_c0,
                 Y => tile_14_Y_c0,
                 R => tile_14_output_c0);

   tile_14_filtered_output_c0 <= unsigned(tile_14_output_c0(4 downto 0));
   bh7_w34_2_c0 <= tile_14_filtered_output_c0(0);
   bh7_w35_3_c0 <= tile_14_filtered_output_c0(1);
   bh7_w36_4_c0 <= tile_14_filtered_output_c0(2);
   bh7_w37_6_c0 <= tile_14_filtered_output_c0(3);
   bh7_w38_6_c0 <= tile_14_filtered_output_c0(4);
   tile_15_X_c0 <= X(19 downto 17);
   tile_15_Y_c0 <= Y(15 downto 14);
   tile_15_mult: IntMultiplierLUT_3x2_Freq800_uid66
      port map ( clk  => clk,
                 X => tile_15_X_c0,
                 Y => tile_15_Y_c0,
                 R => tile_15_output_c0);

   tile_15_filtered_output_c0 <= unsigned(tile_15_output_c0(4 downto 0));
   bh7_w31_1_c0 <= tile_15_filtered_output_c0(0);
   bh7_w32_1_c0 <= tile_15_filtered_output_c0(1);
   bh7_w33_2_c0 <= tile_15_filtered_output_c0(2);
   bh7_w34_3_c0 <= tile_15_filtered_output_c0(3);
   bh7_w35_4_c0 <= tile_15_filtered_output_c0(4);
   tile_16_X_c0 <= X(23 downto 23);
   tile_16_Y_c0 <= Y(13 downto 12);
   tile_16_mult: IntMultiplierLUT_1x2_Freq800_uid71
      port map ( clk  => clk,
                 X => tile_16_X_c0,
                 Y => tile_16_Y_c0,
                 R => tile_16_output_c0);

   tile_16_filtered_output_c0 <= unsigned(tile_16_output_c0(1 downto 0));
   bh7_w35_5_c0 <= tile_16_filtered_output_c0(0);
   bh7_w36_5_c0 <= tile_16_filtered_output_c0(1);
   tile_17_X_c0 <= X(22 downto 20);
   tile_17_Y_c0 <= Y(13 downto 12);
   tile_17_mult: IntMultiplierLUT_3x2_Freq800_uid73
      port map ( clk  => clk,
                 X => tile_17_X_c0,
                 Y => tile_17_Y_c0,
                 R => tile_17_output_c0);

   tile_17_filtered_output_c0 <= unsigned(tile_17_output_c0(4 downto 0));
   bh7_w32_2_c0 <= tile_17_filtered_output_c0(0);
   bh7_w33_3_c0 <= tile_17_filtered_output_c0(1);
   bh7_w34_4_c0 <= tile_17_filtered_output_c0(2);
   bh7_w35_6_c0 <= tile_17_filtered_output_c0(3);
   bh7_w36_6_c0 <= tile_17_filtered_output_c0(4);
   tile_18_X_c0 <= X(19 downto 17);
   tile_18_Y_c0 <= Y(13 downto 12);
   tile_18_mult: IntMultiplierLUT_3x2_Freq800_uid78
      port map ( clk  => clk,
                 X => tile_18_X_c0,
                 Y => tile_18_Y_c0,
                 R => tile_18_output_c0);

   tile_18_filtered_output_c0 <= unsigned(tile_18_output_c0(4 downto 0));
   bh7_w29_1_c0 <= tile_18_filtered_output_c0(0);
   bh7_w30_1_c0 <= tile_18_filtered_output_c0(1);
   bh7_w31_2_c0 <= tile_18_filtered_output_c0(2);
   bh7_w32_3_c0 <= tile_18_filtered_output_c0(3);
   bh7_w33_4_c0 <= tile_18_filtered_output_c0(4);
   tile_19_X_c0 <= X(23 downto 23);
   tile_19_Y_c0 <= Y(11 downto 10);
   tile_19_mult: IntMultiplierLUT_1x2_Freq800_uid83
      port map ( clk  => clk,
                 X => tile_19_X_c0,
                 Y => tile_19_Y_c0,
                 R => tile_19_output_c0);

   tile_19_filtered_output_c0 <= unsigned(tile_19_output_c0(1 downto 0));
   bh7_w33_5_c0 <= tile_19_filtered_output_c0(0);
   bh7_w34_5_c0 <= tile_19_filtered_output_c0(1);
   tile_20_X_c0 <= X(22 downto 20);
   tile_20_Y_c0 <= Y(11 downto 10);
   tile_20_mult: IntMultiplierLUT_3x2_Freq800_uid85
      port map ( clk  => clk,
                 X => tile_20_X_c0,
                 Y => tile_20_Y_c0,
                 R => tile_20_output_c0);

   tile_20_filtered_output_c0 <= unsigned(tile_20_output_c0(4 downto 0));
   bh7_w30_2_c0 <= tile_20_filtered_output_c0(0);
   bh7_w31_3_c0 <= tile_20_filtered_output_c0(1);
   bh7_w32_4_c0 <= tile_20_filtered_output_c0(2);
   bh7_w33_6_c0 <= tile_20_filtered_output_c0(3);
   bh7_w34_6_c0 <= tile_20_filtered_output_c0(4);
   tile_21_X_c0 <= X(19 downto 17);
   tile_21_Y_c0 <= Y(11 downto 10);
   tile_21_mult: IntMultiplierLUT_3x2_Freq800_uid90
      port map ( clk  => clk,
                 X => tile_21_X_c0,
                 Y => tile_21_Y_c0,
                 R => tile_21_output_c0);

   tile_21_filtered_output_c0 <= unsigned(tile_21_output_c0(4 downto 0));
   bh7_w27_1_c0 <= tile_21_filtered_output_c0(0);
   bh7_w28_1_c0 <= tile_21_filtered_output_c0(1);
   bh7_w29_2_c0 <= tile_21_filtered_output_c0(2);
   bh7_w30_3_c0 <= tile_21_filtered_output_c0(3);
   bh7_w31_4_c0 <= tile_21_filtered_output_c0(4);
   tile_22_X_c0 <= X(23 downto 23);
   tile_22_Y_c0 <= Y(9 downto 8);
   tile_22_mult: IntMultiplierLUT_1x2_Freq800_uid95
      port map ( clk  => clk,
                 X => tile_22_X_c0,
                 Y => tile_22_Y_c0,
                 R => tile_22_output_c0);

   tile_22_filtered_output_c0 <= unsigned(tile_22_output_c0(1 downto 0));
   bh7_w31_5_c0 <= tile_22_filtered_output_c0(0);
   bh7_w32_5_c0 <= tile_22_filtered_output_c0(1);
   tile_23_X_c0 <= X(22 downto 20);
   tile_23_Y_c0 <= Y(9 downto 8);
   tile_23_mult: IntMultiplierLUT_3x2_Freq800_uid97
      port map ( clk  => clk,
                 X => tile_23_X_c0,
                 Y => tile_23_Y_c0,
                 R => tile_23_output_c0);

   tile_23_filtered_output_c0 <= unsigned(tile_23_output_c0(4 downto 0));
   bh7_w28_2_c0 <= tile_23_filtered_output_c0(0);
   bh7_w29_3_c0 <= tile_23_filtered_output_c0(1);
   bh7_w30_4_c0 <= tile_23_filtered_output_c0(2);
   bh7_w31_6_c0 <= tile_23_filtered_output_c0(3);
   bh7_w32_6_c0 <= tile_23_filtered_output_c0(4);
   tile_24_X_c0 <= X(19 downto 17);
   tile_24_Y_c0 <= Y(9 downto 8);
   tile_24_mult: IntMultiplierLUT_3x2_Freq800_uid102
      port map ( clk  => clk,
                 X => tile_24_X_c0,
                 Y => tile_24_Y_c0,
                 R => tile_24_output_c0);

   tile_24_filtered_output_c0 <= unsigned(tile_24_output_c0(4 downto 0));
   bh7_w25_1_c0 <= tile_24_filtered_output_c0(0);
   bh7_w26_1_c0 <= tile_24_filtered_output_c0(1);
   bh7_w27_2_c0 <= tile_24_filtered_output_c0(2);
   bh7_w28_3_c0 <= tile_24_filtered_output_c0(3);
   bh7_w29_4_c0 <= tile_24_filtered_output_c0(4);
   tile_25_X_c0 <= X(23 downto 23);
   tile_25_Y_c0 <= Y(7 downto 6);
   tile_25_mult: IntMultiplierLUT_1x2_Freq800_uid107
      port map ( clk  => clk,
                 X => tile_25_X_c0,
                 Y => tile_25_Y_c0,
                 R => tile_25_output_c0);

   tile_25_filtered_output_c0 <= unsigned(tile_25_output_c0(1 downto 0));
   bh7_w29_5_c0 <= tile_25_filtered_output_c0(0);
   bh7_w30_5_c0 <= tile_25_filtered_output_c0(1);
   tile_26_X_c0 <= X(22 downto 20);
   tile_26_Y_c0 <= Y(7 downto 6);
   tile_26_mult: IntMultiplierLUT_3x2_Freq800_uid109
      port map ( clk  => clk,
                 X => tile_26_X_c0,
                 Y => tile_26_Y_c0,
                 R => tile_26_output_c0);

   tile_26_filtered_output_c0 <= unsigned(tile_26_output_c0(4 downto 0));
   bh7_w26_2_c0 <= tile_26_filtered_output_c0(0);
   bh7_w27_3_c0 <= tile_26_filtered_output_c0(1);
   bh7_w28_4_c0 <= tile_26_filtered_output_c0(2);
   bh7_w29_6_c0 <= tile_26_filtered_output_c0(3);
   bh7_w30_6_c0 <= tile_26_filtered_output_c0(4);
   tile_27_X_c0 <= X(19 downto 17);
   tile_27_Y_c0 <= Y(7 downto 6);
   tile_27_mult: IntMultiplierLUT_3x2_Freq800_uid114
      port map ( clk  => clk,
                 X => tile_27_X_c0,
                 Y => tile_27_Y_c0,
                 R => tile_27_output_c0);

   tile_27_filtered_output_c0 <= unsigned(tile_27_output_c0(4 downto 0));
   bh7_w23_1_c0 <= tile_27_filtered_output_c0(0);
   bh7_w24_1_c0 <= tile_27_filtered_output_c0(1);
   bh7_w25_2_c0 <= tile_27_filtered_output_c0(2);
   bh7_w26_3_c0 <= tile_27_filtered_output_c0(3);
   bh7_w27_4_c0 <= tile_27_filtered_output_c0(4);
   tile_28_X_c0 <= X(23 downto 23);
   tile_28_Y_c0 <= Y(5 downto 4);
   tile_28_mult: IntMultiplierLUT_1x2_Freq800_uid119
      port map ( clk  => clk,
                 X => tile_28_X_c0,
                 Y => tile_28_Y_c0,
                 R => tile_28_output_c0);

   tile_28_filtered_output_c0 <= unsigned(tile_28_output_c0(1 downto 0));
   bh7_w27_5_c0 <= tile_28_filtered_output_c0(0);
   bh7_w28_5_c0 <= tile_28_filtered_output_c0(1);
   tile_29_X_c0 <= X(22 downto 20);
   tile_29_Y_c0 <= Y(5 downto 4);
   tile_29_mult: IntMultiplierLUT_3x2_Freq800_uid121
      port map ( clk  => clk,
                 X => tile_29_X_c0,
                 Y => tile_29_Y_c0,
                 R => tile_29_output_c0);

   tile_29_filtered_output_c0 <= unsigned(tile_29_output_c0(4 downto 0));
   bh7_w24_2_c0 <= tile_29_filtered_output_c0(0);
   bh7_w25_3_c0 <= tile_29_filtered_output_c0(1);
   bh7_w26_4_c0 <= tile_29_filtered_output_c0(2);
   bh7_w27_6_c0 <= tile_29_filtered_output_c0(3);
   bh7_w28_6_c0 <= tile_29_filtered_output_c0(4);
   tile_30_X_c0 <= X(19 downto 17);
   tile_30_Y_c0 <= Y(5 downto 4);
   tile_30_mult: IntMultiplierLUT_3x2_Freq800_uid126
      port map ( clk  => clk,
                 X => tile_30_X_c0,
                 Y => tile_30_Y_c0,
                 R => tile_30_output_c0);

   tile_30_filtered_output_c0 <= unsigned(tile_30_output_c0(4 downto 0));
   bh7_w21_1_c0 <= tile_30_filtered_output_c0(0);
   bh7_w22_1_c0 <= tile_30_filtered_output_c0(1);
   bh7_w23_2_c0 <= tile_30_filtered_output_c0(2);
   bh7_w24_3_c0 <= tile_30_filtered_output_c0(3);
   bh7_w25_4_c0 <= tile_30_filtered_output_c0(4);
   tile_31_X_c0 <= X(23 downto 23);
   tile_31_Y_c0 <= Y(3 downto 2);
   tile_31_mult: IntMultiplierLUT_1x2_Freq800_uid131
      port map ( clk  => clk,
                 X => tile_31_X_c0,
                 Y => tile_31_Y_c0,
                 R => tile_31_output_c0);

   tile_31_filtered_output_c0 <= unsigned(tile_31_output_c0(1 downto 0));
   bh7_w25_5_c0 <= tile_31_filtered_output_c0(0);
   bh7_w26_5_c0 <= tile_31_filtered_output_c0(1);
   tile_32_X_c0 <= X(22 downto 20);
   tile_32_Y_c0 <= Y(3 downto 2);
   tile_32_mult: IntMultiplierLUT_3x2_Freq800_uid133
      port map ( clk  => clk,
                 X => tile_32_X_c0,
                 Y => tile_32_Y_c0,
                 R => tile_32_output_c0);

   tile_32_filtered_output_c0 <= unsigned(tile_32_output_c0(4 downto 0));
   bh7_w22_2_c0 <= tile_32_filtered_output_c0(0);
   bh7_w23_3_c0 <= tile_32_filtered_output_c0(1);
   bh7_w24_4_c0 <= tile_32_filtered_output_c0(2);
   bh7_w25_6_c0 <= tile_32_filtered_output_c0(3);
   bh7_w26_6_c0 <= tile_32_filtered_output_c0(4);
   tile_33_X_c0 <= X(19 downto 17);
   tile_33_Y_c0 <= Y(3 downto 2);
   tile_33_mult: IntMultiplierLUT_3x2_Freq800_uid138
      port map ( clk  => clk,
                 X => tile_33_X_c0,
                 Y => tile_33_Y_c0,
                 R => tile_33_output_c0);

   tile_33_filtered_output_c0 <= unsigned(tile_33_output_c0(4 downto 0));
   bh7_w19_1_c0 <= tile_33_filtered_output_c0(0);
   bh7_w20_1_c0 <= tile_33_filtered_output_c0(1);
   bh7_w21_2_c0 <= tile_33_filtered_output_c0(2);
   bh7_w22_3_c0 <= tile_33_filtered_output_c0(3);
   bh7_w23_4_c0 <= tile_33_filtered_output_c0(4);
   tile_34_X_c0 <= X(23 downto 23);
   tile_34_Y_c0 <= Y(1 downto 0);
   tile_34_mult: IntMultiplierLUT_1x2_Freq800_uid143
      port map ( clk  => clk,
                 X => tile_34_X_c0,
                 Y => tile_34_Y_c0,
                 R => tile_34_output_c0);

   tile_34_filtered_output_c0 <= unsigned(tile_34_output_c0(1 downto 0));
   bh7_w23_5_c0 <= tile_34_filtered_output_c0(0);
   bh7_w24_5_c0 <= tile_34_filtered_output_c0(1);
   tile_35_X_c0 <= X(22 downto 20);
   tile_35_Y_c0 <= Y(1 downto 0);
   tile_35_mult: IntMultiplierLUT_3x2_Freq800_uid145
      port map ( clk  => clk,
                 X => tile_35_X_c0,
                 Y => tile_35_Y_c0,
                 R => tile_35_output_c0);

   tile_35_filtered_output_c0 <= unsigned(tile_35_output_c0(4 downto 0));
   bh7_w20_2_c0 <= tile_35_filtered_output_c0(0);
   bh7_w21_3_c0 <= tile_35_filtered_output_c0(1);
   bh7_w22_4_c0 <= tile_35_filtered_output_c0(2);
   bh7_w23_6_c0 <= tile_35_filtered_output_c0(3);
   bh7_w24_6_c0 <= tile_35_filtered_output_c0(4);
   tile_36_X_c0 <= X(19 downto 17);
   tile_36_Y_c0 <= Y(1 downto 0);
   tile_36_mult: IntMultiplierLUT_3x2_Freq800_uid150
      port map ( clk  => clk,
                 X => tile_36_X_c0,
                 Y => tile_36_Y_c0,
                 R => tile_36_output_c0);

   tile_36_filtered_output_c0 <= unsigned(tile_36_output_c0(4 downto 0));
   bh7_w17_1_c0 <= tile_36_filtered_output_c0(0);
   bh7_w18_1_c0 <= tile_36_filtered_output_c0(1);
   bh7_w19_2_c0 <= tile_36_filtered_output_c0(2);
   bh7_w20_3_c0 <= tile_36_filtered_output_c0(3);
   bh7_w21_4_c0 <= tile_36_filtered_output_c0(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq800_uid156_bh7_uid157_In0_c0 <= "" & bh7_w18_1_c0 & "0" & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid157_In1_c0 <= "" & bh7_w19_1_c0 & bh7_w19_2_c0;
   bh7_w18_2_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_c1(0);
   bh7_w19_3_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_c1(1);
   bh7_w20_4_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid157: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid157_In0_c0,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid157_In1_c0,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_copy158_c0);
   Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid157_Out0_copy158_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid160_bh7_uid161_In0_c0 <= "" & bh7_w20_1_c0 & bh7_w20_2_c0 & bh7_w20_3_c0;
   bh7_w20_5_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_c1(0);
   bh7_w21_5_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_c1(1);
   Compressor_3_2_Freq800_uid160_uid161: Compressor_3_2_Freq800_uid160
      port map ( X0 => Compressor_3_2_Freq800_uid160_bh7_uid161_In0_c0,
                 R => Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_copy162_c0);
   Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid161_Out0_copy162_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid165_In0_c0 <= "" & bh7_w21_1_c0 & bh7_w21_2_c0 & bh7_w21_3_c0 & bh7_w21_4_c0;
   Compressor_14_3_Freq800_uid164_bh7_uid165_In1_c0 <= "" & bh7_w22_1_c0;
   bh7_w21_6_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_c1(0);
   bh7_w22_5_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_c1(1);
   bh7_w23_7_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_c1(2);
   Compressor_14_3_Freq800_uid164_uid165: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid165_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid165_In1_c0,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_copy166_c0);
   Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid165_Out0_copy166_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid160_bh7_uid167_In0_c0 <= "" & bh7_w22_2_c0 & bh7_w22_3_c0 & bh7_w22_4_c0;
   bh7_w22_6_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_c1(0);
   bh7_w23_8_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_c1(1);
   Compressor_3_2_Freq800_uid160_uid167: Compressor_3_2_Freq800_uid160
      port map ( X0 => Compressor_3_2_Freq800_uid160_bh7_uid167_In0_c0,
                 R => Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_copy168_c0);
   Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid167_Out0_copy168_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid171_In0_c0 <= "" & bh7_w23_1_c0 & bh7_w23_2_c0 & bh7_w23_3_c0 & bh7_w23_4_c0 & bh7_w23_5_c0 & bh7_w23_6_c0;
   bh7_w23_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_c1(0);
   bh7_w24_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_c1(1);
   bh7_w25_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid171: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid171_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_copy172_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid171_Out0_copy172_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid173_In0_c0 <= "" & bh7_w24_1_c0 & bh7_w24_2_c0 & bh7_w24_3_c0 & bh7_w24_4_c0 & bh7_w24_5_c0 & bh7_w24_6_c0;
   bh7_w24_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_c1(0);
   bh7_w25_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_c1(1);
   bh7_w26_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid173: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid173_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_copy174_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid173_Out0_copy174_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid175_In0_c0 <= "" & bh7_w25_1_c0 & bh7_w25_2_c0 & bh7_w25_3_c0 & bh7_w25_4_c0 & bh7_w25_5_c0 & bh7_w25_6_c0;
   bh7_w25_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_c1(0);
   bh7_w26_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_c1(1);
   bh7_w27_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid175: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid175_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_copy176_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid175_Out0_copy176_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid177_In0_c0 <= "" & bh7_w26_1_c0 & bh7_w26_2_c0 & bh7_w26_3_c0 & bh7_w26_4_c0 & bh7_w26_5_c0 & bh7_w26_6_c0;
   bh7_w26_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_c1(0);
   bh7_w27_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_c1(1);
   bh7_w28_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid177: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid177_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_copy178_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid177_Out0_copy178_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid179_In0_c0 <= "" & bh7_w27_1_c0 & bh7_w27_2_c0 & bh7_w27_3_c0 & bh7_w27_4_c0 & bh7_w27_5_c0 & bh7_w27_6_c0;
   bh7_w27_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_c1(0);
   bh7_w28_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_c1(1);
   bh7_w29_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid179: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid179_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_copy180_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid179_Out0_copy180_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid181_In0_c0 <= "" & bh7_w28_1_c0 & bh7_w28_2_c0 & bh7_w28_3_c0 & bh7_w28_4_c0 & bh7_w28_5_c0 & bh7_w28_6_c0;
   bh7_w28_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_c1(0);
   bh7_w29_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_c1(1);
   bh7_w30_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid181: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid181_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_copy182_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid181_Out0_copy182_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid183_In0_c0 <= "" & bh7_w29_1_c0 & bh7_w29_2_c0 & bh7_w29_3_c0 & bh7_w29_4_c0 & bh7_w29_5_c0 & bh7_w29_6_c0;
   bh7_w29_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_c1(0);
   bh7_w30_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_c1(1);
   bh7_w31_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid183: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid183_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_copy184_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid183_Out0_copy184_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid185_In0_c0 <= "" & bh7_w30_1_c0 & bh7_w30_2_c0 & bh7_w30_3_c0 & bh7_w30_4_c0 & bh7_w30_5_c0 & bh7_w30_6_c0;
   bh7_w30_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_c1(0);
   bh7_w31_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_c1(1);
   bh7_w32_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid185: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid185_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_copy186_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid185_Out0_copy186_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid187_In0_c0 <= "" & bh7_w31_1_c0 & bh7_w31_2_c0 & bh7_w31_3_c0 & bh7_w31_4_c0 & bh7_w31_5_c0 & bh7_w31_6_c0;
   bh7_w31_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_c1(0);
   bh7_w32_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_c1(1);
   bh7_w33_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid187: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid187_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_copy188_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid187_Out0_copy188_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid189_In0_c0 <= "" & bh7_w32_1_c0 & bh7_w32_2_c0 & bh7_w32_3_c0 & bh7_w32_4_c0 & bh7_w32_5_c0 & bh7_w32_6_c0;
   bh7_w32_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_c1(0);
   bh7_w33_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_c1(1);
   bh7_w34_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid189: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid189_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_copy190_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid189_Out0_copy190_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid191_In0_c0 <= "" & bh7_w33_1_c0 & bh7_w33_2_c0 & bh7_w33_3_c0 & bh7_w33_4_c0 & bh7_w33_5_c0 & bh7_w33_6_c0;
   bh7_w33_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_c1(0);
   bh7_w34_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_c1(1);
   bh7_w35_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid191: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid191_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_copy192_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid191_Out0_copy192_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid193_In0_c0 <= "" & bh7_w34_1_c0 & bh7_w34_2_c0 & bh7_w34_3_c0 & bh7_w34_4_c0 & bh7_w34_5_c0 & bh7_w34_6_c0;
   bh7_w34_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_c1(0);
   bh7_w35_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_c1(1);
   bh7_w36_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid193: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid193_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_copy194_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid193_Out0_copy194_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid195_In0_c0 <= "" & bh7_w35_1_c0 & bh7_w35_2_c0 & bh7_w35_3_c0 & bh7_w35_4_c0 & bh7_w35_5_c0 & bh7_w35_6_c0;
   bh7_w35_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_c1(0);
   bh7_w36_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_c1(1);
   bh7_w37_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid195: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid195_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_copy196_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid195_Out0_copy196_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid197_In0_c0 <= "" & bh7_w36_1_c0 & bh7_w36_2_c0 & bh7_w36_3_c0 & bh7_w36_4_c0 & bh7_w36_5_c0 & bh7_w36_6_c0;
   bh7_w36_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_c1(0);
   bh7_w37_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_c1(1);
   bh7_w38_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid197: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid197_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_copy198_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid197_Out0_copy198_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid199_In0_c0 <= "" & bh7_w37_1_c0 & bh7_w37_2_c0 & bh7_w37_3_c0 & bh7_w37_4_c0 & bh7_w37_5_c0 & bh7_w37_6_c0;
   bh7_w37_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_c1(0);
   bh7_w38_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_c1(1);
   bh7_w39_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid199: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid199_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_copy200_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid199_Out0_copy200_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid201_In0_c0 <= "" & bh7_w38_1_c0 & bh7_w38_2_c0 & bh7_w38_3_c0 & bh7_w38_4_c0 & bh7_w38_5_c0 & bh7_w38_6_c0;
   bh7_w38_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_c1(0);
   bh7_w39_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_c1(1);
   bh7_w40_7_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid201: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid201_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_copy202_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid201_Out0_copy202_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid203_In0_c0 <= "" & bh7_w39_1_c0 & bh7_w39_2_c0 & bh7_w39_3_c0 & bh7_w39_4_c0 & bh7_w39_5_c0 & bh7_w39_6_c0;
   bh7_w39_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_c1(0);
   bh7_w40_8_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_c1(1);
   bh7_w41_5_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid203: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid203_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_copy204_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid203_Out0_copy204_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid170_bh7_uid205_In0_c0 <= "" & bh7_w40_1_c0 & bh7_w40_2_c0 & bh7_w40_3_c0 & bh7_w40_4_c0 & bh7_w40_5_c0 & bh7_w40_6_c0;
   bh7_w40_9_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_c1(0);
   bh7_w41_6_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_c1(1);
   bh7_w42_5_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_c1(2);
   Compressor_6_3_Freq800_uid170_uid205: Compressor_6_3_Freq800_uid170
      port map ( X0 => Compressor_6_3_Freq800_uid170_bh7_uid205_In0_c0,
                 R => Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_copy206_c0);
   Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_c1 <= Compressor_6_3_Freq800_uid170_bh7_uid205_Out0_copy206_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid207_In0_c0 <= "" & bh7_w41_0_c0 & bh7_w41_1_c0 & bh7_w41_2_c0 & bh7_w41_3_c0;
   Compressor_14_3_Freq800_uid164_bh7_uid207_In1_c0 <= "" & bh7_w42_0_c0;
   bh7_w41_7_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_c1(0);
   bh7_w42_6_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_c1(1);
   bh7_w43_4_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_c1(2);
   Compressor_14_3_Freq800_uid164_uid207: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid207_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid207_In1_c0,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_copy208_c0);
   Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid207_Out0_copy208_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid209_In0_c0 <= "" & bh7_w42_1_c0 & bh7_w42_2_c0 & bh7_w42_3_c0 & bh7_w42_4_c0;
   Compressor_14_3_Freq800_uid164_bh7_uid209_In1_c0 <= "" & bh7_w43_0_c0;
   bh7_w42_7_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_c1(0);
   bh7_w43_5_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_c1(1);
   bh7_w44_3_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_c1(2);
   Compressor_14_3_Freq800_uid164_uid209: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid209_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid209_In1_c0,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_copy210_c0);
   Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid209_Out0_copy210_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid211_In0_c0 <= "" & bh7_w43_1_c0 & bh7_w43_2_c0 & bh7_w43_3_c0;
   Compressor_23_3_Freq800_uid156_bh7_uid211_In1_c0 <= "" & bh7_w44_0_c0 & bh7_w44_1_c0;
   bh7_w43_6_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_c1(0);
   bh7_w44_4_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_c1(1);
   bh7_w45_2_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid211: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid211_In0_c0,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid211_In1_c0,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_copy212_c0);
   Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid211_Out0_copy212_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid213_In0_c0 <= "" & bh7_w45_0_c0 & bh7_w45_1_c0 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid213_In1_c0 <= "" & bh7_w46_0_c0 & bh7_w46_1_c0;
   bh7_w45_3_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_c1(0);
   bh7_w46_2_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_c1(1);
   bh7_w47_0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid213: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid213_In0_c0,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid213_In1_c0,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_copy214_c0);
   Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid213_Out0_copy214_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid215_In0_c1 <= "" & bh7_w20_5_c1 & bh7_w20_4_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid215_In1_c1 <= "" & bh7_w21_6_c1 & bh7_w21_5_c1;
   bh7_w20_6_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid215_Out0_c1(0);
   bh7_w21_7_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid215_Out0_c1(1);
   bh7_w22_7_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid215_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid215: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid215_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid215_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid215_Out0_copy216_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid215_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid215_Out0_copy216_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid160_bh7_uid217_In0_c1 <= "" & bh7_w22_6_c1 & bh7_w22_5_c1 & "0";
   bh7_w22_8_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid217_Out0_c1(0);
   bh7_w23_10_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid217_Out0_c1(1);
   Compressor_3_2_Freq800_uid160_uid217: Compressor_3_2_Freq800_uid160
      port map ( X0 => Compressor_3_2_Freq800_uid160_bh7_uid217_In0_c1,
                 R => Compressor_3_2_Freq800_uid160_bh7_uid217_Out0_copy218_c1);
   Compressor_3_2_Freq800_uid160_bh7_uid217_Out0_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid217_Out0_copy218_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid219_In0_c1 <= "" & bh7_w23_8_c1 & bh7_w23_7_c1 & bh7_w23_9_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid219_In1_c1 <= "" & bh7_w24_8_c1 & bh7_w24_7_c1;
   bh7_w23_11_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid219_Out0_c1(0);
   bh7_w24_9_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid219_Out0_c1(1);
   bh7_w25_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid219_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid219: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid219_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid219_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid219_Out0_copy220_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid219_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid219_Out0_copy220_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid221_In0_c1 <= "" & bh7_w25_9_c1 & bh7_w25_8_c1 & bh7_w25_7_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid221_In1_c1 <= "" & bh7_w26_9_c1 & bh7_w26_8_c1;
   bh7_w25_11_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid221_Out0_c1(0);
   bh7_w26_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid221_Out0_c1(1);
   bh7_w27_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid221_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid221: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid221_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid221_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid221_Out0_copy222_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid221_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid221_Out0_copy222_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid223_In0_c1 <= "" & bh7_w27_9_c1 & bh7_w27_8_c1 & bh7_w27_7_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid223_In1_c1 <= "" & bh7_w28_9_c1 & bh7_w28_8_c1;
   bh7_w27_11_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid223_Out0_c1(0);
   bh7_w28_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid223_Out0_c1(1);
   bh7_w29_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid223_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid223: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid223_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid223_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid223_Out0_copy224_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid223_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid223_Out0_copy224_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid225_In0_c1 <= "" & bh7_w29_9_c1 & bh7_w29_8_c1 & bh7_w29_7_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid225_In1_c1 <= "" & bh7_w30_9_c1 & bh7_w30_8_c1;
   bh7_w29_11_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid225_Out0_c1(0);
   bh7_w30_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid225_Out0_c1(1);
   bh7_w31_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid225_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid225: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid225_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid225_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid225_Out0_copy226_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid225_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid225_Out0_copy226_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid227_In0_c1 <= "" & bh7_w31_9_c1 & bh7_w31_8_c1 & bh7_w31_7_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid227_In1_c1 <= "" & bh7_w32_9_c1 & bh7_w32_8_c1;
   bh7_w31_11_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid227_Out0_c1(0);
   bh7_w32_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid227_Out0_c1(1);
   bh7_w33_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid227_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid227: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid227_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid227_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid227_Out0_copy228_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid227_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid227_Out0_copy228_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid229_In0_c1 <= "" & bh7_w33_9_c1 & bh7_w33_8_c1 & bh7_w33_7_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid229_In1_c1 <= "" & bh7_w34_9_c1 & bh7_w34_8_c1;
   bh7_w33_11_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid229_Out0_c1(0);
   bh7_w34_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid229_Out0_c1(1);
   bh7_w35_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid229_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid229: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid229_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid229_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid229_Out0_copy230_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid229_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid229_Out0_copy230_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid231_In0_c1 <= "" & bh7_w35_9_c1 & bh7_w35_8_c1 & bh7_w35_7_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid231_In1_c1 <= "" & bh7_w36_9_c1 & bh7_w36_8_c1;
   bh7_w35_11_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid231_Out0_c1(0);
   bh7_w36_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid231_Out0_c1(1);
   bh7_w37_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid231_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid231: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid231_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid231_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid231_Out0_copy232_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid231_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid231_Out0_copy232_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid233_In0_c1 <= "" & bh7_w37_9_c1 & bh7_w37_8_c1 & bh7_w37_7_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid233_In1_c1 <= "" & bh7_w38_9_c1 & bh7_w38_8_c1;
   bh7_w37_11_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid233_Out0_c1(0);
   bh7_w38_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid233_Out0_c1(1);
   bh7_w39_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid233_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid233: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid233_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid233_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid233_Out0_copy234_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid233_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid233_Out0_copy234_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid235_In0_c1 <= "" & bh7_w39_9_c1 & bh7_w39_8_c1 & bh7_w39_7_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid235_In1_c1 <= "" & bh7_w40_9_c1 & bh7_w40_8_c1;
   bh7_w39_11_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid235_Out0_c1(0);
   bh7_w40_10_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid235_Out0_c1(1);
   bh7_w41_8_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid235_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid235: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid235_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid235_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid235_Out0_copy236_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid235_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid235_Out0_copy236_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid237_In0_c1 <= "" & bh7_w41_4_c1 & bh7_w41_7_c1 & bh7_w41_6_c1 & bh7_w41_5_c1;
   Compressor_14_3_Freq800_uid164_bh7_uid237_In1_c0 <= "" & "0";
   bh7_w41_9_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid237_Out0_c1(0);
   bh7_w42_8_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid237_Out0_c1(1);
   bh7_w43_7_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid237_Out0_c1(2);
   Compressor_14_3_Freq800_uid164_uid237: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid237_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid237_In1_c1,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid237_Out0_copy238_c1);
   Compressor_14_3_Freq800_uid164_bh7_uid237_Out0_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid237_Out0_copy238_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid160_bh7_uid239_In0_c1 <= "" & bh7_w42_7_c1 & bh7_w42_6_c1 & bh7_w42_5_c1;
   bh7_w42_9_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid239_Out0_c1(0);
   bh7_w43_8_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid239_Out0_c1(1);
   Compressor_3_2_Freq800_uid160_uid239: Compressor_3_2_Freq800_uid160
      port map ( X0 => Compressor_3_2_Freq800_uid160_bh7_uid239_In0_c1,
                 R => Compressor_3_2_Freq800_uid160_bh7_uid239_Out0_copy240_c1);
   Compressor_3_2_Freq800_uid160_bh7_uid239_Out0_c1 <= Compressor_3_2_Freq800_uid160_bh7_uid239_Out0_copy240_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid241_In0_c1 <= "" & bh7_w43_6_c1 & bh7_w43_5_c1 & bh7_w43_4_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid241_In1_c1 <= "" & bh7_w44_2_c1 & bh7_w44_4_c1;
   bh7_w43_9_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid241_Out0_c1(0);
   bh7_w44_5_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid241_Out0_c1(1);
   bh7_w45_4_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid241_Out0_c1(2);
   Compressor_23_3_Freq800_uid156_uid241: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid241_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid241_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid241_Out0_copy242_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid241_Out0_c1 <= Compressor_23_3_Freq800_uid156_bh7_uid241_Out0_copy242_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid243_In0_c1 <= "" & bh7_w45_3_c1 & bh7_w45_2_c1 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid243_In1_c1 <= "" & bh7_w46_2_c1;
   bh7_w45_5_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid243_Out0_c1(0);
   bh7_w46_3_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid243_Out0_c1(1);
   bh7_w47_1_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid243_Out0_c1(2);
   Compressor_14_3_Freq800_uid164_uid243: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid243_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid243_In1_c1,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid243_Out0_copy244_c1);
   Compressor_14_3_Freq800_uid164_bh7_uid243_Out0_c1 <= Compressor_14_3_Freq800_uid164_bh7_uid243_Out0_copy244_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid245_In0_c1 <= "" & bh7_w22_8_c1 & bh7_w22_7_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid245_In1_c1 <= "" & bh7_w23_10_c1 & bh7_w23_11_c1;
   bh7_w22_9_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_c2(0);
   bh7_w23_12_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_c2(1);
   bh7_w24_10_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid245: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid245_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid245_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_copy246_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid245_Out0_copy246_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid247_In0_c1 <= "" & bh7_w25_11_c1 & bh7_w25_10_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid247_In1_c1 <= "" & bh7_w26_7_c1 & bh7_w26_10_c1;
   bh7_w25_12_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_c2(0);
   bh7_w26_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_c2(1);
   bh7_w27_12_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid247: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid247_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid247_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_copy248_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid247_Out0_copy248_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid249_In0_c1 <= "" & bh7_w27_11_c1 & bh7_w27_10_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid249_In1_c1 <= "" & bh7_w28_7_c1 & bh7_w28_10_c1;
   bh7_w27_13_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_c2(0);
   bh7_w28_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_c2(1);
   bh7_w29_12_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid249: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid249_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid249_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_copy250_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid249_Out0_copy250_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid251_In0_c1 <= "" & bh7_w29_11_c1 & bh7_w29_10_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid251_In1_c1 <= "" & bh7_w30_7_c1 & bh7_w30_10_c1;
   bh7_w29_13_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_c2(0);
   bh7_w30_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_c2(1);
   bh7_w31_12_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid251: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid251_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid251_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_copy252_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid251_Out0_copy252_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid253_In0_c1 <= "" & bh7_w31_11_c1 & bh7_w31_10_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid253_In1_c1 <= "" & bh7_w32_7_c1 & bh7_w32_10_c1;
   bh7_w31_13_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_c2(0);
   bh7_w32_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_c2(1);
   bh7_w33_12_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid253: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid253_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid253_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_copy254_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid253_Out0_copy254_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid255_In0_c1 <= "" & bh7_w33_11_c1 & bh7_w33_10_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid255_In1_c1 <= "" & bh7_w34_7_c1 & bh7_w34_10_c1;
   bh7_w33_13_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_c2(0);
   bh7_w34_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_c2(1);
   bh7_w35_12_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid255: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid255_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid255_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_copy256_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid255_Out0_copy256_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid257_In0_c1 <= "" & bh7_w35_11_c1 & bh7_w35_10_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid257_In1_c1 <= "" & bh7_w36_7_c1 & bh7_w36_10_c1;
   bh7_w35_13_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_c2(0);
   bh7_w36_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_c2(1);
   bh7_w37_12_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid257: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid257_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid257_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_copy258_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid257_Out0_copy258_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid259_In0_c1 <= "" & bh7_w37_11_c1 & bh7_w37_10_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid259_In1_c1 <= "" & bh7_w38_7_c1 & bh7_w38_10_c1;
   bh7_w37_13_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_c2(0);
   bh7_w38_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_c2(1);
   bh7_w39_12_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid259: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid259_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid259_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_copy260_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid259_Out0_copy260_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid261_In0_c1 <= "" & bh7_w39_11_c1 & bh7_w39_10_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid261_In1_c1 <= "" & bh7_w40_7_c1 & bh7_w40_10_c1;
   bh7_w39_13_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_c2(0);
   bh7_w40_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_c2(1);
   bh7_w41_10_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid261: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid261_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid261_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_copy262_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid261_Out0_copy262_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid263_In0_c1 <= "" & bh7_w41_9_c1 & bh7_w41_8_c1 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid263_In1_c1 <= "" & bh7_w42_8_c1 & bh7_w42_9_c1;
   bh7_w41_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_c2(0);
   bh7_w42_10_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_c2(1);
   bh7_w43_10_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid263: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid263_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid263_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_copy264_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid263_Out0_copy264_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid265_In0_c1 <= "" & bh7_w43_7_c1 & bh7_w43_9_c1 & bh7_w43_8_c1;
   Compressor_23_3_Freq800_uid156_bh7_uid265_In1_c1 <= "" & bh7_w44_3_c1 & bh7_w44_5_c1;
   bh7_w43_11_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_c2(0);
   bh7_w44_6_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_c2(1);
   bh7_w45_6_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_c2(2);
   Compressor_23_3_Freq800_uid156_uid265: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid265_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid265_In1_c1,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_copy266_c1);
   Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_c2 <= Compressor_23_3_Freq800_uid156_bh7_uid265_Out0_copy266_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid267_In0_c1 <= "" & bh7_w45_5_c1 & bh7_w45_4_c1 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid267_In1_c1 <= "" & bh7_w46_3_c1;
   bh7_w45_7_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_c2(0);
   bh7_w46_4_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_c2(1);
   bh7_w47_2_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid267: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid267_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid267_In1_c1,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_copy268_c1);
   Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid267_Out0_copy268_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid160_bh7_uid269_In0_c1 <= "" & bh7_w47_0_c1 & bh7_w47_1_c1 & "0";
   bh7_w47_3_c2 <= Compressor_3_2_Freq800_uid160_bh7_uid269_Out0_c2(0);
   Compressor_3_2_Freq800_uid160_uid269: Compressor_3_2_Freq800_uid160
      port map ( X0 => Compressor_3_2_Freq800_uid160_bh7_uid269_In0_c1,
                 R => Compressor_3_2_Freq800_uid160_bh7_uid269_Out0_copy270_c1);
   Compressor_3_2_Freq800_uid160_bh7_uid269_Out0_c2 <= Compressor_3_2_Freq800_uid160_bh7_uid269_Out0_copy270_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid271_In0_c2 <= "" & bh7_w24_9_c2 & bh7_w24_10_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid271_In1_c2 <= "" & bh7_w25_12_c2;
   bh7_w24_11_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid271_Out0_c2(0);
   bh7_w25_13_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid271_Out0_c2(1);
   bh7_w26_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid271_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid271: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid271_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid271_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid271_Out0_copy272_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid271_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid271_Out0_copy272_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid273_In0_c2 <= "" & bh7_w27_13_c2 & bh7_w27_12_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid273_In1_c2 <= "" & bh7_w28_11_c2;
   bh7_w27_14_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid273_Out0_c2(0);
   bh7_w28_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid273_Out0_c2(1);
   bh7_w29_14_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid273_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid273: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid273_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid273_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid273_Out0_copy274_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid273_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid273_Out0_copy274_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid275_In0_c2 <= "" & bh7_w29_13_c2 & bh7_w29_12_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid275_In1_c2 <= "" & bh7_w30_11_c2;
   bh7_w29_15_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid275_Out0_c2(0);
   bh7_w30_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid275_Out0_c2(1);
   bh7_w31_14_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid275_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid275: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid275_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid275_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid275_Out0_copy276_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid275_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid275_Out0_copy276_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid277_In0_c2 <= "" & bh7_w31_13_c2 & bh7_w31_12_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid277_In1_c2 <= "" & bh7_w32_11_c2;
   bh7_w31_15_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid277_Out0_c2(0);
   bh7_w32_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid277_Out0_c2(1);
   bh7_w33_14_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid277_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid277: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid277_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid277_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid277_Out0_copy278_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid277_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid277_Out0_copy278_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid279_In0_c2 <= "" & bh7_w33_13_c2 & bh7_w33_12_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid279_In1_c2 <= "" & bh7_w34_11_c2;
   bh7_w33_15_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid279_Out0_c2(0);
   bh7_w34_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid279_Out0_c2(1);
   bh7_w35_14_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid279_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid279: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid279_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid279_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid279_Out0_copy280_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid279_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid279_Out0_copy280_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid281_In0_c2 <= "" & bh7_w35_13_c2 & bh7_w35_12_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid281_In1_c2 <= "" & bh7_w36_11_c2;
   bh7_w35_15_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid281_Out0_c2(0);
   bh7_w36_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid281_Out0_c2(1);
   bh7_w37_14_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid281_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid281: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid281_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid281_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid281_Out0_copy282_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid281_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid281_Out0_copy282_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid283_In0_c2 <= "" & bh7_w37_13_c2 & bh7_w37_12_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid283_In1_c2 <= "" & bh7_w38_11_c2;
   bh7_w37_15_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid283_Out0_c2(0);
   bh7_w38_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid283_Out0_c2(1);
   bh7_w39_14_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid283_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid283: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid283_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid283_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid283_Out0_copy284_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid283_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid283_Out0_copy284_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid285_In0_c2 <= "" & bh7_w39_13_c2 & bh7_w39_12_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid285_In1_c2 <= "" & bh7_w40_11_c2;
   bh7_w39_15_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid285_Out0_c2(0);
   bh7_w40_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid285_Out0_c2(1);
   bh7_w41_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid285_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid285: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid285_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid285_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid285_Out0_copy286_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid285_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid285_Out0_copy286_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid287_In0_c2 <= "" & bh7_w41_11_c2 & bh7_w41_10_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid287_In1_c2 <= "" & bh7_w42_10_c2;
   bh7_w41_13_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid287_Out0_c2(0);
   bh7_w42_11_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid287_Out0_c2(1);
   bh7_w43_12_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid287_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid287: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid287_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid287_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid287_Out0_copy288_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid287_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid287_Out0_copy288_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid289_In0_c2 <= "" & bh7_w43_10_c2 & bh7_w43_11_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid289_In1_c2 <= "" & bh7_w44_6_c2;
   bh7_w43_13_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid289_Out0_c2(0);
   bh7_w44_7_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid289_Out0_c2(1);
   bh7_w45_8_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid289_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid289: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid289_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid289_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid289_Out0_copy290_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid289_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid289_Out0_copy290_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid291_In0_c2 <= "" & bh7_w45_6_c2 & bh7_w45_7_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid291_In1_c2 <= "" & bh7_w46_4_c2;
   bh7_w45_9_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid291_Out0_c2(0);
   bh7_w46_5_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid291_Out0_c2(1);
   bh7_w47_4_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid291_Out0_c2(2);
   Compressor_14_3_Freq800_uid164_uid291: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid291_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid291_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid291_Out0_copy292_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid291_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid291_Out0_copy292_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid293_In0_c2 <= "" & bh7_w47_3_c2 & bh7_w47_2_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid293_In1_c0 <= "" & "0";
   bh7_w47_5_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid293_Out0_c2(0);
   Compressor_14_3_Freq800_uid164_uid293: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid293_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid293_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid293_Out0_copy294_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid293_Out0_c2 <= Compressor_14_3_Freq800_uid164_bh7_uid293_Out0_copy294_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid295_In0_c2 <= "" & bh7_w26_11_c2 & bh7_w26_12_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid295_In1_c2 <= "" & bh7_w27_14_c2;
   bh7_w26_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_c3(0);
   bh7_w27_15_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_c3(1);
   bh7_w28_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid295: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid295_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid295_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_copy296_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid295_Out0_copy296_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid297_In0_c2 <= "" & bh7_w29_15_c2 & bh7_w29_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid297_In1_c2 <= "" & bh7_w30_12_c2;
   bh7_w29_16_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_c3(0);
   bh7_w30_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_c3(1);
   bh7_w31_16_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid297: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid297_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid297_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_copy298_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid297_Out0_copy298_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid299_In0_c2 <= "" & bh7_w31_15_c2 & bh7_w31_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid299_In1_c2 <= "" & bh7_w32_12_c2;
   bh7_w31_17_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_c3(0);
   bh7_w32_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_c3(1);
   bh7_w33_16_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid299: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid299_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid299_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_copy300_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid299_Out0_copy300_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid301_In0_c2 <= "" & bh7_w33_15_c2 & bh7_w33_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid301_In1_c2 <= "" & bh7_w34_12_c2;
   bh7_w33_17_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_c3(0);
   bh7_w34_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_c3(1);
   bh7_w35_16_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid301: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid301_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid301_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_copy302_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid301_Out0_copy302_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid303_In0_c2 <= "" & bh7_w35_15_c2 & bh7_w35_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid303_In1_c2 <= "" & bh7_w36_12_c2;
   bh7_w35_17_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_c3(0);
   bh7_w36_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_c3(1);
   bh7_w37_16_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid303: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid303_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid303_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_copy304_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid303_Out0_copy304_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid305_In0_c2 <= "" & bh7_w37_15_c2 & bh7_w37_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid305_In1_c2 <= "" & bh7_w38_12_c2;
   bh7_w37_17_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_c3(0);
   bh7_w38_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_c3(1);
   bh7_w39_16_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid305: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid305_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid305_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_copy306_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid305_Out0_copy306_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid307_In0_c2 <= "" & bh7_w39_15_c2 & bh7_w39_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid307_In1_c2 <= "" & bh7_w40_12_c2;
   bh7_w39_17_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_c3(0);
   bh7_w40_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_c3(1);
   bh7_w41_14_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid307: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid307_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid307_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_copy308_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid307_Out0_copy308_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid309_In0_c2 <= "" & bh7_w41_13_c2 & bh7_w41_12_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid309_In1_c2 <= "" & bh7_w42_11_c2;
   bh7_w41_15_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_c3(0);
   bh7_w42_12_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_c3(1);
   bh7_w43_14_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid309: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid309_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid309_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_copy310_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid309_Out0_copy310_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid311_In0_c2 <= "" & bh7_w43_12_c2 & bh7_w43_13_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid311_In1_c2 <= "" & bh7_w44_7_c2;
   bh7_w43_15_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_c3(0);
   bh7_w44_8_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_c3(1);
   bh7_w45_10_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid311: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid311_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid311_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_copy312_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid311_Out0_copy312_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid313_In0_c2 <= "" & bh7_w45_8_c2 & bh7_w45_9_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid313_In1_c2 <= "" & bh7_w46_5_c2;
   bh7_w45_11_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_c3(0);
   bh7_w46_6_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_c3(1);
   bh7_w47_6_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid313: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid313_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid313_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_copy314_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid313_Out0_copy314_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid315_In0_c2 <= "" & bh7_w47_4_c2 & bh7_w47_5_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid315_In1_c0 <= "" & "0";
   bh7_w47_7_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid315_Out0_c3(0);
   Compressor_14_3_Freq800_uid164_uid315: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid315_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid315_In1_c2,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid315_Out0_copy316_c2);
   Compressor_14_3_Freq800_uid164_bh7_uid315_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid315_Out0_copy316_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid317_In0_c2 <= "" & bh7_w17_1_c2 & bh7_w17_0_c2 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid317_In1_c2 <= "" & bh7_w18_2_c2 & bh7_w18_0_c2;
   bh7_w17_2_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_c3(0);
   bh7_w18_3_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_c3(1);
   bh7_w19_4_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid317: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid317_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid317_In1_c2,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_copy318_c2);
   Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid317_Out0_copy318_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid319_In0_c2 <= "" & bh7_w19_3_c2 & bh7_w19_0_c2 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid319_In1_c2 <= "" & bh7_w20_6_c2 & bh7_w20_0_c2;
   bh7_w19_5_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_c3(0);
   bh7_w20_7_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_c3(1);
   bh7_w21_8_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid319: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid319_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid319_In1_c2,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_copy320_c2);
   Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid319_Out0_copy320_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid321_In0_c2 <= "" & bh7_w21_7_c2 & bh7_w21_0_c2 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid321_In1_c2 <= "" & bh7_w22_9_c2 & bh7_w22_0_c2;
   bh7_w21_9_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_c3(0);
   bh7_w22_10_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_c3(1);
   bh7_w23_13_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid321: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid321_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid321_In1_c2,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_copy322_c2);
   Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid321_Out0_copy322_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid323_In0_c2 <= "" & bh7_w23_12_c2 & bh7_w23_0_c2 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid323_In1_c2 <= "" & bh7_w24_11_c2 & bh7_w24_0_c2;
   bh7_w23_14_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_c3(0);
   bh7_w24_12_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_c3(1);
   bh7_w25_14_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid323: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid323_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid323_In1_c2,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_copy324_c2);
   Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid323_Out0_copy324_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid325_In0_c2 <= "" & bh7_w25_13_c2 & bh7_w25_0_c2 & "0";
   Compressor_23_3_Freq800_uid156_bh7_uid325_In1_c3 <= "" & bh7_w26_0_c3 & bh7_w26_13_c3;
   bh7_w25_15_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid325_Out0_c3(0);
   bh7_w26_14_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid325_Out0_c3(1);
   bh7_w27_16_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid325_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid325: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid325_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid325_In1_c3,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid325_Out0_copy326_c3);
   Compressor_23_3_Freq800_uid156_bh7_uid325_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid325_Out0_copy326_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid160_bh7_uid327_In0_c3 <= "" & bh7_w27_0_c3 & bh7_w27_15_c3 & "0";
   bh7_w27_17_c3 <= Compressor_3_2_Freq800_uid160_bh7_uid327_Out0_c3(0);
   bh7_w28_14_c3 <= Compressor_3_2_Freq800_uid160_bh7_uid327_Out0_c3(1);
   Compressor_3_2_Freq800_uid160_uid327: Compressor_3_2_Freq800_uid160
      port map ( X0 => Compressor_3_2_Freq800_uid160_bh7_uid327_In0_c3,
                 R => Compressor_3_2_Freq800_uid160_bh7_uid327_Out0_copy328_c3);
   Compressor_3_2_Freq800_uid160_bh7_uid327_Out0_c3 <= Compressor_3_2_Freq800_uid160_bh7_uid327_Out0_copy328_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid329_In0_c3 <= "" & bh7_w28_12_c3 & bh7_w28_0_c3 & bh7_w28_13_c3;
   Compressor_23_3_Freq800_uid156_bh7_uid329_In1_c3 <= "" & bh7_w29_0_c3 & bh7_w29_16_c3;
   bh7_w28_15_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid329_Out0_c3(0);
   bh7_w29_17_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid329_Out0_c3(1);
   bh7_w30_14_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid329_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid329: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid329_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid329_In1_c3,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid329_Out0_copy330_c3);
   Compressor_23_3_Freq800_uid156_bh7_uid329_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid329_Out0_copy330_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid160_bh7_uid331_In0_c3 <= "" & bh7_w30_0_c3 & bh7_w30_13_c3 & "0";
   bh7_w30_15_c3 <= Compressor_3_2_Freq800_uid160_bh7_uid331_Out0_c3(0);
   bh7_w31_18_c3 <= Compressor_3_2_Freq800_uid160_bh7_uid331_Out0_c3(1);
   Compressor_3_2_Freq800_uid160_uid331: Compressor_3_2_Freq800_uid160
      port map ( X0 => Compressor_3_2_Freq800_uid160_bh7_uid331_In0_c3,
                 R => Compressor_3_2_Freq800_uid160_bh7_uid331_Out0_copy332_c3);
   Compressor_3_2_Freq800_uid160_bh7_uid331_Out0_c3 <= Compressor_3_2_Freq800_uid160_bh7_uid331_Out0_copy332_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid333_In0_c3 <= "" & bh7_w31_0_c3 & bh7_w31_17_c3 & bh7_w31_16_c3;
   Compressor_23_3_Freq800_uid156_bh7_uid333_In1_c3 <= "" & bh7_w32_0_c3 & bh7_w32_13_c3;
   bh7_w31_19_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid333_Out0_c3(0);
   bh7_w32_14_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid333_Out0_c3(1);
   bh7_w33_18_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid333_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid333: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid333_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid333_In1_c3,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid333_Out0_copy334_c3);
   Compressor_23_3_Freq800_uid156_bh7_uid333_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid333_Out0_copy334_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid335_In0_c3 <= "" & bh7_w33_0_c3 & bh7_w33_17_c3 & bh7_w33_16_c3;
   Compressor_23_3_Freq800_uid156_bh7_uid335_In1_c3 <= "" & bh7_w34_0_c3 & bh7_w34_13_c3;
   bh7_w33_19_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid335_Out0_c3(0);
   bh7_w34_14_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid335_Out0_c3(1);
   bh7_w35_18_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid335_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid335: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid335_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid335_In1_c3,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid335_Out0_copy336_c3);
   Compressor_23_3_Freq800_uid156_bh7_uid335_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid335_Out0_copy336_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid337_In0_c3 <= "" & bh7_w35_0_c3 & bh7_w35_17_c3 & bh7_w35_16_c3;
   Compressor_23_3_Freq800_uid156_bh7_uid337_In1_c3 <= "" & bh7_w36_0_c3 & bh7_w36_13_c3;
   bh7_w35_19_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid337_Out0_c3(0);
   bh7_w36_14_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid337_Out0_c3(1);
   bh7_w37_18_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid337_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid337: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid337_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid337_In1_c3,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid337_Out0_copy338_c3);
   Compressor_23_3_Freq800_uid156_bh7_uid337_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid337_Out0_copy338_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid339_In0_c3 <= "" & bh7_w37_0_c3 & bh7_w37_17_c3 & bh7_w37_16_c3;
   Compressor_23_3_Freq800_uid156_bh7_uid339_In1_c3 <= "" & bh7_w38_0_c3 & bh7_w38_13_c3;
   bh7_w37_19_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid339_Out0_c3(0);
   bh7_w38_14_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid339_Out0_c3(1);
   bh7_w39_18_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid339_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid339: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid339_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid339_In1_c3,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid339_Out0_copy340_c3);
   Compressor_23_3_Freq800_uid156_bh7_uid339_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid339_Out0_copy340_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid156_bh7_uid341_In0_c3 <= "" & bh7_w39_0_c3 & bh7_w39_17_c3 & bh7_w39_16_c3;
   Compressor_23_3_Freq800_uid156_bh7_uid341_In1_c3 <= "" & bh7_w40_0_c3 & bh7_w40_13_c3;
   bh7_w39_19_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid341_Out0_c3(0);
   bh7_w40_14_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid341_Out0_c3(1);
   bh7_w41_16_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid341_Out0_c3(2);
   Compressor_23_3_Freq800_uid156_uid341: Compressor_23_3_Freq800_uid156
      port map ( X0 => Compressor_23_3_Freq800_uid156_bh7_uid341_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid156_bh7_uid341_In1_c3,
                 R => Compressor_23_3_Freq800_uid156_bh7_uid341_Out0_copy342_c3);
   Compressor_23_3_Freq800_uid156_bh7_uid341_Out0_c3 <= Compressor_23_3_Freq800_uid156_bh7_uid341_Out0_copy342_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid343_In0_c3 <= "" & bh7_w41_15_c3 & bh7_w41_14_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid343_In1_c3 <= "" & bh7_w42_12_c3;
   bh7_w41_17_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid343_Out0_c3(0);
   bh7_w42_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid343_Out0_c3(1);
   bh7_w43_16_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid343_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid343: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid343_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid343_In1_c3,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid343_Out0_copy344_c3);
   Compressor_14_3_Freq800_uid164_bh7_uid343_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid343_Out0_copy344_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid345_In0_c3 <= "" & bh7_w43_14_c3 & bh7_w43_15_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid345_In1_c3 <= "" & bh7_w44_8_c3;
   bh7_w43_17_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid345_Out0_c3(0);
   bh7_w44_9_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid345_Out0_c3(1);
   bh7_w45_12_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid345_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid345: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid345_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid345_In1_c3,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid345_Out0_copy346_c3);
   Compressor_14_3_Freq800_uid164_bh7_uid345_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid345_Out0_copy346_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid347_In0_c3 <= "" & bh7_w45_10_c3 & bh7_w45_11_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid347_In1_c3 <= "" & bh7_w46_6_c3;
   bh7_w45_13_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid347_Out0_c3(0);
   bh7_w46_7_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid347_Out0_c3(1);
   bh7_w47_8_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid347_Out0_c3(2);
   Compressor_14_3_Freq800_uid164_uid347: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid347_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid347_In1_c3,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid347_Out0_copy348_c3);
   Compressor_14_3_Freq800_uid164_bh7_uid347_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid347_Out0_copy348_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid164_bh7_uid349_In0_c3 <= "" & bh7_w47_6_c3 & bh7_w47_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c0 <= "" & "0";
   bh7_w47_9_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid349_Out0_c3(0);
   Compressor_14_3_Freq800_uid164_uid349: Compressor_14_3_Freq800_uid164
      port map ( X0 => Compressor_14_3_Freq800_uid164_bh7_uid349_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid164_bh7_uid349_In1_c3,
                 R => Compressor_14_3_Freq800_uid164_bh7_uid349_Out0_copy350_c3);
   Compressor_14_3_Freq800_uid164_bh7_uid349_Out0_c3 <= Compressor_14_3_Freq800_uid164_bh7_uid349_Out0_copy350_c3; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh7_18_c3 <= bh7_w18_3_c3 & bh7_w17_2_c3 & bh7_w16_0_c3 & bh7_w15_0_c3 & bh7_w14_0_c3 & bh7_w13_0_c3 & bh7_w12_0_c3 & bh7_w11_0_c3 & bh7_w10_0_c3 & bh7_w9_0_c3 & bh7_w8_0_c3 & bh7_w7_0_c3 & bh7_w6_0_c3 & bh7_w5_0_c3 & bh7_w4_0_c3 & bh7_w3_0_c3 & bh7_w2_0_c3 & bh7_w1_0_c3 & bh7_w0_0_c3;

   bitheapFinalAdd_bh7_In0_c3 <= "0" & bh7_w47_8_c3 & bh7_w46_7_c3 & bh7_w45_12_c3 & bh7_w44_9_c3 & bh7_w43_16_c3 & bh7_w42_13_c3 & bh7_w41_17_c3 & bh7_w40_14_c3 & bh7_w39_19_c3 & bh7_w38_14_c3 & bh7_w37_19_c3 & bh7_w36_14_c3 & bh7_w35_19_c3 & bh7_w34_14_c3 & bh7_w33_19_c3 & bh7_w32_14_c3 & bh7_w31_19_c3 & bh7_w30_15_c3 & bh7_w29_17_c3 & bh7_w28_15_c3 & bh7_w27_17_c3 & bh7_w26_14_c3 & bh7_w25_14_c3 & bh7_w24_12_c3 & bh7_w23_14_c3 & bh7_w22_10_c3 & bh7_w21_9_c3 & bh7_w20_7_c3 & bh7_w19_5_c3;
   bitheapFinalAdd_bh7_In1_c3 <= "0" & bh7_w47_9_c3 & "0" & bh7_w45_13_c3 & "0" & bh7_w43_17_c3 & "0" & bh7_w41_16_c3 & "0" & bh7_w39_18_c3 & "0" & bh7_w37_18_c3 & "0" & bh7_w35_18_c3 & "0" & bh7_w33_18_c3 & "0" & bh7_w31_18_c3 & bh7_w30_14_c3 & "0" & bh7_w28_14_c3 & bh7_w27_16_c3 & "0" & bh7_w25_15_c3 & "0" & bh7_w23_13_c3 & "0" & bh7_w21_8_c3 & "0" & bh7_w19_4_c3;
   bitheapFinalAdd_bh7_Cin_c0 <= '0';

   bitheapFinalAdd_bh7: IntAdder_30_Freq800_uid352
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 Cin => bitheapFinalAdd_bh7_Cin_c0,
                 X => bitheapFinalAdd_bh7_In0_c3,
                 Y => bitheapFinalAdd_bh7_In1_c3,
                 R => bitheapFinalAdd_bh7_Out_c13);
   bitheapResult_bh7_c13 <= bitheapFinalAdd_bh7_Out_c13(28 downto 0) & tmp_bitheapResult_bh7_18_c13;
   R <= bitheapResult_bh7_c13(47 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_Freq800_uid355
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_Freq800_uid355 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26 : in std_logic;
          X : in  std_logic_vector(32 downto 0);
          Y : in  std_logic_vector(32 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_Freq800_uid355 is
signal Cin_1_c15, Cin_1_c16 :  std_logic;
signal X_1_c14, X_1_c15, X_1_c16 :  std_logic_vector(3 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3, Y_1_c4, Y_1_c5, Y_1_c6, Y_1_c7, Y_1_c8, Y_1_c9, Y_1_c10, Y_1_c11, Y_1_c12, Y_1_c13, Y_1_c14, Y_1_c15, Y_1_c16 :  std_logic_vector(3 downto 0);
signal S_1_c16 :  std_logic_vector(3 downto 0);
signal R_1_c16, R_1_c17, R_1_c18, R_1_c19, R_1_c20, R_1_c21, R_1_c22, R_1_c23, R_1_c24, R_1_c25, R_1_c26 :  std_logic_vector(2 downto 0);
signal Cin_2_c16, Cin_2_c17 :  std_logic;
signal X_2_c14, X_2_c15, X_2_c16, X_2_c17 :  std_logic_vector(3 downto 0);
signal Y_2_c0, Y_2_c1, Y_2_c2, Y_2_c3, Y_2_c4, Y_2_c5, Y_2_c6, Y_2_c7, Y_2_c8, Y_2_c9, Y_2_c10, Y_2_c11, Y_2_c12, Y_2_c13, Y_2_c14, Y_2_c15, Y_2_c16, Y_2_c17 :  std_logic_vector(3 downto 0);
signal S_2_c17 :  std_logic_vector(3 downto 0);
signal R_2_c17, R_2_c18, R_2_c19, R_2_c20, R_2_c21, R_2_c22, R_2_c23, R_2_c24, R_2_c25, R_2_c26 :  std_logic_vector(2 downto 0);
signal Cin_3_c17, Cin_3_c18 :  std_logic;
signal X_3_c14, X_3_c15, X_3_c16, X_3_c17, X_3_c18 :  std_logic_vector(3 downto 0);
signal Y_3_c0, Y_3_c1, Y_3_c2, Y_3_c3, Y_3_c4, Y_3_c5, Y_3_c6, Y_3_c7, Y_3_c8, Y_3_c9, Y_3_c10, Y_3_c11, Y_3_c12, Y_3_c13, Y_3_c14, Y_3_c15, Y_3_c16, Y_3_c17, Y_3_c18 :  std_logic_vector(3 downto 0);
signal S_3_c18 :  std_logic_vector(3 downto 0);
signal R_3_c18, R_3_c19, R_3_c20, R_3_c21, R_3_c22, R_3_c23, R_3_c24, R_3_c25, R_3_c26 :  std_logic_vector(2 downto 0);
signal Cin_4_c18, Cin_4_c19 :  std_logic;
signal X_4_c14, X_4_c15, X_4_c16, X_4_c17, X_4_c18, X_4_c19 :  std_logic_vector(3 downto 0);
signal Y_4_c0, Y_4_c1, Y_4_c2, Y_4_c3, Y_4_c4, Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8, Y_4_c9, Y_4_c10, Y_4_c11, Y_4_c12, Y_4_c13, Y_4_c14, Y_4_c15, Y_4_c16, Y_4_c17, Y_4_c18, Y_4_c19 :  std_logic_vector(3 downto 0);
signal S_4_c19 :  std_logic_vector(3 downto 0);
signal R_4_c19, R_4_c20, R_4_c21, R_4_c22, R_4_c23, R_4_c24, R_4_c25, R_4_c26 :  std_logic_vector(2 downto 0);
signal Cin_5_c19, Cin_5_c20 :  std_logic;
signal X_5_c14, X_5_c15, X_5_c16, X_5_c17, X_5_c18, X_5_c19, X_5_c20 :  std_logic_vector(3 downto 0);
signal Y_5_c0, Y_5_c1, Y_5_c2, Y_5_c3, Y_5_c4, Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9, Y_5_c10, Y_5_c11, Y_5_c12, Y_5_c13, Y_5_c14, Y_5_c15, Y_5_c16, Y_5_c17, Y_5_c18, Y_5_c19, Y_5_c20 :  std_logic_vector(3 downto 0);
signal S_5_c20 :  std_logic_vector(3 downto 0);
signal R_5_c20, R_5_c21, R_5_c22, R_5_c23, R_5_c24, R_5_c25, R_5_c26 :  std_logic_vector(2 downto 0);
signal Cin_6_c20, Cin_6_c21 :  std_logic;
signal X_6_c14, X_6_c15, X_6_c16, X_6_c17, X_6_c18, X_6_c19, X_6_c20, X_6_c21 :  std_logic_vector(3 downto 0);
signal Y_6_c0, Y_6_c1, Y_6_c2, Y_6_c3, Y_6_c4, Y_6_c5, Y_6_c6, Y_6_c7, Y_6_c8, Y_6_c9, Y_6_c10, Y_6_c11, Y_6_c12, Y_6_c13, Y_6_c14, Y_6_c15, Y_6_c16, Y_6_c17, Y_6_c18, Y_6_c19, Y_6_c20, Y_6_c21 :  std_logic_vector(3 downto 0);
signal S_6_c21 :  std_logic_vector(3 downto 0);
signal R_6_c21, R_6_c22, R_6_c23, R_6_c24, R_6_c25, R_6_c26 :  std_logic_vector(2 downto 0);
signal Cin_7_c21, Cin_7_c22 :  std_logic;
signal X_7_c14, X_7_c15, X_7_c16, X_7_c17, X_7_c18, X_7_c19, X_7_c20, X_7_c21, X_7_c22 :  std_logic_vector(3 downto 0);
signal Y_7_c0, Y_7_c1, Y_7_c2, Y_7_c3, Y_7_c4, Y_7_c5, Y_7_c6, Y_7_c7, Y_7_c8, Y_7_c9, Y_7_c10, Y_7_c11, Y_7_c12, Y_7_c13, Y_7_c14, Y_7_c15, Y_7_c16, Y_7_c17, Y_7_c18, Y_7_c19, Y_7_c20, Y_7_c21, Y_7_c22 :  std_logic_vector(3 downto 0);
signal S_7_c22 :  std_logic_vector(3 downto 0);
signal R_7_c22, R_7_c23, R_7_c24, R_7_c25, R_7_c26 :  std_logic_vector(2 downto 0);
signal Cin_8_c22, Cin_8_c23 :  std_logic;
signal X_8_c14, X_8_c15, X_8_c16, X_8_c17, X_8_c18, X_8_c19, X_8_c20, X_8_c21, X_8_c22, X_8_c23 :  std_logic_vector(3 downto 0);
signal Y_8_c0, Y_8_c1, Y_8_c2, Y_8_c3, Y_8_c4, Y_8_c5, Y_8_c6, Y_8_c7, Y_8_c8, Y_8_c9, Y_8_c10, Y_8_c11, Y_8_c12, Y_8_c13, Y_8_c14, Y_8_c15, Y_8_c16, Y_8_c17, Y_8_c18, Y_8_c19, Y_8_c20, Y_8_c21, Y_8_c22, Y_8_c23 :  std_logic_vector(3 downto 0);
signal S_8_c23 :  std_logic_vector(3 downto 0);
signal R_8_c23, R_8_c24, R_8_c25, R_8_c26 :  std_logic_vector(2 downto 0);
signal Cin_9_c23, Cin_9_c24 :  std_logic;
signal X_9_c14, X_9_c15, X_9_c16, X_9_c17, X_9_c18, X_9_c19, X_9_c20, X_9_c21, X_9_c22, X_9_c23, X_9_c24 :  std_logic_vector(3 downto 0);
signal Y_9_c0, Y_9_c1, Y_9_c2, Y_9_c3, Y_9_c4, Y_9_c5, Y_9_c6, Y_9_c7, Y_9_c8, Y_9_c9, Y_9_c10, Y_9_c11, Y_9_c12, Y_9_c13, Y_9_c14, Y_9_c15, Y_9_c16, Y_9_c17, Y_9_c18, Y_9_c19, Y_9_c20, Y_9_c21, Y_9_c22, Y_9_c23, Y_9_c24 :  std_logic_vector(3 downto 0);
signal S_9_c24 :  std_logic_vector(3 downto 0);
signal R_9_c24, R_9_c25, R_9_c26 :  std_logic_vector(2 downto 0);
signal Cin_10_c24, Cin_10_c25 :  std_logic;
signal X_10_c14, X_10_c15, X_10_c16, X_10_c17, X_10_c18, X_10_c19, X_10_c20, X_10_c21, X_10_c22, X_10_c23, X_10_c24, X_10_c25 :  std_logic_vector(3 downto 0);
signal Y_10_c0, Y_10_c1, Y_10_c2, Y_10_c3, Y_10_c4, Y_10_c5, Y_10_c6, Y_10_c7, Y_10_c8, Y_10_c9, Y_10_c10, Y_10_c11, Y_10_c12, Y_10_c13, Y_10_c14, Y_10_c15, Y_10_c16, Y_10_c17, Y_10_c18, Y_10_c19, Y_10_c20, Y_10_c21, Y_10_c22, Y_10_c23, Y_10_c24, Y_10_c25 :  std_logic_vector(3 downto 0);
signal S_10_c25 :  std_logic_vector(3 downto 0);
signal R_10_c25, R_10_c26 :  std_logic_vector(2 downto 0);
signal Cin_11_c25, Cin_11_c26 :  std_logic;
signal X_11_c14, X_11_c15, X_11_c16, X_11_c17, X_11_c18, X_11_c19, X_11_c20, X_11_c21, X_11_c22, X_11_c23, X_11_c24, X_11_c25, X_11_c26 :  std_logic_vector(3 downto 0);
signal Y_11_c0, Y_11_c1, Y_11_c2, Y_11_c3, Y_11_c4, Y_11_c5, Y_11_c6, Y_11_c7, Y_11_c8, Y_11_c9, Y_11_c10, Y_11_c11, Y_11_c12, Y_11_c13, Y_11_c14, Y_11_c15, Y_11_c16, Y_11_c17, Y_11_c18, Y_11_c19, Y_11_c20, Y_11_c21, Y_11_c22, Y_11_c23, Y_11_c24, Y_11_c25, Y_11_c26 :  std_logic_vector(3 downto 0);
signal S_11_c26 :  std_logic_vector(3 downto 0);
signal R_11_c26 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_1_c1 <= Y_1_c0;
               Y_2_c1 <= Y_2_c0;
               Y_3_c1 <= Y_3_c0;
               Y_4_c1 <= Y_4_c0;
               Y_5_c1 <= Y_5_c0;
               Y_6_c1 <= Y_6_c0;
               Y_7_c1 <= Y_7_c0;
               Y_8_c1 <= Y_8_c0;
               Y_9_c1 <= Y_9_c0;
               Y_10_c1 <= Y_10_c0;
               Y_11_c1 <= Y_11_c0;
            end if;
            if ce_2 = '1' then
               Y_1_c2 <= Y_1_c1;
               Y_2_c2 <= Y_2_c1;
               Y_3_c2 <= Y_3_c1;
               Y_4_c2 <= Y_4_c1;
               Y_5_c2 <= Y_5_c1;
               Y_6_c2 <= Y_6_c1;
               Y_7_c2 <= Y_7_c1;
               Y_8_c2 <= Y_8_c1;
               Y_9_c2 <= Y_9_c1;
               Y_10_c2 <= Y_10_c1;
               Y_11_c2 <= Y_11_c1;
            end if;
            if ce_3 = '1' then
               Y_1_c3 <= Y_1_c2;
               Y_2_c3 <= Y_2_c2;
               Y_3_c3 <= Y_3_c2;
               Y_4_c3 <= Y_4_c2;
               Y_5_c3 <= Y_5_c2;
               Y_6_c3 <= Y_6_c2;
               Y_7_c3 <= Y_7_c2;
               Y_8_c3 <= Y_8_c2;
               Y_9_c3 <= Y_9_c2;
               Y_10_c3 <= Y_10_c2;
               Y_11_c3 <= Y_11_c2;
            end if;
            if ce_4 = '1' then
               Y_1_c4 <= Y_1_c3;
               Y_2_c4 <= Y_2_c3;
               Y_3_c4 <= Y_3_c3;
               Y_4_c4 <= Y_4_c3;
               Y_5_c4 <= Y_5_c3;
               Y_6_c4 <= Y_6_c3;
               Y_7_c4 <= Y_7_c3;
               Y_8_c4 <= Y_8_c3;
               Y_9_c4 <= Y_9_c3;
               Y_10_c4 <= Y_10_c3;
               Y_11_c4 <= Y_11_c3;
            end if;
            if ce_5 = '1' then
               Y_1_c5 <= Y_1_c4;
               Y_2_c5 <= Y_2_c4;
               Y_3_c5 <= Y_3_c4;
               Y_4_c5 <= Y_4_c4;
               Y_5_c5 <= Y_5_c4;
               Y_6_c5 <= Y_6_c4;
               Y_7_c5 <= Y_7_c4;
               Y_8_c5 <= Y_8_c4;
               Y_9_c5 <= Y_9_c4;
               Y_10_c5 <= Y_10_c4;
               Y_11_c5 <= Y_11_c4;
            end if;
            if ce_6 = '1' then
               Y_1_c6 <= Y_1_c5;
               Y_2_c6 <= Y_2_c5;
               Y_3_c6 <= Y_3_c5;
               Y_4_c6 <= Y_4_c5;
               Y_5_c6 <= Y_5_c5;
               Y_6_c6 <= Y_6_c5;
               Y_7_c6 <= Y_7_c5;
               Y_8_c6 <= Y_8_c5;
               Y_9_c6 <= Y_9_c5;
               Y_10_c6 <= Y_10_c5;
               Y_11_c6 <= Y_11_c5;
            end if;
            if ce_7 = '1' then
               Y_1_c7 <= Y_1_c6;
               Y_2_c7 <= Y_2_c6;
               Y_3_c7 <= Y_3_c6;
               Y_4_c7 <= Y_4_c6;
               Y_5_c7 <= Y_5_c6;
               Y_6_c7 <= Y_6_c6;
               Y_7_c7 <= Y_7_c6;
               Y_8_c7 <= Y_8_c6;
               Y_9_c7 <= Y_9_c6;
               Y_10_c7 <= Y_10_c6;
               Y_11_c7 <= Y_11_c6;
            end if;
            if ce_8 = '1' then
               Y_1_c8 <= Y_1_c7;
               Y_2_c8 <= Y_2_c7;
               Y_3_c8 <= Y_3_c7;
               Y_4_c8 <= Y_4_c7;
               Y_5_c8 <= Y_5_c7;
               Y_6_c8 <= Y_6_c7;
               Y_7_c8 <= Y_7_c7;
               Y_8_c8 <= Y_8_c7;
               Y_9_c8 <= Y_9_c7;
               Y_10_c8 <= Y_10_c7;
               Y_11_c8 <= Y_11_c7;
            end if;
            if ce_9 = '1' then
               Y_1_c9 <= Y_1_c8;
               Y_2_c9 <= Y_2_c8;
               Y_3_c9 <= Y_3_c8;
               Y_4_c9 <= Y_4_c8;
               Y_5_c9 <= Y_5_c8;
               Y_6_c9 <= Y_6_c8;
               Y_7_c9 <= Y_7_c8;
               Y_8_c9 <= Y_8_c8;
               Y_9_c9 <= Y_9_c8;
               Y_10_c9 <= Y_10_c8;
               Y_11_c9 <= Y_11_c8;
            end if;
            if ce_10 = '1' then
               Y_1_c10 <= Y_1_c9;
               Y_2_c10 <= Y_2_c9;
               Y_3_c10 <= Y_3_c9;
               Y_4_c10 <= Y_4_c9;
               Y_5_c10 <= Y_5_c9;
               Y_6_c10 <= Y_6_c9;
               Y_7_c10 <= Y_7_c9;
               Y_8_c10 <= Y_8_c9;
               Y_9_c10 <= Y_9_c9;
               Y_10_c10 <= Y_10_c9;
               Y_11_c10 <= Y_11_c9;
            end if;
            if ce_11 = '1' then
               Y_1_c11 <= Y_1_c10;
               Y_2_c11 <= Y_2_c10;
               Y_3_c11 <= Y_3_c10;
               Y_4_c11 <= Y_4_c10;
               Y_5_c11 <= Y_5_c10;
               Y_6_c11 <= Y_6_c10;
               Y_7_c11 <= Y_7_c10;
               Y_8_c11 <= Y_8_c10;
               Y_9_c11 <= Y_9_c10;
               Y_10_c11 <= Y_10_c10;
               Y_11_c11 <= Y_11_c10;
            end if;
            if ce_12 = '1' then
               Y_1_c12 <= Y_1_c11;
               Y_2_c12 <= Y_2_c11;
               Y_3_c12 <= Y_3_c11;
               Y_4_c12 <= Y_4_c11;
               Y_5_c12 <= Y_5_c11;
               Y_6_c12 <= Y_6_c11;
               Y_7_c12 <= Y_7_c11;
               Y_8_c12 <= Y_8_c11;
               Y_9_c12 <= Y_9_c11;
               Y_10_c12 <= Y_10_c11;
               Y_11_c12 <= Y_11_c11;
            end if;
            if ce_13 = '1' then
               Y_1_c13 <= Y_1_c12;
               Y_2_c13 <= Y_2_c12;
               Y_3_c13 <= Y_3_c12;
               Y_4_c13 <= Y_4_c12;
               Y_5_c13 <= Y_5_c12;
               Y_6_c13 <= Y_6_c12;
               Y_7_c13 <= Y_7_c12;
               Y_8_c13 <= Y_8_c12;
               Y_9_c13 <= Y_9_c12;
               Y_10_c13 <= Y_10_c12;
               Y_11_c13 <= Y_11_c12;
            end if;
            if ce_14 = '1' then
               Y_1_c14 <= Y_1_c13;
               Y_2_c14 <= Y_2_c13;
               Y_3_c14 <= Y_3_c13;
               Y_4_c14 <= Y_4_c13;
               Y_5_c14 <= Y_5_c13;
               Y_6_c14 <= Y_6_c13;
               Y_7_c14 <= Y_7_c13;
               Y_8_c14 <= Y_8_c13;
               Y_9_c14 <= Y_9_c13;
               Y_10_c14 <= Y_10_c13;
               Y_11_c14 <= Y_11_c13;
            end if;
            if ce_15 = '1' then
               X_1_c15 <= X_1_c14;
               Y_1_c15 <= Y_1_c14;
               X_2_c15 <= X_2_c14;
               Y_2_c15 <= Y_2_c14;
               X_3_c15 <= X_3_c14;
               Y_3_c15 <= Y_3_c14;
               X_4_c15 <= X_4_c14;
               Y_4_c15 <= Y_4_c14;
               X_5_c15 <= X_5_c14;
               Y_5_c15 <= Y_5_c14;
               X_6_c15 <= X_6_c14;
               Y_6_c15 <= Y_6_c14;
               X_7_c15 <= X_7_c14;
               Y_7_c15 <= Y_7_c14;
               X_8_c15 <= X_8_c14;
               Y_8_c15 <= Y_8_c14;
               X_9_c15 <= X_9_c14;
               Y_9_c15 <= Y_9_c14;
               X_10_c15 <= X_10_c14;
               Y_10_c15 <= Y_10_c14;
               X_11_c15 <= X_11_c14;
               Y_11_c15 <= Y_11_c14;
            end if;
            if ce_16 = '1' then
               Cin_1_c16 <= Cin_1_c15;
               X_1_c16 <= X_1_c15;
               Y_1_c16 <= Y_1_c15;
               X_2_c16 <= X_2_c15;
               Y_2_c16 <= Y_2_c15;
               X_3_c16 <= X_3_c15;
               Y_3_c16 <= Y_3_c15;
               X_4_c16 <= X_4_c15;
               Y_4_c16 <= Y_4_c15;
               X_5_c16 <= X_5_c15;
               Y_5_c16 <= Y_5_c15;
               X_6_c16 <= X_6_c15;
               Y_6_c16 <= Y_6_c15;
               X_7_c16 <= X_7_c15;
               Y_7_c16 <= Y_7_c15;
               X_8_c16 <= X_8_c15;
               Y_8_c16 <= Y_8_c15;
               X_9_c16 <= X_9_c15;
               Y_9_c16 <= Y_9_c15;
               X_10_c16 <= X_10_c15;
               Y_10_c16 <= Y_10_c15;
               X_11_c16 <= X_11_c15;
               Y_11_c16 <= Y_11_c15;
            end if;
            if ce_17 = '1' then
               R_1_c17 <= R_1_c16;
               Cin_2_c17 <= Cin_2_c16;
               X_2_c17 <= X_2_c16;
               Y_2_c17 <= Y_2_c16;
               X_3_c17 <= X_3_c16;
               Y_3_c17 <= Y_3_c16;
               X_4_c17 <= X_4_c16;
               Y_4_c17 <= Y_4_c16;
               X_5_c17 <= X_5_c16;
               Y_5_c17 <= Y_5_c16;
               X_6_c17 <= X_6_c16;
               Y_6_c17 <= Y_6_c16;
               X_7_c17 <= X_7_c16;
               Y_7_c17 <= Y_7_c16;
               X_8_c17 <= X_8_c16;
               Y_8_c17 <= Y_8_c16;
               X_9_c17 <= X_9_c16;
               Y_9_c17 <= Y_9_c16;
               X_10_c17 <= X_10_c16;
               Y_10_c17 <= Y_10_c16;
               X_11_c17 <= X_11_c16;
               Y_11_c17 <= Y_11_c16;
            end if;
            if ce_18 = '1' then
               R_1_c18 <= R_1_c17;
               R_2_c18 <= R_2_c17;
               Cin_3_c18 <= Cin_3_c17;
               X_3_c18 <= X_3_c17;
               Y_3_c18 <= Y_3_c17;
               X_4_c18 <= X_4_c17;
               Y_4_c18 <= Y_4_c17;
               X_5_c18 <= X_5_c17;
               Y_5_c18 <= Y_5_c17;
               X_6_c18 <= X_6_c17;
               Y_6_c18 <= Y_6_c17;
               X_7_c18 <= X_7_c17;
               Y_7_c18 <= Y_7_c17;
               X_8_c18 <= X_8_c17;
               Y_8_c18 <= Y_8_c17;
               X_9_c18 <= X_9_c17;
               Y_9_c18 <= Y_9_c17;
               X_10_c18 <= X_10_c17;
               Y_10_c18 <= Y_10_c17;
               X_11_c18 <= X_11_c17;
               Y_11_c18 <= Y_11_c17;
            end if;
            if ce_19 = '1' then
               R_1_c19 <= R_1_c18;
               R_2_c19 <= R_2_c18;
               R_3_c19 <= R_3_c18;
               Cin_4_c19 <= Cin_4_c18;
               X_4_c19 <= X_4_c18;
               Y_4_c19 <= Y_4_c18;
               X_5_c19 <= X_5_c18;
               Y_5_c19 <= Y_5_c18;
               X_6_c19 <= X_6_c18;
               Y_6_c19 <= Y_6_c18;
               X_7_c19 <= X_7_c18;
               Y_7_c19 <= Y_7_c18;
               X_8_c19 <= X_8_c18;
               Y_8_c19 <= Y_8_c18;
               X_9_c19 <= X_9_c18;
               Y_9_c19 <= Y_9_c18;
               X_10_c19 <= X_10_c18;
               Y_10_c19 <= Y_10_c18;
               X_11_c19 <= X_11_c18;
               Y_11_c19 <= Y_11_c18;
            end if;
            if ce_20 = '1' then
               R_1_c20 <= R_1_c19;
               R_2_c20 <= R_2_c19;
               R_3_c20 <= R_3_c19;
               R_4_c20 <= R_4_c19;
               Cin_5_c20 <= Cin_5_c19;
               X_5_c20 <= X_5_c19;
               Y_5_c20 <= Y_5_c19;
               X_6_c20 <= X_6_c19;
               Y_6_c20 <= Y_6_c19;
               X_7_c20 <= X_7_c19;
               Y_7_c20 <= Y_7_c19;
               X_8_c20 <= X_8_c19;
               Y_8_c20 <= Y_8_c19;
               X_9_c20 <= X_9_c19;
               Y_9_c20 <= Y_9_c19;
               X_10_c20 <= X_10_c19;
               Y_10_c20 <= Y_10_c19;
               X_11_c20 <= X_11_c19;
               Y_11_c20 <= Y_11_c19;
            end if;
            if ce_21 = '1' then
               R_1_c21 <= R_1_c20;
               R_2_c21 <= R_2_c20;
               R_3_c21 <= R_3_c20;
               R_4_c21 <= R_4_c20;
               R_5_c21 <= R_5_c20;
               Cin_6_c21 <= Cin_6_c20;
               X_6_c21 <= X_6_c20;
               Y_6_c21 <= Y_6_c20;
               X_7_c21 <= X_7_c20;
               Y_7_c21 <= Y_7_c20;
               X_8_c21 <= X_8_c20;
               Y_8_c21 <= Y_8_c20;
               X_9_c21 <= X_9_c20;
               Y_9_c21 <= Y_9_c20;
               X_10_c21 <= X_10_c20;
               Y_10_c21 <= Y_10_c20;
               X_11_c21 <= X_11_c20;
               Y_11_c21 <= Y_11_c20;
            end if;
            if ce_22 = '1' then
               R_1_c22 <= R_1_c21;
               R_2_c22 <= R_2_c21;
               R_3_c22 <= R_3_c21;
               R_4_c22 <= R_4_c21;
               R_5_c22 <= R_5_c21;
               R_6_c22 <= R_6_c21;
               Cin_7_c22 <= Cin_7_c21;
               X_7_c22 <= X_7_c21;
               Y_7_c22 <= Y_7_c21;
               X_8_c22 <= X_8_c21;
               Y_8_c22 <= Y_8_c21;
               X_9_c22 <= X_9_c21;
               Y_9_c22 <= Y_9_c21;
               X_10_c22 <= X_10_c21;
               Y_10_c22 <= Y_10_c21;
               X_11_c22 <= X_11_c21;
               Y_11_c22 <= Y_11_c21;
            end if;
            if ce_23 = '1' then
               R_1_c23 <= R_1_c22;
               R_2_c23 <= R_2_c22;
               R_3_c23 <= R_3_c22;
               R_4_c23 <= R_4_c22;
               R_5_c23 <= R_5_c22;
               R_6_c23 <= R_6_c22;
               R_7_c23 <= R_7_c22;
               Cin_8_c23 <= Cin_8_c22;
               X_8_c23 <= X_8_c22;
               Y_8_c23 <= Y_8_c22;
               X_9_c23 <= X_9_c22;
               Y_9_c23 <= Y_9_c22;
               X_10_c23 <= X_10_c22;
               Y_10_c23 <= Y_10_c22;
               X_11_c23 <= X_11_c22;
               Y_11_c23 <= Y_11_c22;
            end if;
            if ce_24 = '1' then
               R_1_c24 <= R_1_c23;
               R_2_c24 <= R_2_c23;
               R_3_c24 <= R_3_c23;
               R_4_c24 <= R_4_c23;
               R_5_c24 <= R_5_c23;
               R_6_c24 <= R_6_c23;
               R_7_c24 <= R_7_c23;
               R_8_c24 <= R_8_c23;
               Cin_9_c24 <= Cin_9_c23;
               X_9_c24 <= X_9_c23;
               Y_9_c24 <= Y_9_c23;
               X_10_c24 <= X_10_c23;
               Y_10_c24 <= Y_10_c23;
               X_11_c24 <= X_11_c23;
               Y_11_c24 <= Y_11_c23;
            end if;
            if ce_25 = '1' then
               R_1_c25 <= R_1_c24;
               R_2_c25 <= R_2_c24;
               R_3_c25 <= R_3_c24;
               R_4_c25 <= R_4_c24;
               R_5_c25 <= R_5_c24;
               R_6_c25 <= R_6_c24;
               R_7_c25 <= R_7_c24;
               R_8_c25 <= R_8_c24;
               R_9_c25 <= R_9_c24;
               Cin_10_c25 <= Cin_10_c24;
               X_10_c25 <= X_10_c24;
               Y_10_c25 <= Y_10_c24;
               X_11_c25 <= X_11_c24;
               Y_11_c25 <= Y_11_c24;
            end if;
            if ce_26 = '1' then
               R_1_c26 <= R_1_c25;
               R_2_c26 <= R_2_c25;
               R_3_c26 <= R_3_c25;
               R_4_c26 <= R_4_c25;
               R_5_c26 <= R_5_c25;
               R_6_c26 <= R_6_c25;
               R_7_c26 <= R_7_c25;
               R_8_c26 <= R_8_c25;
               R_9_c26 <= R_9_c25;
               R_10_c26 <= R_10_c25;
               Cin_11_c26 <= Cin_11_c25;
               X_11_c26 <= X_11_c25;
               Y_11_c26 <= Y_11_c25;
            end if;
         end if;
      end process;
   Cin_1_c15 <= Cin;
   X_1_c14 <= '0' & X(2 downto 0);
   Y_1_c0 <= '0' & Y(2 downto 0);
   S_1_c16 <= X_1_c16 + Y_1_c16 + Cin_1_c16;
   R_1_c16 <= S_1_c16(2 downto 0);
   Cin_2_c16 <= S_1_c16(3);
   X_2_c14 <= '0' & X(5 downto 3);
   Y_2_c0 <= '0' & Y(5 downto 3);
   S_2_c17 <= X_2_c17 + Y_2_c17 + Cin_2_c17;
   R_2_c17 <= S_2_c17(2 downto 0);
   Cin_3_c17 <= S_2_c17(3);
   X_3_c14 <= '0' & X(8 downto 6);
   Y_3_c0 <= '0' & Y(8 downto 6);
   S_3_c18 <= X_3_c18 + Y_3_c18 + Cin_3_c18;
   R_3_c18 <= S_3_c18(2 downto 0);
   Cin_4_c18 <= S_3_c18(3);
   X_4_c14 <= '0' & X(11 downto 9);
   Y_4_c0 <= '0' & Y(11 downto 9);
   S_4_c19 <= X_4_c19 + Y_4_c19 + Cin_4_c19;
   R_4_c19 <= S_4_c19(2 downto 0);
   Cin_5_c19 <= S_4_c19(3);
   X_5_c14 <= '0' & X(14 downto 12);
   Y_5_c0 <= '0' & Y(14 downto 12);
   S_5_c20 <= X_5_c20 + Y_5_c20 + Cin_5_c20;
   R_5_c20 <= S_5_c20(2 downto 0);
   Cin_6_c20 <= S_5_c20(3);
   X_6_c14 <= '0' & X(17 downto 15);
   Y_6_c0 <= '0' & Y(17 downto 15);
   S_6_c21 <= X_6_c21 + Y_6_c21 + Cin_6_c21;
   R_6_c21 <= S_6_c21(2 downto 0);
   Cin_7_c21 <= S_6_c21(3);
   X_7_c14 <= '0' & X(20 downto 18);
   Y_7_c0 <= '0' & Y(20 downto 18);
   S_7_c22 <= X_7_c22 + Y_7_c22 + Cin_7_c22;
   R_7_c22 <= S_7_c22(2 downto 0);
   Cin_8_c22 <= S_7_c22(3);
   X_8_c14 <= '0' & X(23 downto 21);
   Y_8_c0 <= '0' & Y(23 downto 21);
   S_8_c23 <= X_8_c23 + Y_8_c23 + Cin_8_c23;
   R_8_c23 <= S_8_c23(2 downto 0);
   Cin_9_c23 <= S_8_c23(3);
   X_9_c14 <= '0' & X(26 downto 24);
   Y_9_c0 <= '0' & Y(26 downto 24);
   S_9_c24 <= X_9_c24 + Y_9_c24 + Cin_9_c24;
   R_9_c24 <= S_9_c24(2 downto 0);
   Cin_10_c24 <= S_9_c24(3);
   X_10_c14 <= '0' & X(29 downto 27);
   Y_10_c0 <= '0' & Y(29 downto 27);
   S_10_c25 <= X_10_c25 + Y_10_c25 + Cin_10_c25;
   R_10_c25 <= S_10_c25(2 downto 0);
   Cin_11_c25 <= S_10_c25(3);
   X_11_c14 <= '0' & X(32 downto 30);
   Y_11_c0 <= '0' & Y(32 downto 30);
   S_11_c26 <= X_11_c26 + Y_11_c26 + Cin_11_c26;
   R_11_c26 <= S_11_c26(2 downto 0);
   R <= R_11_c26 & R_10_c26 & R_9_c26 & R_8_c26 & R_7_c26 & R_6_c26 & R_5_c26 & R_4_c26 & R_3_c26 & R_2_c26 & R_1_c26 ;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointMultiplier
--                      (FPMult_8_23_uid2_Freq800_uid3)
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 26 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointMultiplier_32_2_034000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointMultiplier_32_2_034000 is
   component IntMultiplier_24x24_48_Freq800_uid5 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13 : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_Freq800_uid355 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26 : in std_logic;
             X : in  std_logic_vector(32 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(32 downto 0)   );
   end component;

signal sign_c0, sign_c1, sign_c2, sign_c3, sign_c4, sign_c5, sign_c6, sign_c7, sign_c8, sign_c9, sign_c10, sign_c11, sign_c12, sign_c13, sign_c14, sign_c15, sign_c16, sign_c17, sign_c18, sign_c19, sign_c20, sign_c21, sign_c22, sign_c23, sign_c24, sign_c25, sign_c26 :  std_logic;
signal expX_c0, expX_c1 :  std_logic_vector(7 downto 0);
signal expY_c0, expY_c1 :  std_logic_vector(7 downto 0);
signal expSumPreSub_c1, expSumPreSub_c2 :  std_logic_vector(9 downto 0);
signal bias_c0, bias_c1, bias_c2 :  std_logic_vector(9 downto 0);
signal expSum_c2, expSum_c3, expSum_c4, expSum_c5, expSum_c6, expSum_c7, expSum_c8, expSum_c9, expSum_c10, expSum_c11, expSum_c12, expSum_c13 :  std_logic_vector(9 downto 0);
signal sigX_c0 :  std_logic_vector(23 downto 0);
signal sigY_c0 :  std_logic_vector(23 downto 0);
signal sigProd_c13, sigProd_c14 :  std_logic_vector(47 downto 0);
signal excSel_c0 :  std_logic_vector(3 downto 0);
signal exc_c0, exc_c1, exc_c2, exc_c3, exc_c4, exc_c5, exc_c6, exc_c7, exc_c8, exc_c9, exc_c10, exc_c11, exc_c12, exc_c13, exc_c14, exc_c15, exc_c16, exc_c17, exc_c18, exc_c19, exc_c20, exc_c21, exc_c22, exc_c23, exc_c24, exc_c25, exc_c26 :  std_logic_vector(1 downto 0);
signal norm_c13, norm_c14 :  std_logic;
signal expPostNorm_c13, expPostNorm_c14 :  std_logic_vector(9 downto 0);
signal sigProdExt_c14, sigProdExt_c15 :  std_logic_vector(47 downto 0);
signal expSig_c14 :  std_logic_vector(32 downto 0);
signal sticky_c14, sticky_c15 :  std_logic;
signal guard_c14, guard_c15 :  std_logic;
signal round_c15 :  std_logic;
signal expSigPostRound_c26 :  std_logic_vector(32 downto 0);
signal excPostNorm_c26 :  std_logic_vector(1 downto 0);
signal finalExc_c26 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               sign_c1 <= sign_c0;
               expX_c1 <= expX_c0;
               expY_c1 <= expY_c0;
               bias_c1 <= bias_c0;
               exc_c1 <= exc_c0;
            end if;
            if ce_2 = '1' then
               sign_c2 <= sign_c1;
               expSumPreSub_c2 <= expSumPreSub_c1;
               bias_c2 <= bias_c1;
               exc_c2 <= exc_c1;
            end if;
            if ce_3 = '1' then
               sign_c3 <= sign_c2;
               expSum_c3 <= expSum_c2;
               exc_c3 <= exc_c2;
            end if;
            if ce_4 = '1' then
               sign_c4 <= sign_c3;
               expSum_c4 <= expSum_c3;
               exc_c4 <= exc_c3;
            end if;
            if ce_5 = '1' then
               sign_c5 <= sign_c4;
               expSum_c5 <= expSum_c4;
               exc_c5 <= exc_c4;
            end if;
            if ce_6 = '1' then
               sign_c6 <= sign_c5;
               expSum_c6 <= expSum_c5;
               exc_c6 <= exc_c5;
            end if;
            if ce_7 = '1' then
               sign_c7 <= sign_c6;
               expSum_c7 <= expSum_c6;
               exc_c7 <= exc_c6;
            end if;
            if ce_8 = '1' then
               sign_c8 <= sign_c7;
               expSum_c8 <= expSum_c7;
               exc_c8 <= exc_c7;
            end if;
            if ce_9 = '1' then
               sign_c9 <= sign_c8;
               expSum_c9 <= expSum_c8;
               exc_c9 <= exc_c8;
            end if;
            if ce_10 = '1' then
               sign_c10 <= sign_c9;
               expSum_c10 <= expSum_c9;
               exc_c10 <= exc_c9;
            end if;
            if ce_11 = '1' then
               sign_c11 <= sign_c10;
               expSum_c11 <= expSum_c10;
               exc_c11 <= exc_c10;
            end if;
            if ce_12 = '1' then
               sign_c12 <= sign_c11;
               expSum_c12 <= expSum_c11;
               exc_c12 <= exc_c11;
            end if;
            if ce_13 = '1' then
               sign_c13 <= sign_c12;
               expSum_c13 <= expSum_c12;
               exc_c13 <= exc_c12;
            end if;
            if ce_14 = '1' then
               sign_c14 <= sign_c13;
               sigProd_c14 <= sigProd_c13;
               exc_c14 <= exc_c13;
               norm_c14 <= norm_c13;
               expPostNorm_c14 <= expPostNorm_c13;
            end if;
            if ce_15 = '1' then
               sign_c15 <= sign_c14;
               exc_c15 <= exc_c14;
               sigProdExt_c15 <= sigProdExt_c14;
               sticky_c15 <= sticky_c14;
               guard_c15 <= guard_c14;
            end if;
            if ce_16 = '1' then
               sign_c16 <= sign_c15;
               exc_c16 <= exc_c15;
            end if;
            if ce_17 = '1' then
               sign_c17 <= sign_c16;
               exc_c17 <= exc_c16;
            end if;
            if ce_18 = '1' then
               sign_c18 <= sign_c17;
               exc_c18 <= exc_c17;
            end if;
            if ce_19 = '1' then
               sign_c19 <= sign_c18;
               exc_c19 <= exc_c18;
            end if;
            if ce_20 = '1' then
               sign_c20 <= sign_c19;
               exc_c20 <= exc_c19;
            end if;
            if ce_21 = '1' then
               sign_c21 <= sign_c20;
               exc_c21 <= exc_c20;
            end if;
            if ce_22 = '1' then
               sign_c22 <= sign_c21;
               exc_c22 <= exc_c21;
            end if;
            if ce_23 = '1' then
               sign_c23 <= sign_c22;
               exc_c23 <= exc_c22;
            end if;
            if ce_24 = '1' then
               sign_c24 <= sign_c23;
               exc_c24 <= exc_c23;
            end if;
            if ce_25 = '1' then
               sign_c25 <= sign_c24;
               exc_c25 <= exc_c24;
            end if;
            if ce_26 = '1' then
               sign_c26 <= sign_c25;
               exc_c26 <= exc_c25;
            end if;
         end if;
      end process;
   sign_c0 <= X(31) xor Y(31);
   expX_c0 <= X(30 downto 23);
   expY_c0 <= Y(30 downto 23);
   expSumPreSub_c1 <= ("00" & expX_c1) + ("00" & expY_c1);
   bias_c0 <= CONV_STD_LOGIC_VECTOR(127,10);
   expSum_c2 <= expSumPreSub_c2 - bias_c2;
   sigX_c0 <= "1" & X(22 downto 0);
   sigY_c0 <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_24x24_48_Freq800_uid5
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 X => sigX_c0,
                 Y => sigY_c0,
                 R => sigProd_c13);
   excSel_c0 <= X(33 downto 32) & Y(33 downto 32);
   with excSel_c0  select  
   exc_c0 <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm_c13 <= sigProd_c13(47);
   -- exponent update
   expPostNorm_c13 <= expSum_c13 + ("000000000" & norm_c13);
   -- significand normalization shift
   sigProdExt_c14 <= sigProd_c14(46 downto 0) & "0" when norm_c14='1' else
                         sigProd_c14(45 downto 0) & "00";
   expSig_c14 <= expPostNorm_c14 & sigProdExt_c14(47 downto 25);
   sticky_c14 <= sigProdExt_c14(24);
   guard_c14 <= '0' when sigProdExt_c14(23 downto 0)="000000000000000000000000" else '1';
   round_c15 <= sticky_c15 and ( (guard_c15 and not(sigProdExt_c15(25))) or (sigProdExt_c15(25) ))  ;
   RoundingAdder: IntAdder_33_Freq800_uid355
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 Cin => round_c15,
                 X => expSig_c14,
                 Y => "000000000000000000000000000000000",
                 R => expSigPostRound_c26);
   with expSigPostRound_c26(32 downto 31)  select 
   excPostNorm_c26 <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_c26  select  
   finalExc_c26 <= exc_c26 when  "11"|"10"|"00",
                       excPostNorm_c26 when others; 
   R <= finalExc_c26 & sign_c26 & expSigPostRound_c26(30 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid15
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid15 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid15 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid20
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid20 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid20 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid27
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid27 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid27 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid32
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid32 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid32 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid39
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid39 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid39 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid44
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid44 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid44 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid51
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid51 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid51 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid56
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid56 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid56 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid63
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid63 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid63 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid68
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid68 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid68 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid75
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid75 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid75 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid80
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid80 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid80 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid87
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid87 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid87 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid92
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid92 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid92 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid99
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid99 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid99 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid104
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid104 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid104 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid111
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid111 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid111 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid116
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid116 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid116 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid123
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid128
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid128 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid128 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid135
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid135 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid135 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid140
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid140 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid140 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid147
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid147 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid147 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid152
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid152 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid152 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq500_uid156
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq500_uid156 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq500_uid156 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq500_uid160
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq500_uid160 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq500_uid160 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq500_uid164
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq500_uid164 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq500_uid164 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq500_uid170
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq500_uid170 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq500_uid170 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq500_uid9
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq500_uid9 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq500_uid9 is
signal Mfull_c0, Mfull_c1 :  std_logic_vector(40 downto 0);
signal M_c1 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c1 <= Mfull_c1(40 downto 0);
   R <= M_c1;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq500_uid11
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid11 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid11 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid13
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid13 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid13 is
   component MultTable_Freq500_uid15 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy16_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid15
      port map ( X => Xtable_c0,
                 Y => Y1_copy16_c0);
   Y1_c0 <= Y1_copy16_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid18
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid18 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid18 is
   component MultTable_Freq500_uid20 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy21_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid20
      port map ( X => Xtable_c0,
                 Y => Y1_copy21_c0);
   Y1_c0 <= Y1_copy21_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq500_uid23
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid23 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid23 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid25
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid25 is
   component MultTable_Freq500_uid27 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy28_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid27
      port map ( X => Xtable_c0,
                 Y => Y1_copy28_c0);
   Y1_c0 <= Y1_copy28_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid30
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid30 is
   component MultTable_Freq500_uid32 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy33_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid32
      port map ( X => Xtable_c0,
                 Y => Y1_copy33_c0);
   Y1_c0 <= Y1_copy33_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq500_uid35
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid35 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid35 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid37
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid37 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid37 is
   component MultTable_Freq500_uid39 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy40_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid39
      port map ( X => Xtable_c0,
                 Y => Y1_copy40_c0);
   Y1_c0 <= Y1_copy40_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid42
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid42 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid42 is
   component MultTable_Freq500_uid44 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy45_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid44
      port map ( X => Xtable_c0,
                 Y => Y1_copy45_c0);
   Y1_c0 <= Y1_copy45_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq500_uid47
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid47 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid47 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid49
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid49 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid49 is
   component MultTable_Freq500_uid51 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy52_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid51
      port map ( X => Xtable_c0,
                 Y => Y1_copy52_c0);
   Y1_c0 <= Y1_copy52_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid54
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid54 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid54 is
   component MultTable_Freq500_uid56 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy57_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid56
      port map ( X => Xtable_c0,
                 Y => Y1_copy57_c0);
   Y1_c0 <= Y1_copy57_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq500_uid59
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid59 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid59 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid61
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid61 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid61 is
   component MultTable_Freq500_uid63 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy64_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid63
      port map ( X => Xtable_c0,
                 Y => Y1_copy64_c0);
   Y1_c0 <= Y1_copy64_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid66
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid66 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid66 is
   component MultTable_Freq500_uid68 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy69_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid68
      port map ( X => Xtable_c0,
                 Y => Y1_copy69_c0);
   Y1_c0 <= Y1_copy69_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq500_uid71
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid71 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid73
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid73 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid73 is
   component MultTable_Freq500_uid75 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy76_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid75
      port map ( X => Xtable_c0,
                 Y => Y1_copy76_c0);
   Y1_c0 <= Y1_copy76_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid78
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid78 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid78 is
   component MultTable_Freq500_uid80 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy81_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid80
      port map ( X => Xtable_c0,
                 Y => Y1_copy81_c0);
   Y1_c0 <= Y1_copy81_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq500_uid83
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid83 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid83 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid85
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid85 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid85 is
   component MultTable_Freq500_uid87 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy88_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid87
      port map ( X => Xtable_c0,
                 Y => Y1_copy88_c0);
   Y1_c0 <= Y1_copy88_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid90
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid90 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid90 is
   component MultTable_Freq500_uid92 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy93_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid92
      port map ( X => Xtable_c0,
                 Y => Y1_copy93_c0);
   Y1_c0 <= Y1_copy93_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq500_uid95
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid95 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid95 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq500_uid97
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid97 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid97 is
   component MultTable_Freq500_uid99 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy100_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid99
      port map ( X => Xtable_c0,
                 Y => Y1_copy100_c0);
   Y1_c0 <= Y1_copy100_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid102
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid102 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid102 is
   component MultTable_Freq500_uid104 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy105_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid104
      port map ( X => Xtable_c0,
                 Y => Y1_copy105_c0);
   Y1_c0 <= Y1_copy105_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq500_uid107
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid107 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid107 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid109
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid109 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid109 is
   component MultTable_Freq500_uid111 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy112_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid111
      port map ( X => Xtable_c0,
                 Y => Y1_copy112_c0);
   Y1_c0 <= Y1_copy112_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid114
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid114 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid114 is
   component MultTable_Freq500_uid116 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy117_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid116
      port map ( X => Xtable_c0,
                 Y => Y1_copy117_c0);
   Y1_c0 <= Y1_copy117_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq500_uid119
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid119 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid119 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid121
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid121 is
   component MultTable_Freq500_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy124_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid123
      port map ( X => Xtable_c0,
                 Y => Y1_copy124_c0);
   Y1_c0 <= Y1_copy124_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid126
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid126 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid126 is
   component MultTable_Freq500_uid128 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy129_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid128
      port map ( X => Xtable_c0,
                 Y => Y1_copy129_c0);
   Y1_c0 <= Y1_copy129_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq500_uid131
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid131 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid131 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid133
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid133 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid133 is
   component MultTable_Freq500_uid135 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy136_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid135
      port map ( X => Xtable_c0,
                 Y => Y1_copy136_c0);
   Y1_c0 <= Y1_copy136_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid138
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid138 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid138 is
   component MultTable_Freq500_uid140 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy141_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid140
      port map ( X => Xtable_c0,
                 Y => Y1_copy141_c0);
   Y1_c0 <= Y1_copy141_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq500_uid143
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq500_uid143 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq500_uid143 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid145
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid145 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid145 is
   component MultTable_Freq500_uid147 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy148_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid147
      port map ( X => Xtable_c0,
                 Y => Y1_copy148_c0);
   Y1_c0 <= Y1_copy148_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid150
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid150 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid150 is
   component MultTable_Freq500_uid152 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy153_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid152
      port map ( X => Xtable_c0,
                 Y => Y1_copy153_c0);
   Y1_c0 <= Y1_copy153_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_30_Freq500_uid330
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_30_Freq500_uid330 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(29 downto 0);
          Y : in  std_logic_vector(29 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of IntAdder_30_Freq500_uid330 is
signal Rtmp_c2 :  std_logic_vector(29 downto 0);
signal X_c2 :  std_logic_vector(29 downto 0);
signal Y_c2 :  std_logic_vector(29 downto 0);
signal Cin_c1, Cin_c2 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               X_c2 <= X;
               Y_c2 <= Y;
               Cin_c2 <= Cin_c1;
            end if;
         end if;
      end process;
   Rtmp_c2 <= X_c2 + Y_c2 + Cin_c2;
   R <= Rtmp_c2;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_24x24_48_Freq500_uid5
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_24x24_48_Freq500_uid5 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_24x24_48_Freq500_uid5 is
   component DSPBlock_17x24_Freq500_uid9 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid11 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid13 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid18 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid23 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid35 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid37 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid42 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid47 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid49 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid54 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid59 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid61 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid66 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid73 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid78 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid83 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid85 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid90 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid95 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid97 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid102 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid107 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid109 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid114 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid119 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid126 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid131 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid133 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid138 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq500_uid143 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid145 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid150 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq500_uid156 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq500_uid160 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_14_3_Freq500_uid164 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq500_uid170 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_30_Freq500_uid330 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(29 downto 0);
             Y : in  std_logic_vector(29 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(29 downto 0)   );
   end component;

signal XX_m6_c0 :  std_logic_vector(23 downto 0);
signal YY_m6_c0 :  std_logic_vector(23 downto 0);
signal tile_0_X_c0 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_0_output_c1 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c1 :  unsigned(40-0 downto 0);
signal bh7_w0_0_c1 :  std_logic;
signal bh7_w1_0_c1 :  std_logic;
signal bh7_w2_0_c1 :  std_logic;
signal bh7_w3_0_c1 :  std_logic;
signal bh7_w4_0_c1 :  std_logic;
signal bh7_w5_0_c1 :  std_logic;
signal bh7_w6_0_c1 :  std_logic;
signal bh7_w7_0_c1 :  std_logic;
signal bh7_w8_0_c1 :  std_logic;
signal bh7_w9_0_c1 :  std_logic;
signal bh7_w10_0_c1 :  std_logic;
signal bh7_w11_0_c1 :  std_logic;
signal bh7_w12_0_c1 :  std_logic;
signal bh7_w13_0_c1 :  std_logic;
signal bh7_w14_0_c1 :  std_logic;
signal bh7_w15_0_c1 :  std_logic;
signal bh7_w16_0_c1 :  std_logic;
signal bh7_w17_0_c1 :  std_logic;
signal bh7_w18_0_c1 :  std_logic;
signal bh7_w19_0_c1 :  std_logic;
signal bh7_w20_0_c1 :  std_logic;
signal bh7_w21_0_c1 :  std_logic;
signal bh7_w22_0_c1 :  std_logic;
signal bh7_w23_0_c1 :  std_logic;
signal bh7_w24_0_c1 :  std_logic;
signal bh7_w25_0_c1 :  std_logic;
signal bh7_w26_0_c1 :  std_logic;
signal bh7_w27_0_c1 :  std_logic;
signal bh7_w28_0_c1 :  std_logic;
signal bh7_w29_0_c1 :  std_logic;
signal bh7_w30_0_c1 :  std_logic;
signal bh7_w31_0_c1 :  std_logic;
signal bh7_w32_0_c1 :  std_logic;
signal bh7_w33_0_c1 :  std_logic;
signal bh7_w34_0_c1 :  std_logic;
signal bh7_w35_0_c1 :  std_logic;
signal bh7_w36_0_c1 :  std_logic;
signal bh7_w37_0_c1 :  std_logic;
signal bh7_w38_0_c1 :  std_logic;
signal bh7_w39_0_c1 :  std_logic;
signal bh7_w40_0_c1 :  std_logic;
signal tile_1_X_c0 :  std_logic_vector(0 downto 0);
signal tile_1_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_1_output_c0 :  std_logic_vector(1 downto 0);
signal tile_1_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w45_0_c0 :  std_logic;
signal bh7_w46_0_c0 :  std_logic;
signal tile_2_X_c0 :  std_logic_vector(2 downto 0);
signal tile_2_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_2_output_c0 :  std_logic_vector(4 downto 0);
signal tile_2_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w42_0_c0 :  std_logic;
signal bh7_w43_0_c0 :  std_logic;
signal bh7_w44_0_c0 :  std_logic;
signal bh7_w45_1_c0 :  std_logic;
signal bh7_w46_1_c0 :  std_logic;
signal tile_3_X_c0 :  std_logic_vector(2 downto 0);
signal tile_3_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_3_output_c0 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w39_1_c0 :  std_logic;
signal bh7_w40_1_c0 :  std_logic;
signal bh7_w41_0_c0 :  std_logic;
signal bh7_w42_1_c0 :  std_logic;
signal bh7_w43_1_c0 :  std_logic;
signal tile_4_X_c0 :  std_logic_vector(0 downto 0);
signal tile_4_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_4_output_c0 :  std_logic_vector(1 downto 0);
signal tile_4_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w43_2_c0 :  std_logic;
signal bh7_w44_1_c0 :  std_logic;
signal tile_5_X_c0 :  std_logic_vector(2 downto 0);
signal tile_5_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_5_output_c0 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w40_2_c0 :  std_logic;
signal bh7_w41_1_c0 :  std_logic;
signal bh7_w42_2_c0 :  std_logic;
signal bh7_w43_3_c0 :  std_logic;
signal bh7_w44_2_c0 :  std_logic;
signal tile_6_X_c0 :  std_logic_vector(2 downto 0);
signal tile_6_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_6_output_c0 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w37_1_c0 :  std_logic;
signal bh7_w38_1_c0 :  std_logic;
signal bh7_w39_2_c0 :  std_logic;
signal bh7_w40_3_c0 :  std_logic;
signal bh7_w41_2_c0 :  std_logic;
signal tile_7_X_c0 :  std_logic_vector(0 downto 0);
signal tile_7_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_7_output_c0 :  std_logic_vector(1 downto 0);
signal tile_7_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w41_3_c0 :  std_logic;
signal bh7_w42_3_c0 :  std_logic;
signal tile_8_X_c0 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_8_output_c0 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w38_2_c0 :  std_logic;
signal bh7_w39_3_c0 :  std_logic;
signal bh7_w40_4_c0 :  std_logic;
signal bh7_w41_4_c0 :  std_logic;
signal bh7_w42_4_c0 :  std_logic;
signal tile_9_X_c0 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_9_output_c0 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w35_1_c0 :  std_logic;
signal bh7_w36_1_c0 :  std_logic;
signal bh7_w37_2_c0 :  std_logic;
signal bh7_w38_3_c0 :  std_logic;
signal bh7_w39_4_c0 :  std_logic;
signal tile_10_X_c0 :  std_logic_vector(0 downto 0);
signal tile_10_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_10_output_c0 :  std_logic_vector(1 downto 0);
signal tile_10_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w39_5_c0 :  std_logic;
signal bh7_w40_5_c0 :  std_logic;
signal tile_11_X_c0 :  std_logic_vector(2 downto 0);
signal tile_11_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_11_output_c0 :  std_logic_vector(4 downto 0);
signal tile_11_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w36_2_c0 :  std_logic;
signal bh7_w37_3_c0 :  std_logic;
signal bh7_w38_4_c0 :  std_logic;
signal bh7_w39_6_c0 :  std_logic;
signal bh7_w40_6_c0 :  std_logic;
signal tile_12_X_c0 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_12_output_c0 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w33_1_c0 :  std_logic;
signal bh7_w34_1_c0 :  std_logic;
signal bh7_w35_2_c0 :  std_logic;
signal bh7_w36_3_c0 :  std_logic;
signal bh7_w37_4_c0 :  std_logic;
signal tile_13_X_c0 :  std_logic_vector(0 downto 0);
signal tile_13_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_13_output_c0 :  std_logic_vector(1 downto 0);
signal tile_13_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w37_5_c0 :  std_logic;
signal bh7_w38_5_c0 :  std_logic;
signal tile_14_X_c0 :  std_logic_vector(2 downto 0);
signal tile_14_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_14_output_c0 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w34_2_c0 :  std_logic;
signal bh7_w35_3_c0 :  std_logic;
signal bh7_w36_4_c0 :  std_logic;
signal bh7_w37_6_c0 :  std_logic;
signal bh7_w38_6_c0 :  std_logic;
signal tile_15_X_c0 :  std_logic_vector(2 downto 0);
signal tile_15_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_15_output_c0 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w31_1_c0 :  std_logic;
signal bh7_w32_1_c0 :  std_logic;
signal bh7_w33_2_c0 :  std_logic;
signal bh7_w34_3_c0 :  std_logic;
signal bh7_w35_4_c0 :  std_logic;
signal tile_16_X_c0 :  std_logic_vector(0 downto 0);
signal tile_16_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_16_output_c0 :  std_logic_vector(1 downto 0);
signal tile_16_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w35_5_c0 :  std_logic;
signal bh7_w36_5_c0 :  std_logic;
signal tile_17_X_c0 :  std_logic_vector(2 downto 0);
signal tile_17_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_17_output_c0 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w32_2_c0 :  std_logic;
signal bh7_w33_3_c0 :  std_logic;
signal bh7_w34_4_c0 :  std_logic;
signal bh7_w35_6_c0 :  std_logic;
signal bh7_w36_6_c0 :  std_logic;
signal tile_18_X_c0 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_18_output_c0 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w29_1_c0 :  std_logic;
signal bh7_w30_1_c0 :  std_logic;
signal bh7_w31_2_c0 :  std_logic;
signal bh7_w32_3_c0 :  std_logic;
signal bh7_w33_4_c0 :  std_logic;
signal tile_19_X_c0 :  std_logic_vector(0 downto 0);
signal tile_19_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_19_output_c0 :  std_logic_vector(1 downto 0);
signal tile_19_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w33_5_c0 :  std_logic;
signal bh7_w34_5_c0 :  std_logic;
signal tile_20_X_c0 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_20_output_c0 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w30_2_c0 :  std_logic;
signal bh7_w31_3_c0 :  std_logic;
signal bh7_w32_4_c0 :  std_logic;
signal bh7_w33_6_c0 :  std_logic;
signal bh7_w34_6_c0 :  std_logic;
signal tile_21_X_c0 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_21_output_c0 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w27_1_c0 :  std_logic;
signal bh7_w28_1_c0 :  std_logic;
signal bh7_w29_2_c0 :  std_logic;
signal bh7_w30_3_c0 :  std_logic;
signal bh7_w31_4_c0 :  std_logic;
signal tile_22_X_c0 :  std_logic_vector(0 downto 0);
signal tile_22_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_22_output_c0 :  std_logic_vector(1 downto 0);
signal tile_22_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w31_5_c0 :  std_logic;
signal bh7_w32_5_c0 :  std_logic;
signal tile_23_X_c0 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_23_output_c0 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w28_2_c0 :  std_logic;
signal bh7_w29_3_c0 :  std_logic;
signal bh7_w30_4_c0 :  std_logic;
signal bh7_w31_6_c0 :  std_logic;
signal bh7_w32_6_c0 :  std_logic;
signal tile_24_X_c0 :  std_logic_vector(2 downto 0);
signal tile_24_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_24_output_c0 :  std_logic_vector(4 downto 0);
signal tile_24_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w25_1_c0 :  std_logic;
signal bh7_w26_1_c0 :  std_logic;
signal bh7_w27_2_c0 :  std_logic;
signal bh7_w28_3_c0 :  std_logic;
signal bh7_w29_4_c0 :  std_logic;
signal tile_25_X_c0 :  std_logic_vector(0 downto 0);
signal tile_25_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_25_output_c0 :  std_logic_vector(1 downto 0);
signal tile_25_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w29_5_c0 :  std_logic;
signal bh7_w30_5_c0 :  std_logic;
signal tile_26_X_c0 :  std_logic_vector(2 downto 0);
signal tile_26_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_26_output_c0 :  std_logic_vector(4 downto 0);
signal tile_26_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w26_2_c0 :  std_logic;
signal bh7_w27_3_c0 :  std_logic;
signal bh7_w28_4_c0 :  std_logic;
signal bh7_w29_6_c0 :  std_logic;
signal bh7_w30_6_c0 :  std_logic;
signal tile_27_X_c0 :  std_logic_vector(2 downto 0);
signal tile_27_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_27_output_c0 :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w23_1_c0 :  std_logic;
signal bh7_w24_1_c0 :  std_logic;
signal bh7_w25_2_c0 :  std_logic;
signal bh7_w26_3_c0 :  std_logic;
signal bh7_w27_4_c0 :  std_logic;
signal tile_28_X_c0 :  std_logic_vector(0 downto 0);
signal tile_28_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_28_output_c0 :  std_logic_vector(1 downto 0);
signal tile_28_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w27_5_c0 :  std_logic;
signal bh7_w28_5_c0 :  std_logic;
signal tile_29_X_c0 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_29_output_c0 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w24_2_c0 :  std_logic;
signal bh7_w25_3_c0 :  std_logic;
signal bh7_w26_4_c0 :  std_logic;
signal bh7_w27_6_c0 :  std_logic;
signal bh7_w28_6_c0 :  std_logic;
signal tile_30_X_c0 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_30_output_c0 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w21_1_c0 :  std_logic;
signal bh7_w22_1_c0 :  std_logic;
signal bh7_w23_2_c0 :  std_logic;
signal bh7_w24_3_c0 :  std_logic;
signal bh7_w25_4_c0 :  std_logic;
signal tile_31_X_c0 :  std_logic_vector(0 downto 0);
signal tile_31_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_31_output_c0 :  std_logic_vector(1 downto 0);
signal tile_31_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w25_5_c0 :  std_logic;
signal bh7_w26_5_c0 :  std_logic;
signal tile_32_X_c0 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_32_output_c0 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w22_2_c0 :  std_logic;
signal bh7_w23_3_c0 :  std_logic;
signal bh7_w24_4_c0 :  std_logic;
signal bh7_w25_6_c0 :  std_logic;
signal bh7_w26_6_c0 :  std_logic;
signal tile_33_X_c0 :  std_logic_vector(2 downto 0);
signal tile_33_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_33_output_c0 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w19_1_c0 :  std_logic;
signal bh7_w20_1_c0 :  std_logic;
signal bh7_w21_2_c0 :  std_logic;
signal bh7_w22_3_c0 :  std_logic;
signal bh7_w23_4_c0 :  std_logic;
signal tile_34_X_c0 :  std_logic_vector(0 downto 0);
signal tile_34_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_34_output_c0 :  std_logic_vector(1 downto 0);
signal tile_34_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w23_5_c0 :  std_logic;
signal bh7_w24_5_c0 :  std_logic;
signal tile_35_X_c0 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_35_output_c0 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w20_2_c0 :  std_logic;
signal bh7_w21_3_c0 :  std_logic;
signal bh7_w22_4_c0 :  std_logic;
signal bh7_w23_6_c0 :  std_logic;
signal bh7_w24_6_c0 :  std_logic;
signal tile_36_X_c0 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_36_output_c0 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w17_1_c0, bh7_w17_1_c1 :  std_logic;
signal bh7_w18_1_c0 :  std_logic;
signal bh7_w19_2_c0 :  std_logic;
signal bh7_w20_3_c0 :  std_logic;
signal bh7_w21_4_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid157_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid157_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid157_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w18_2_c0, bh7_w18_2_c1 :  std_logic;
signal bh7_w19_3_c0, bh7_w19_3_c1 :  std_logic;
signal bh7_w20_4_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid157_Out0_copy158_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid161_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid161_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w20_5_c0 :  std_logic;
signal bh7_w21_5_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid160_bh7_uid161_Out0_copy162_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid165_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid165_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid165_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w21_6_c0 :  std_logic;
signal bh7_w22_5_c0 :  std_logic;
signal bh7_w23_7_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid165_Out0_copy166_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid167_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid167_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w22_6_c0 :  std_logic;
signal bh7_w23_8_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid160_bh7_uid167_Out0_copy168_c0 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid171_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid171_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w23_9_c0 :  std_logic;
signal bh7_w24_7_c0 :  std_logic;
signal bh7_w25_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid171_Out0_copy172_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid173_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid173_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w24_8_c0 :  std_logic;
signal bh7_w25_8_c0 :  std_logic;
signal bh7_w26_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid173_Out0_copy174_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid175_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid175_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w25_9_c0 :  std_logic;
signal bh7_w26_8_c0 :  std_logic;
signal bh7_w27_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid175_Out0_copy176_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid177_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid177_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w26_9_c0 :  std_logic;
signal bh7_w27_8_c0 :  std_logic;
signal bh7_w28_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid177_Out0_copy178_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid179_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid179_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w27_9_c0 :  std_logic;
signal bh7_w28_8_c0 :  std_logic;
signal bh7_w29_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid179_Out0_copy180_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid181_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid181_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w28_9_c0 :  std_logic;
signal bh7_w29_8_c0 :  std_logic;
signal bh7_w30_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid181_Out0_copy182_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid183_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid183_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w29_9_c0 :  std_logic;
signal bh7_w30_8_c0 :  std_logic;
signal bh7_w31_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid183_Out0_copy184_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid185_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid185_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w30_9_c0 :  std_logic;
signal bh7_w31_8_c0 :  std_logic;
signal bh7_w32_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid185_Out0_copy186_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid187_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid187_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w31_9_c0 :  std_logic;
signal bh7_w32_8_c0 :  std_logic;
signal bh7_w33_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid187_Out0_copy188_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid189_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid189_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w32_9_c0 :  std_logic;
signal bh7_w33_8_c0 :  std_logic;
signal bh7_w34_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid189_Out0_copy190_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid191_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid191_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w33_9_c0 :  std_logic;
signal bh7_w34_8_c0 :  std_logic;
signal bh7_w35_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid191_Out0_copy192_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid193_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid193_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w34_9_c0 :  std_logic;
signal bh7_w35_8_c0 :  std_logic;
signal bh7_w36_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid193_Out0_copy194_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid195_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid195_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w35_9_c0 :  std_logic;
signal bh7_w36_8_c0 :  std_logic;
signal bh7_w37_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid195_Out0_copy196_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid197_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid197_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w36_9_c0 :  std_logic;
signal bh7_w37_8_c0 :  std_logic;
signal bh7_w38_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid197_Out0_copy198_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid199_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid199_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w37_9_c0 :  std_logic;
signal bh7_w38_8_c0 :  std_logic;
signal bh7_w39_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid199_Out0_copy200_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid201_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid201_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w38_9_c0 :  std_logic;
signal bh7_w39_8_c0 :  std_logic;
signal bh7_w40_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid201_Out0_copy202_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid203_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid203_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w39_9_c0 :  std_logic;
signal bh7_w40_8_c0 :  std_logic;
signal bh7_w41_5_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid203_Out0_copy204_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid205_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid170_bh7_uid205_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w40_9_c0 :  std_logic;
signal bh7_w41_6_c0 :  std_logic;
signal bh7_w42_5_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid170_bh7_uid205_Out0_copy206_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid207_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid207_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid207_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w41_7_c0 :  std_logic;
signal bh7_w42_6_c0 :  std_logic;
signal bh7_w43_4_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid207_Out0_copy208_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid209_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid209_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid209_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w42_7_c0 :  std_logic;
signal bh7_w43_5_c0 :  std_logic;
signal bh7_w44_3_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid209_Out0_copy210_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid211_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid211_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid211_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w43_6_c0 :  std_logic;
signal bh7_w44_4_c0 :  std_logic;
signal bh7_w45_2_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid211_Out0_copy212_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid213_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid213_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid213_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w45_3_c0 :  std_logic;
signal bh7_w46_2_c0 :  std_logic;
signal bh7_w47_0_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid213_Out0_copy214_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid215_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid215_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid215_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w20_6_c0, bh7_w20_6_c1 :  std_logic;
signal bh7_w21_7_c0, bh7_w21_7_c1 :  std_logic;
signal bh7_w22_7_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid215_Out0_copy216_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid217_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid217_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w22_8_c0 :  std_logic;
signal bh7_w23_10_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid160_bh7_uid217_Out0_copy218_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid219_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid219_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid219_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w23_11_c0 :  std_logic;
signal bh7_w24_9_c0, bh7_w24_9_c1 :  std_logic;
signal bh7_w25_10_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid219_Out0_copy220_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid221_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid221_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid221_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w25_11_c0 :  std_logic;
signal bh7_w26_10_c0 :  std_logic;
signal bh7_w27_10_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid221_Out0_copy222_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid223_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid223_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid223_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w27_11_c0 :  std_logic;
signal bh7_w28_10_c0 :  std_logic;
signal bh7_w29_10_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid223_Out0_copy224_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid225_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid225_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid225_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w29_11_c0 :  std_logic;
signal bh7_w30_10_c0 :  std_logic;
signal bh7_w31_10_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid225_Out0_copy226_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid227_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid227_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid227_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w31_11_c0 :  std_logic;
signal bh7_w32_10_c0 :  std_logic;
signal bh7_w33_10_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid227_Out0_copy228_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid229_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid229_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid229_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w33_11_c0 :  std_logic;
signal bh7_w34_10_c0 :  std_logic;
signal bh7_w35_10_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid229_Out0_copy230_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid231_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid231_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid231_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w35_11_c0 :  std_logic;
signal bh7_w36_10_c0 :  std_logic;
signal bh7_w37_10_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid231_Out0_copy232_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid233_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid233_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid233_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w37_11_c0 :  std_logic;
signal bh7_w38_10_c0 :  std_logic;
signal bh7_w39_10_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid233_Out0_copy234_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid235_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid235_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid235_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w39_11_c0 :  std_logic;
signal bh7_w40_10_c0 :  std_logic;
signal bh7_w41_8_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid235_Out0_copy236_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid237_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid237_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid237_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w41_9_c0 :  std_logic;
signal bh7_w42_8_c0 :  std_logic;
signal bh7_w43_7_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid237_Out0_copy238_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid239_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid239_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w42_9_c0 :  std_logic;
signal bh7_w43_8_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid160_bh7_uid239_Out0_copy240_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid241_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid241_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid241_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w43_9_c0 :  std_logic;
signal bh7_w44_5_c0 :  std_logic;
signal bh7_w45_4_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid241_Out0_copy242_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid243_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid243_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid243_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w45_5_c0 :  std_logic;
signal bh7_w46_3_c0 :  std_logic;
signal bh7_w47_1_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid243_Out0_copy244_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid245_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid245_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w22_9_c1 :  std_logic;
signal bh7_w23_12_c1 :  std_logic;
signal bh7_w24_10_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_copy246_c0, Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_copy246_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid247_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid247_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w25_12_c1 :  std_logic;
signal bh7_w26_11_c1 :  std_logic;
signal bh7_w27_12_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_copy248_c0, Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_copy248_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid249_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid249_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w27_13_c1 :  std_logic;
signal bh7_w28_11_c1 :  std_logic;
signal bh7_w29_12_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_copy250_c0, Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_copy250_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid251_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid251_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_13_c1 :  std_logic;
signal bh7_w30_11_c1 :  std_logic;
signal bh7_w31_12_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_copy252_c0, Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_copy252_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid253_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid253_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_13_c1 :  std_logic;
signal bh7_w32_11_c1 :  std_logic;
signal bh7_w33_12_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_copy254_c0, Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_copy254_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid255_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid255_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_13_c1 :  std_logic;
signal bh7_w34_11_c1 :  std_logic;
signal bh7_w35_12_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_copy256_c0, Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_copy256_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid257_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid257_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w35_13_c1 :  std_logic;
signal bh7_w36_11_c1 :  std_logic;
signal bh7_w37_12_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_copy258_c0, Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_copy258_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid259_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid259_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w37_13_c1 :  std_logic;
signal bh7_w38_11_c1 :  std_logic;
signal bh7_w39_12_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_copy260_c0, Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_copy260_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid261_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid261_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w39_13_c1 :  std_logic;
signal bh7_w40_11_c1 :  std_logic;
signal bh7_w41_10_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_copy262_c0, Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_copy262_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid263_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid263_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w41_11_c1 :  std_logic;
signal bh7_w42_10_c1 :  std_logic;
signal bh7_w43_10_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_copy264_c0, Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_copy264_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid265_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid265_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w43_11_c1 :  std_logic;
signal bh7_w44_6_c1 :  std_logic;
signal bh7_w45_6_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_copy266_c0, Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_copy266_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid267_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid267_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w45_7_c1 :  std_logic;
signal bh7_w46_4_c1 :  std_logic;
signal bh7_w47_2_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_copy268_c0, Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_copy268_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid269_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid269_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w47_3_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid160_bh7_uid269_Out0_copy270_c0, Compressor_3_2_Freq500_uid160_bh7_uid269_Out0_copy270_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid271_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid271_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid271_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w24_11_c1 :  std_logic;
signal bh7_w25_13_c1 :  std_logic;
signal bh7_w26_12_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid271_Out0_copy272_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid273_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid273_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid273_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w27_14_c1 :  std_logic;
signal bh7_w28_12_c1 :  std_logic;
signal bh7_w29_14_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid273_Out0_copy274_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid275_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid275_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid275_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_15_c1 :  std_logic;
signal bh7_w30_12_c1 :  std_logic;
signal bh7_w31_14_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid275_Out0_copy276_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid277_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid277_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid277_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_15_c1 :  std_logic;
signal bh7_w32_12_c1 :  std_logic;
signal bh7_w33_14_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid277_Out0_copy278_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid279_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid279_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid279_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_15_c1 :  std_logic;
signal bh7_w34_12_c1 :  std_logic;
signal bh7_w35_14_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid279_Out0_copy280_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid281_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid281_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid281_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w35_15_c1 :  std_logic;
signal bh7_w36_12_c1 :  std_logic;
signal bh7_w37_14_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid281_Out0_copy282_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid283_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid283_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid283_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w37_15_c1 :  std_logic;
signal bh7_w38_12_c1 :  std_logic;
signal bh7_w39_14_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid283_Out0_copy284_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid285_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid285_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid285_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w39_15_c1 :  std_logic;
signal bh7_w40_12_c1 :  std_logic;
signal bh7_w41_12_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid285_Out0_copy286_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid287_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid287_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid287_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w41_13_c1 :  std_logic;
signal bh7_w42_11_c1 :  std_logic;
signal bh7_w43_12_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid287_Out0_copy288_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid289_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid289_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid289_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w43_13_c1 :  std_logic;
signal bh7_w44_7_c1 :  std_logic;
signal bh7_w45_8_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid289_Out0_copy290_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid291_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid291_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid291_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w45_9_c1 :  std_logic;
signal bh7_w46_5_c1 :  std_logic;
signal bh7_w47_4_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid291_Out0_copy292_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid293_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid293_In1_c0, Compressor_14_3_Freq500_uid164_bh7_uid293_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid293_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w47_5_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid293_Out0_copy294_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid295_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid295_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid295_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w17_2_c1 :  std_logic;
signal bh7_w18_3_c1 :  std_logic;
signal bh7_w19_4_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid295_Out0_copy296_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid297_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid297_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid297_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w19_5_c1 :  std_logic;
signal bh7_w20_7_c1 :  std_logic;
signal bh7_w21_8_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid297_Out0_copy298_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid299_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid299_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid299_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_9_c1 :  std_logic;
signal bh7_w22_10_c1 :  std_logic;
signal bh7_w23_13_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid299_Out0_copy300_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid301_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid301_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid301_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w23_14_c1 :  std_logic;
signal bh7_w24_12_c1 :  std_logic;
signal bh7_w25_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid301_Out0_copy302_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid303_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid303_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w25_15_c1 :  std_logic;
signal bh7_w26_13_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid160_bh7_uid303_Out0_copy304_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid305_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid305_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid305_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w26_14_c1 :  std_logic;
signal bh7_w27_15_c1 :  std_logic;
signal bh7_w28_13_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid305_Out0_copy306_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid307_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid160_bh7_uid307_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w28_14_c1 :  std_logic;
signal bh7_w29_16_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid160_bh7_uid307_Out0_copy308_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid309_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid309_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid309_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_17_c1 :  std_logic;
signal bh7_w30_13_c1 :  std_logic;
signal bh7_w31_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid309_Out0_copy310_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid311_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid311_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid311_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_17_c1 :  std_logic;
signal bh7_w32_13_c1 :  std_logic;
signal bh7_w33_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid311_Out0_copy312_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid313_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid313_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid313_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_17_c1 :  std_logic;
signal bh7_w34_13_c1 :  std_logic;
signal bh7_w35_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid313_Out0_copy314_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid315_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid315_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid315_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w35_17_c1 :  std_logic;
signal bh7_w36_13_c1 :  std_logic;
signal bh7_w37_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid315_Out0_copy316_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid317_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid317_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid317_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w37_17_c1 :  std_logic;
signal bh7_w38_13_c1 :  std_logic;
signal bh7_w39_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid317_Out0_copy318_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid319_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid319_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid156_bh7_uid319_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w39_17_c1 :  std_logic;
signal bh7_w40_13_c1 :  std_logic;
signal bh7_w41_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid156_bh7_uid319_Out0_copy320_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid321_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid321_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid321_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w41_15_c1 :  std_logic;
signal bh7_w42_12_c1 :  std_logic;
signal bh7_w43_14_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid321_Out0_copy322_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid323_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid323_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid323_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w43_15_c1 :  std_logic;
signal bh7_w44_8_c1 :  std_logic;
signal bh7_w45_10_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid323_Out0_copy324_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid325_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid325_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid325_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w45_11_c1 :  std_logic;
signal bh7_w46_6_c1 :  std_logic;
signal bh7_w47_6_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid325_Out0_copy326_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid327_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid327_In1_c0, Compressor_14_3_Freq500_uid164_bh7_uid327_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid164_bh7_uid327_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w47_7_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid164_bh7_uid327_Out0_copy328_c1 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh7_18_c1, tmp_bitheapResult_bh7_18_c2 :  std_logic_vector(18 downto 0);
signal bitheapFinalAdd_bh7_In0_c1 :  std_logic_vector(29 downto 0);
signal bitheapFinalAdd_bh7_In1_c1 :  std_logic_vector(29 downto 0);
signal bitheapFinalAdd_bh7_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh7_Out_c2 :  std_logic_vector(29 downto 0);
signal bitheapResult_bh7_c2 :  std_logic_vector(47 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               bh7_w17_1_c1 <= bh7_w17_1_c0;
               bh7_w18_2_c1 <= bh7_w18_2_c0;
               bh7_w19_3_c1 <= bh7_w19_3_c0;
               bh7_w20_6_c1 <= bh7_w20_6_c0;
               bh7_w21_7_c1 <= bh7_w21_7_c0;
               bh7_w24_9_c1 <= bh7_w24_9_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_copy246_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_copy246_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_copy248_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_copy248_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_copy250_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_copy250_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_copy252_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_copy252_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_copy254_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_copy254_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_copy256_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_copy256_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_copy258_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_copy258_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_copy260_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_copy260_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_copy262_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_copy262_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_copy264_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_copy264_c0;
               Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_copy266_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_copy266_c0;
               Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_copy268_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_copy268_c0;
               Compressor_3_2_Freq500_uid160_bh7_uid269_Out0_copy270_c1 <= Compressor_3_2_Freq500_uid160_bh7_uid269_Out0_copy270_c0;
               Compressor_14_3_Freq500_uid164_bh7_uid293_In1_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid293_In1_c0;
               Compressor_14_3_Freq500_uid164_bh7_uid327_In1_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid327_In1_c0;
            end if;
            if ce_2 = '1' then
               tmp_bitheapResult_bh7_18_c2 <= tmp_bitheapResult_bh7_18_c1;
            end if;
         end if;
      end process;
   XX_m6_c0 <= X ;
   YY_m6_c0 <= Y ;
   tile_0_X_c0 <= X(16 downto 0);
   tile_0_Y_c0 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq500_uid9
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 X => tile_0_X_c0,
                 Y => tile_0_Y_c0,
                 R => tile_0_output_c1);

   tile_0_filtered_output_c1 <= unsigned(tile_0_output_c1(40 downto 0));
   bh7_w0_0_c1 <= tile_0_filtered_output_c1(0);
   bh7_w1_0_c1 <= tile_0_filtered_output_c1(1);
   bh7_w2_0_c1 <= tile_0_filtered_output_c1(2);
   bh7_w3_0_c1 <= tile_0_filtered_output_c1(3);
   bh7_w4_0_c1 <= tile_0_filtered_output_c1(4);
   bh7_w5_0_c1 <= tile_0_filtered_output_c1(5);
   bh7_w6_0_c1 <= tile_0_filtered_output_c1(6);
   bh7_w7_0_c1 <= tile_0_filtered_output_c1(7);
   bh7_w8_0_c1 <= tile_0_filtered_output_c1(8);
   bh7_w9_0_c1 <= tile_0_filtered_output_c1(9);
   bh7_w10_0_c1 <= tile_0_filtered_output_c1(10);
   bh7_w11_0_c1 <= tile_0_filtered_output_c1(11);
   bh7_w12_0_c1 <= tile_0_filtered_output_c1(12);
   bh7_w13_0_c1 <= tile_0_filtered_output_c1(13);
   bh7_w14_0_c1 <= tile_0_filtered_output_c1(14);
   bh7_w15_0_c1 <= tile_0_filtered_output_c1(15);
   bh7_w16_0_c1 <= tile_0_filtered_output_c1(16);
   bh7_w17_0_c1 <= tile_0_filtered_output_c1(17);
   bh7_w18_0_c1 <= tile_0_filtered_output_c1(18);
   bh7_w19_0_c1 <= tile_0_filtered_output_c1(19);
   bh7_w20_0_c1 <= tile_0_filtered_output_c1(20);
   bh7_w21_0_c1 <= tile_0_filtered_output_c1(21);
   bh7_w22_0_c1 <= tile_0_filtered_output_c1(22);
   bh7_w23_0_c1 <= tile_0_filtered_output_c1(23);
   bh7_w24_0_c1 <= tile_0_filtered_output_c1(24);
   bh7_w25_0_c1 <= tile_0_filtered_output_c1(25);
   bh7_w26_0_c1 <= tile_0_filtered_output_c1(26);
   bh7_w27_0_c1 <= tile_0_filtered_output_c1(27);
   bh7_w28_0_c1 <= tile_0_filtered_output_c1(28);
   bh7_w29_0_c1 <= tile_0_filtered_output_c1(29);
   bh7_w30_0_c1 <= tile_0_filtered_output_c1(30);
   bh7_w31_0_c1 <= tile_0_filtered_output_c1(31);
   bh7_w32_0_c1 <= tile_0_filtered_output_c1(32);
   bh7_w33_0_c1 <= tile_0_filtered_output_c1(33);
   bh7_w34_0_c1 <= tile_0_filtered_output_c1(34);
   bh7_w35_0_c1 <= tile_0_filtered_output_c1(35);
   bh7_w36_0_c1 <= tile_0_filtered_output_c1(36);
   bh7_w37_0_c1 <= tile_0_filtered_output_c1(37);
   bh7_w38_0_c1 <= tile_0_filtered_output_c1(38);
   bh7_w39_0_c1 <= tile_0_filtered_output_c1(39);
   bh7_w40_0_c1 <= tile_0_filtered_output_c1(40);
   tile_1_X_c0 <= X(23 downto 23);
   tile_1_Y_c0 <= Y(23 downto 22);
   tile_1_mult: IntMultiplierLUT_1x2_Freq500_uid11
      port map ( clk  => clk,
                 X => tile_1_X_c0,
                 Y => tile_1_Y_c0,
                 R => tile_1_output_c0);

   tile_1_filtered_output_c0 <= unsigned(tile_1_output_c0(1 downto 0));
   bh7_w45_0_c0 <= tile_1_filtered_output_c0(0);
   bh7_w46_0_c0 <= tile_1_filtered_output_c0(1);
   tile_2_X_c0 <= X(22 downto 20);
   tile_2_Y_c0 <= Y(23 downto 22);
   tile_2_mult: IntMultiplierLUT_3x2_Freq500_uid13
      port map ( clk  => clk,
                 X => tile_2_X_c0,
                 Y => tile_2_Y_c0,
                 R => tile_2_output_c0);

   tile_2_filtered_output_c0 <= unsigned(tile_2_output_c0(4 downto 0));
   bh7_w42_0_c0 <= tile_2_filtered_output_c0(0);
   bh7_w43_0_c0 <= tile_2_filtered_output_c0(1);
   bh7_w44_0_c0 <= tile_2_filtered_output_c0(2);
   bh7_w45_1_c0 <= tile_2_filtered_output_c0(3);
   bh7_w46_1_c0 <= tile_2_filtered_output_c0(4);
   tile_3_X_c0 <= X(19 downto 17);
   tile_3_Y_c0 <= Y(23 downto 22);
   tile_3_mult: IntMultiplierLUT_3x2_Freq500_uid18
      port map ( clk  => clk,
                 X => tile_3_X_c0,
                 Y => tile_3_Y_c0,
                 R => tile_3_output_c0);

   tile_3_filtered_output_c0 <= unsigned(tile_3_output_c0(4 downto 0));
   bh7_w39_1_c0 <= tile_3_filtered_output_c0(0);
   bh7_w40_1_c0 <= tile_3_filtered_output_c0(1);
   bh7_w41_0_c0 <= tile_3_filtered_output_c0(2);
   bh7_w42_1_c0 <= tile_3_filtered_output_c0(3);
   bh7_w43_1_c0 <= tile_3_filtered_output_c0(4);
   tile_4_X_c0 <= X(23 downto 23);
   tile_4_Y_c0 <= Y(21 downto 20);
   tile_4_mult: IntMultiplierLUT_1x2_Freq500_uid23
      port map ( clk  => clk,
                 X => tile_4_X_c0,
                 Y => tile_4_Y_c0,
                 R => tile_4_output_c0);

   tile_4_filtered_output_c0 <= unsigned(tile_4_output_c0(1 downto 0));
   bh7_w43_2_c0 <= tile_4_filtered_output_c0(0);
   bh7_w44_1_c0 <= tile_4_filtered_output_c0(1);
   tile_5_X_c0 <= X(22 downto 20);
   tile_5_Y_c0 <= Y(21 downto 20);
   tile_5_mult: IntMultiplierLUT_3x2_Freq500_uid25
      port map ( clk  => clk,
                 X => tile_5_X_c0,
                 Y => tile_5_Y_c0,
                 R => tile_5_output_c0);

   tile_5_filtered_output_c0 <= unsigned(tile_5_output_c0(4 downto 0));
   bh7_w40_2_c0 <= tile_5_filtered_output_c0(0);
   bh7_w41_1_c0 <= tile_5_filtered_output_c0(1);
   bh7_w42_2_c0 <= tile_5_filtered_output_c0(2);
   bh7_w43_3_c0 <= tile_5_filtered_output_c0(3);
   bh7_w44_2_c0 <= tile_5_filtered_output_c0(4);
   tile_6_X_c0 <= X(19 downto 17);
   tile_6_Y_c0 <= Y(21 downto 20);
   tile_6_mult: IntMultiplierLUT_3x2_Freq500_uid30
      port map ( clk  => clk,
                 X => tile_6_X_c0,
                 Y => tile_6_Y_c0,
                 R => tile_6_output_c0);

   tile_6_filtered_output_c0 <= unsigned(tile_6_output_c0(4 downto 0));
   bh7_w37_1_c0 <= tile_6_filtered_output_c0(0);
   bh7_w38_1_c0 <= tile_6_filtered_output_c0(1);
   bh7_w39_2_c0 <= tile_6_filtered_output_c0(2);
   bh7_w40_3_c0 <= tile_6_filtered_output_c0(3);
   bh7_w41_2_c0 <= tile_6_filtered_output_c0(4);
   tile_7_X_c0 <= X(23 downto 23);
   tile_7_Y_c0 <= Y(19 downto 18);
   tile_7_mult: IntMultiplierLUT_1x2_Freq500_uid35
      port map ( clk  => clk,
                 X => tile_7_X_c0,
                 Y => tile_7_Y_c0,
                 R => tile_7_output_c0);

   tile_7_filtered_output_c0 <= unsigned(tile_7_output_c0(1 downto 0));
   bh7_w41_3_c0 <= tile_7_filtered_output_c0(0);
   bh7_w42_3_c0 <= tile_7_filtered_output_c0(1);
   tile_8_X_c0 <= X(22 downto 20);
   tile_8_Y_c0 <= Y(19 downto 18);
   tile_8_mult: IntMultiplierLUT_3x2_Freq500_uid37
      port map ( clk  => clk,
                 X => tile_8_X_c0,
                 Y => tile_8_Y_c0,
                 R => tile_8_output_c0);

   tile_8_filtered_output_c0 <= unsigned(tile_8_output_c0(4 downto 0));
   bh7_w38_2_c0 <= tile_8_filtered_output_c0(0);
   bh7_w39_3_c0 <= tile_8_filtered_output_c0(1);
   bh7_w40_4_c0 <= tile_8_filtered_output_c0(2);
   bh7_w41_4_c0 <= tile_8_filtered_output_c0(3);
   bh7_w42_4_c0 <= tile_8_filtered_output_c0(4);
   tile_9_X_c0 <= X(19 downto 17);
   tile_9_Y_c0 <= Y(19 downto 18);
   tile_9_mult: IntMultiplierLUT_3x2_Freq500_uid42
      port map ( clk  => clk,
                 X => tile_9_X_c0,
                 Y => tile_9_Y_c0,
                 R => tile_9_output_c0);

   tile_9_filtered_output_c0 <= unsigned(tile_9_output_c0(4 downto 0));
   bh7_w35_1_c0 <= tile_9_filtered_output_c0(0);
   bh7_w36_1_c0 <= tile_9_filtered_output_c0(1);
   bh7_w37_2_c0 <= tile_9_filtered_output_c0(2);
   bh7_w38_3_c0 <= tile_9_filtered_output_c0(3);
   bh7_w39_4_c0 <= tile_9_filtered_output_c0(4);
   tile_10_X_c0 <= X(23 downto 23);
   tile_10_Y_c0 <= Y(17 downto 16);
   tile_10_mult: IntMultiplierLUT_1x2_Freq500_uid47
      port map ( clk  => clk,
                 X => tile_10_X_c0,
                 Y => tile_10_Y_c0,
                 R => tile_10_output_c0);

   tile_10_filtered_output_c0 <= unsigned(tile_10_output_c0(1 downto 0));
   bh7_w39_5_c0 <= tile_10_filtered_output_c0(0);
   bh7_w40_5_c0 <= tile_10_filtered_output_c0(1);
   tile_11_X_c0 <= X(22 downto 20);
   tile_11_Y_c0 <= Y(17 downto 16);
   tile_11_mult: IntMultiplierLUT_3x2_Freq500_uid49
      port map ( clk  => clk,
                 X => tile_11_X_c0,
                 Y => tile_11_Y_c0,
                 R => tile_11_output_c0);

   tile_11_filtered_output_c0 <= unsigned(tile_11_output_c0(4 downto 0));
   bh7_w36_2_c0 <= tile_11_filtered_output_c0(0);
   bh7_w37_3_c0 <= tile_11_filtered_output_c0(1);
   bh7_w38_4_c0 <= tile_11_filtered_output_c0(2);
   bh7_w39_6_c0 <= tile_11_filtered_output_c0(3);
   bh7_w40_6_c0 <= tile_11_filtered_output_c0(4);
   tile_12_X_c0 <= X(19 downto 17);
   tile_12_Y_c0 <= Y(17 downto 16);
   tile_12_mult: IntMultiplierLUT_3x2_Freq500_uid54
      port map ( clk  => clk,
                 X => tile_12_X_c0,
                 Y => tile_12_Y_c0,
                 R => tile_12_output_c0);

   tile_12_filtered_output_c0 <= unsigned(tile_12_output_c0(4 downto 0));
   bh7_w33_1_c0 <= tile_12_filtered_output_c0(0);
   bh7_w34_1_c0 <= tile_12_filtered_output_c0(1);
   bh7_w35_2_c0 <= tile_12_filtered_output_c0(2);
   bh7_w36_3_c0 <= tile_12_filtered_output_c0(3);
   bh7_w37_4_c0 <= tile_12_filtered_output_c0(4);
   tile_13_X_c0 <= X(23 downto 23);
   tile_13_Y_c0 <= Y(15 downto 14);
   tile_13_mult: IntMultiplierLUT_1x2_Freq500_uid59
      port map ( clk  => clk,
                 X => tile_13_X_c0,
                 Y => tile_13_Y_c0,
                 R => tile_13_output_c0);

   tile_13_filtered_output_c0 <= unsigned(tile_13_output_c0(1 downto 0));
   bh7_w37_5_c0 <= tile_13_filtered_output_c0(0);
   bh7_w38_5_c0 <= tile_13_filtered_output_c0(1);
   tile_14_X_c0 <= X(22 downto 20);
   tile_14_Y_c0 <= Y(15 downto 14);
   tile_14_mult: IntMultiplierLUT_3x2_Freq500_uid61
      port map ( clk  => clk,
                 X => tile_14_X_c0,
                 Y => tile_14_Y_c0,
                 R => tile_14_output_c0);

   tile_14_filtered_output_c0 <= unsigned(tile_14_output_c0(4 downto 0));
   bh7_w34_2_c0 <= tile_14_filtered_output_c0(0);
   bh7_w35_3_c0 <= tile_14_filtered_output_c0(1);
   bh7_w36_4_c0 <= tile_14_filtered_output_c0(2);
   bh7_w37_6_c0 <= tile_14_filtered_output_c0(3);
   bh7_w38_6_c0 <= tile_14_filtered_output_c0(4);
   tile_15_X_c0 <= X(19 downto 17);
   tile_15_Y_c0 <= Y(15 downto 14);
   tile_15_mult: IntMultiplierLUT_3x2_Freq500_uid66
      port map ( clk  => clk,
                 X => tile_15_X_c0,
                 Y => tile_15_Y_c0,
                 R => tile_15_output_c0);

   tile_15_filtered_output_c0 <= unsigned(tile_15_output_c0(4 downto 0));
   bh7_w31_1_c0 <= tile_15_filtered_output_c0(0);
   bh7_w32_1_c0 <= tile_15_filtered_output_c0(1);
   bh7_w33_2_c0 <= tile_15_filtered_output_c0(2);
   bh7_w34_3_c0 <= tile_15_filtered_output_c0(3);
   bh7_w35_4_c0 <= tile_15_filtered_output_c0(4);
   tile_16_X_c0 <= X(23 downto 23);
   tile_16_Y_c0 <= Y(13 downto 12);
   tile_16_mult: IntMultiplierLUT_1x2_Freq500_uid71
      port map ( clk  => clk,
                 X => tile_16_X_c0,
                 Y => tile_16_Y_c0,
                 R => tile_16_output_c0);

   tile_16_filtered_output_c0 <= unsigned(tile_16_output_c0(1 downto 0));
   bh7_w35_5_c0 <= tile_16_filtered_output_c0(0);
   bh7_w36_5_c0 <= tile_16_filtered_output_c0(1);
   tile_17_X_c0 <= X(22 downto 20);
   tile_17_Y_c0 <= Y(13 downto 12);
   tile_17_mult: IntMultiplierLUT_3x2_Freq500_uid73
      port map ( clk  => clk,
                 X => tile_17_X_c0,
                 Y => tile_17_Y_c0,
                 R => tile_17_output_c0);

   tile_17_filtered_output_c0 <= unsigned(tile_17_output_c0(4 downto 0));
   bh7_w32_2_c0 <= tile_17_filtered_output_c0(0);
   bh7_w33_3_c0 <= tile_17_filtered_output_c0(1);
   bh7_w34_4_c0 <= tile_17_filtered_output_c0(2);
   bh7_w35_6_c0 <= tile_17_filtered_output_c0(3);
   bh7_w36_6_c0 <= tile_17_filtered_output_c0(4);
   tile_18_X_c0 <= X(19 downto 17);
   tile_18_Y_c0 <= Y(13 downto 12);
   tile_18_mult: IntMultiplierLUT_3x2_Freq500_uid78
      port map ( clk  => clk,
                 X => tile_18_X_c0,
                 Y => tile_18_Y_c0,
                 R => tile_18_output_c0);

   tile_18_filtered_output_c0 <= unsigned(tile_18_output_c0(4 downto 0));
   bh7_w29_1_c0 <= tile_18_filtered_output_c0(0);
   bh7_w30_1_c0 <= tile_18_filtered_output_c0(1);
   bh7_w31_2_c0 <= tile_18_filtered_output_c0(2);
   bh7_w32_3_c0 <= tile_18_filtered_output_c0(3);
   bh7_w33_4_c0 <= tile_18_filtered_output_c0(4);
   tile_19_X_c0 <= X(23 downto 23);
   tile_19_Y_c0 <= Y(11 downto 10);
   tile_19_mult: IntMultiplierLUT_1x2_Freq500_uid83
      port map ( clk  => clk,
                 X => tile_19_X_c0,
                 Y => tile_19_Y_c0,
                 R => tile_19_output_c0);

   tile_19_filtered_output_c0 <= unsigned(tile_19_output_c0(1 downto 0));
   bh7_w33_5_c0 <= tile_19_filtered_output_c0(0);
   bh7_w34_5_c0 <= tile_19_filtered_output_c0(1);
   tile_20_X_c0 <= X(22 downto 20);
   tile_20_Y_c0 <= Y(11 downto 10);
   tile_20_mult: IntMultiplierLUT_3x2_Freq500_uid85
      port map ( clk  => clk,
                 X => tile_20_X_c0,
                 Y => tile_20_Y_c0,
                 R => tile_20_output_c0);

   tile_20_filtered_output_c0 <= unsigned(tile_20_output_c0(4 downto 0));
   bh7_w30_2_c0 <= tile_20_filtered_output_c0(0);
   bh7_w31_3_c0 <= tile_20_filtered_output_c0(1);
   bh7_w32_4_c0 <= tile_20_filtered_output_c0(2);
   bh7_w33_6_c0 <= tile_20_filtered_output_c0(3);
   bh7_w34_6_c0 <= tile_20_filtered_output_c0(4);
   tile_21_X_c0 <= X(19 downto 17);
   tile_21_Y_c0 <= Y(11 downto 10);
   tile_21_mult: IntMultiplierLUT_3x2_Freq500_uid90
      port map ( clk  => clk,
                 X => tile_21_X_c0,
                 Y => tile_21_Y_c0,
                 R => tile_21_output_c0);

   tile_21_filtered_output_c0 <= unsigned(tile_21_output_c0(4 downto 0));
   bh7_w27_1_c0 <= tile_21_filtered_output_c0(0);
   bh7_w28_1_c0 <= tile_21_filtered_output_c0(1);
   bh7_w29_2_c0 <= tile_21_filtered_output_c0(2);
   bh7_w30_3_c0 <= tile_21_filtered_output_c0(3);
   bh7_w31_4_c0 <= tile_21_filtered_output_c0(4);
   tile_22_X_c0 <= X(23 downto 23);
   tile_22_Y_c0 <= Y(9 downto 8);
   tile_22_mult: IntMultiplierLUT_1x2_Freq500_uid95
      port map ( clk  => clk,
                 X => tile_22_X_c0,
                 Y => tile_22_Y_c0,
                 R => tile_22_output_c0);

   tile_22_filtered_output_c0 <= unsigned(tile_22_output_c0(1 downto 0));
   bh7_w31_5_c0 <= tile_22_filtered_output_c0(0);
   bh7_w32_5_c0 <= tile_22_filtered_output_c0(1);
   tile_23_X_c0 <= X(22 downto 20);
   tile_23_Y_c0 <= Y(9 downto 8);
   tile_23_mult: IntMultiplierLUT_3x2_Freq500_uid97
      port map ( clk  => clk,
                 X => tile_23_X_c0,
                 Y => tile_23_Y_c0,
                 R => tile_23_output_c0);

   tile_23_filtered_output_c0 <= unsigned(tile_23_output_c0(4 downto 0));
   bh7_w28_2_c0 <= tile_23_filtered_output_c0(0);
   bh7_w29_3_c0 <= tile_23_filtered_output_c0(1);
   bh7_w30_4_c0 <= tile_23_filtered_output_c0(2);
   bh7_w31_6_c0 <= tile_23_filtered_output_c0(3);
   bh7_w32_6_c0 <= tile_23_filtered_output_c0(4);
   tile_24_X_c0 <= X(19 downto 17);
   tile_24_Y_c0 <= Y(9 downto 8);
   tile_24_mult: IntMultiplierLUT_3x2_Freq500_uid102
      port map ( clk  => clk,
                 X => tile_24_X_c0,
                 Y => tile_24_Y_c0,
                 R => tile_24_output_c0);

   tile_24_filtered_output_c0 <= unsigned(tile_24_output_c0(4 downto 0));
   bh7_w25_1_c0 <= tile_24_filtered_output_c0(0);
   bh7_w26_1_c0 <= tile_24_filtered_output_c0(1);
   bh7_w27_2_c0 <= tile_24_filtered_output_c0(2);
   bh7_w28_3_c0 <= tile_24_filtered_output_c0(3);
   bh7_w29_4_c0 <= tile_24_filtered_output_c0(4);
   tile_25_X_c0 <= X(23 downto 23);
   tile_25_Y_c0 <= Y(7 downto 6);
   tile_25_mult: IntMultiplierLUT_1x2_Freq500_uid107
      port map ( clk  => clk,
                 X => tile_25_X_c0,
                 Y => tile_25_Y_c0,
                 R => tile_25_output_c0);

   tile_25_filtered_output_c0 <= unsigned(tile_25_output_c0(1 downto 0));
   bh7_w29_5_c0 <= tile_25_filtered_output_c0(0);
   bh7_w30_5_c0 <= tile_25_filtered_output_c0(1);
   tile_26_X_c0 <= X(22 downto 20);
   tile_26_Y_c0 <= Y(7 downto 6);
   tile_26_mult: IntMultiplierLUT_3x2_Freq500_uid109
      port map ( clk  => clk,
                 X => tile_26_X_c0,
                 Y => tile_26_Y_c0,
                 R => tile_26_output_c0);

   tile_26_filtered_output_c0 <= unsigned(tile_26_output_c0(4 downto 0));
   bh7_w26_2_c0 <= tile_26_filtered_output_c0(0);
   bh7_w27_3_c0 <= tile_26_filtered_output_c0(1);
   bh7_w28_4_c0 <= tile_26_filtered_output_c0(2);
   bh7_w29_6_c0 <= tile_26_filtered_output_c0(3);
   bh7_w30_6_c0 <= tile_26_filtered_output_c0(4);
   tile_27_X_c0 <= X(19 downto 17);
   tile_27_Y_c0 <= Y(7 downto 6);
   tile_27_mult: IntMultiplierLUT_3x2_Freq500_uid114
      port map ( clk  => clk,
                 X => tile_27_X_c0,
                 Y => tile_27_Y_c0,
                 R => tile_27_output_c0);

   tile_27_filtered_output_c0 <= unsigned(tile_27_output_c0(4 downto 0));
   bh7_w23_1_c0 <= tile_27_filtered_output_c0(0);
   bh7_w24_1_c0 <= tile_27_filtered_output_c0(1);
   bh7_w25_2_c0 <= tile_27_filtered_output_c0(2);
   bh7_w26_3_c0 <= tile_27_filtered_output_c0(3);
   bh7_w27_4_c0 <= tile_27_filtered_output_c0(4);
   tile_28_X_c0 <= X(23 downto 23);
   tile_28_Y_c0 <= Y(5 downto 4);
   tile_28_mult: IntMultiplierLUT_1x2_Freq500_uid119
      port map ( clk  => clk,
                 X => tile_28_X_c0,
                 Y => tile_28_Y_c0,
                 R => tile_28_output_c0);

   tile_28_filtered_output_c0 <= unsigned(tile_28_output_c0(1 downto 0));
   bh7_w27_5_c0 <= tile_28_filtered_output_c0(0);
   bh7_w28_5_c0 <= tile_28_filtered_output_c0(1);
   tile_29_X_c0 <= X(22 downto 20);
   tile_29_Y_c0 <= Y(5 downto 4);
   tile_29_mult: IntMultiplierLUT_3x2_Freq500_uid121
      port map ( clk  => clk,
                 X => tile_29_X_c0,
                 Y => tile_29_Y_c0,
                 R => tile_29_output_c0);

   tile_29_filtered_output_c0 <= unsigned(tile_29_output_c0(4 downto 0));
   bh7_w24_2_c0 <= tile_29_filtered_output_c0(0);
   bh7_w25_3_c0 <= tile_29_filtered_output_c0(1);
   bh7_w26_4_c0 <= tile_29_filtered_output_c0(2);
   bh7_w27_6_c0 <= tile_29_filtered_output_c0(3);
   bh7_w28_6_c0 <= tile_29_filtered_output_c0(4);
   tile_30_X_c0 <= X(19 downto 17);
   tile_30_Y_c0 <= Y(5 downto 4);
   tile_30_mult: IntMultiplierLUT_3x2_Freq500_uid126
      port map ( clk  => clk,
                 X => tile_30_X_c0,
                 Y => tile_30_Y_c0,
                 R => tile_30_output_c0);

   tile_30_filtered_output_c0 <= unsigned(tile_30_output_c0(4 downto 0));
   bh7_w21_1_c0 <= tile_30_filtered_output_c0(0);
   bh7_w22_1_c0 <= tile_30_filtered_output_c0(1);
   bh7_w23_2_c0 <= tile_30_filtered_output_c0(2);
   bh7_w24_3_c0 <= tile_30_filtered_output_c0(3);
   bh7_w25_4_c0 <= tile_30_filtered_output_c0(4);
   tile_31_X_c0 <= X(23 downto 23);
   tile_31_Y_c0 <= Y(3 downto 2);
   tile_31_mult: IntMultiplierLUT_1x2_Freq500_uid131
      port map ( clk  => clk,
                 X => tile_31_X_c0,
                 Y => tile_31_Y_c0,
                 R => tile_31_output_c0);

   tile_31_filtered_output_c0 <= unsigned(tile_31_output_c0(1 downto 0));
   bh7_w25_5_c0 <= tile_31_filtered_output_c0(0);
   bh7_w26_5_c0 <= tile_31_filtered_output_c0(1);
   tile_32_X_c0 <= X(22 downto 20);
   tile_32_Y_c0 <= Y(3 downto 2);
   tile_32_mult: IntMultiplierLUT_3x2_Freq500_uid133
      port map ( clk  => clk,
                 X => tile_32_X_c0,
                 Y => tile_32_Y_c0,
                 R => tile_32_output_c0);

   tile_32_filtered_output_c0 <= unsigned(tile_32_output_c0(4 downto 0));
   bh7_w22_2_c0 <= tile_32_filtered_output_c0(0);
   bh7_w23_3_c0 <= tile_32_filtered_output_c0(1);
   bh7_w24_4_c0 <= tile_32_filtered_output_c0(2);
   bh7_w25_6_c0 <= tile_32_filtered_output_c0(3);
   bh7_w26_6_c0 <= tile_32_filtered_output_c0(4);
   tile_33_X_c0 <= X(19 downto 17);
   tile_33_Y_c0 <= Y(3 downto 2);
   tile_33_mult: IntMultiplierLUT_3x2_Freq500_uid138
      port map ( clk  => clk,
                 X => tile_33_X_c0,
                 Y => tile_33_Y_c0,
                 R => tile_33_output_c0);

   tile_33_filtered_output_c0 <= unsigned(tile_33_output_c0(4 downto 0));
   bh7_w19_1_c0 <= tile_33_filtered_output_c0(0);
   bh7_w20_1_c0 <= tile_33_filtered_output_c0(1);
   bh7_w21_2_c0 <= tile_33_filtered_output_c0(2);
   bh7_w22_3_c0 <= tile_33_filtered_output_c0(3);
   bh7_w23_4_c0 <= tile_33_filtered_output_c0(4);
   tile_34_X_c0 <= X(23 downto 23);
   tile_34_Y_c0 <= Y(1 downto 0);
   tile_34_mult: IntMultiplierLUT_1x2_Freq500_uid143
      port map ( clk  => clk,
                 X => tile_34_X_c0,
                 Y => tile_34_Y_c0,
                 R => tile_34_output_c0);

   tile_34_filtered_output_c0 <= unsigned(tile_34_output_c0(1 downto 0));
   bh7_w23_5_c0 <= tile_34_filtered_output_c0(0);
   bh7_w24_5_c0 <= tile_34_filtered_output_c0(1);
   tile_35_X_c0 <= X(22 downto 20);
   tile_35_Y_c0 <= Y(1 downto 0);
   tile_35_mult: IntMultiplierLUT_3x2_Freq500_uid145
      port map ( clk  => clk,
                 X => tile_35_X_c0,
                 Y => tile_35_Y_c0,
                 R => tile_35_output_c0);

   tile_35_filtered_output_c0 <= unsigned(tile_35_output_c0(4 downto 0));
   bh7_w20_2_c0 <= tile_35_filtered_output_c0(0);
   bh7_w21_3_c0 <= tile_35_filtered_output_c0(1);
   bh7_w22_4_c0 <= tile_35_filtered_output_c0(2);
   bh7_w23_6_c0 <= tile_35_filtered_output_c0(3);
   bh7_w24_6_c0 <= tile_35_filtered_output_c0(4);
   tile_36_X_c0 <= X(19 downto 17);
   tile_36_Y_c0 <= Y(1 downto 0);
   tile_36_mult: IntMultiplierLUT_3x2_Freq500_uid150
      port map ( clk  => clk,
                 X => tile_36_X_c0,
                 Y => tile_36_Y_c0,
                 R => tile_36_output_c0);

   tile_36_filtered_output_c0 <= unsigned(tile_36_output_c0(4 downto 0));
   bh7_w17_1_c0 <= tile_36_filtered_output_c0(0);
   bh7_w18_1_c0 <= tile_36_filtered_output_c0(1);
   bh7_w19_2_c0 <= tile_36_filtered_output_c0(2);
   bh7_w20_3_c0 <= tile_36_filtered_output_c0(3);
   bh7_w21_4_c0 <= tile_36_filtered_output_c0(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq500_uid156_bh7_uid157_In0_c0 <= "" & bh7_w18_1_c0 & "0" & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid157_In1_c0 <= "" & bh7_w19_1_c0 & bh7_w19_2_c0;
   bh7_w18_2_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid157_Out0_c0(0);
   bh7_w19_3_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid157_Out0_c0(1);
   bh7_w20_4_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid157_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid157: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid157_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid157_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid157_Out0_copy158_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid157_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid157_Out0_copy158_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid160_bh7_uid161_In0_c0 <= "" & bh7_w20_1_c0 & bh7_w20_2_c0 & bh7_w20_3_c0;
   bh7_w20_5_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid161_Out0_c0(0);
   bh7_w21_5_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid161_Out0_c0(1);
   Compressor_3_2_Freq500_uid160_uid161: Compressor_3_2_Freq500_uid160
      port map ( X0 => Compressor_3_2_Freq500_uid160_bh7_uid161_In0_c0,
                 R => Compressor_3_2_Freq500_uid160_bh7_uid161_Out0_copy162_c0);
   Compressor_3_2_Freq500_uid160_bh7_uid161_Out0_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid161_Out0_copy162_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid165_In0_c0 <= "" & bh7_w21_1_c0 & bh7_w21_2_c0 & bh7_w21_3_c0 & bh7_w21_4_c0;
   Compressor_14_3_Freq500_uid164_bh7_uid165_In1_c0 <= "" & bh7_w22_1_c0;
   bh7_w21_6_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid165_Out0_c0(0);
   bh7_w22_5_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid165_Out0_c0(1);
   bh7_w23_7_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid165_Out0_c0(2);
   Compressor_14_3_Freq500_uid164_uid165: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid165_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid165_In1_c0,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid165_Out0_copy166_c0);
   Compressor_14_3_Freq500_uid164_bh7_uid165_Out0_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid165_Out0_copy166_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid160_bh7_uid167_In0_c0 <= "" & bh7_w22_2_c0 & bh7_w22_3_c0 & bh7_w22_4_c0;
   bh7_w22_6_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid167_Out0_c0(0);
   bh7_w23_8_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid167_Out0_c0(1);
   Compressor_3_2_Freq500_uid160_uid167: Compressor_3_2_Freq500_uid160
      port map ( X0 => Compressor_3_2_Freq500_uid160_bh7_uid167_In0_c0,
                 R => Compressor_3_2_Freq500_uid160_bh7_uid167_Out0_copy168_c0);
   Compressor_3_2_Freq500_uid160_bh7_uid167_Out0_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid167_Out0_copy168_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid171_In0_c0 <= "" & bh7_w23_1_c0 & bh7_w23_2_c0 & bh7_w23_3_c0 & bh7_w23_4_c0 & bh7_w23_5_c0 & bh7_w23_6_c0;
   bh7_w23_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid171_Out0_c0(0);
   bh7_w24_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid171_Out0_c0(1);
   bh7_w25_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid171_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid171: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid171_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid171_Out0_copy172_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid171_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid171_Out0_copy172_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid173_In0_c0 <= "" & bh7_w24_1_c0 & bh7_w24_2_c0 & bh7_w24_3_c0 & bh7_w24_4_c0 & bh7_w24_5_c0 & bh7_w24_6_c0;
   bh7_w24_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid173_Out0_c0(0);
   bh7_w25_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid173_Out0_c0(1);
   bh7_w26_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid173_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid173: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid173_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid173_Out0_copy174_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid173_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid173_Out0_copy174_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid175_In0_c0 <= "" & bh7_w25_1_c0 & bh7_w25_2_c0 & bh7_w25_3_c0 & bh7_w25_4_c0 & bh7_w25_5_c0 & bh7_w25_6_c0;
   bh7_w25_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid175_Out0_c0(0);
   bh7_w26_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid175_Out0_c0(1);
   bh7_w27_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid175_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid175: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid175_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid175_Out0_copy176_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid175_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid175_Out0_copy176_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid177_In0_c0 <= "" & bh7_w26_1_c0 & bh7_w26_2_c0 & bh7_w26_3_c0 & bh7_w26_4_c0 & bh7_w26_5_c0 & bh7_w26_6_c0;
   bh7_w26_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid177_Out0_c0(0);
   bh7_w27_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid177_Out0_c0(1);
   bh7_w28_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid177_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid177: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid177_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid177_Out0_copy178_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid177_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid177_Out0_copy178_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid179_In0_c0 <= "" & bh7_w27_1_c0 & bh7_w27_2_c0 & bh7_w27_3_c0 & bh7_w27_4_c0 & bh7_w27_5_c0 & bh7_w27_6_c0;
   bh7_w27_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid179_Out0_c0(0);
   bh7_w28_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid179_Out0_c0(1);
   bh7_w29_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid179_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid179: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid179_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid179_Out0_copy180_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid179_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid179_Out0_copy180_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid181_In0_c0 <= "" & bh7_w28_1_c0 & bh7_w28_2_c0 & bh7_w28_3_c0 & bh7_w28_4_c0 & bh7_w28_5_c0 & bh7_w28_6_c0;
   bh7_w28_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid181_Out0_c0(0);
   bh7_w29_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid181_Out0_c0(1);
   bh7_w30_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid181_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid181: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid181_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid181_Out0_copy182_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid181_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid181_Out0_copy182_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid183_In0_c0 <= "" & bh7_w29_1_c0 & bh7_w29_2_c0 & bh7_w29_3_c0 & bh7_w29_4_c0 & bh7_w29_5_c0 & bh7_w29_6_c0;
   bh7_w29_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid183_Out0_c0(0);
   bh7_w30_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid183_Out0_c0(1);
   bh7_w31_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid183_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid183: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid183_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid183_Out0_copy184_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid183_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid183_Out0_copy184_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid185_In0_c0 <= "" & bh7_w30_1_c0 & bh7_w30_2_c0 & bh7_w30_3_c0 & bh7_w30_4_c0 & bh7_w30_5_c0 & bh7_w30_6_c0;
   bh7_w30_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid185_Out0_c0(0);
   bh7_w31_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid185_Out0_c0(1);
   bh7_w32_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid185_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid185: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid185_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid185_Out0_copy186_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid185_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid185_Out0_copy186_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid187_In0_c0 <= "" & bh7_w31_1_c0 & bh7_w31_2_c0 & bh7_w31_3_c0 & bh7_w31_4_c0 & bh7_w31_5_c0 & bh7_w31_6_c0;
   bh7_w31_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid187_Out0_c0(0);
   bh7_w32_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid187_Out0_c0(1);
   bh7_w33_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid187_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid187: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid187_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid187_Out0_copy188_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid187_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid187_Out0_copy188_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid189_In0_c0 <= "" & bh7_w32_1_c0 & bh7_w32_2_c0 & bh7_w32_3_c0 & bh7_w32_4_c0 & bh7_w32_5_c0 & bh7_w32_6_c0;
   bh7_w32_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid189_Out0_c0(0);
   bh7_w33_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid189_Out0_c0(1);
   bh7_w34_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid189_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid189: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid189_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid189_Out0_copy190_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid189_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid189_Out0_copy190_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid191_In0_c0 <= "" & bh7_w33_1_c0 & bh7_w33_2_c0 & bh7_w33_3_c0 & bh7_w33_4_c0 & bh7_w33_5_c0 & bh7_w33_6_c0;
   bh7_w33_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid191_Out0_c0(0);
   bh7_w34_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid191_Out0_c0(1);
   bh7_w35_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid191_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid191: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid191_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid191_Out0_copy192_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid191_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid191_Out0_copy192_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid193_In0_c0 <= "" & bh7_w34_1_c0 & bh7_w34_2_c0 & bh7_w34_3_c0 & bh7_w34_4_c0 & bh7_w34_5_c0 & bh7_w34_6_c0;
   bh7_w34_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid193_Out0_c0(0);
   bh7_w35_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid193_Out0_c0(1);
   bh7_w36_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid193_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid193: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid193_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid193_Out0_copy194_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid193_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid193_Out0_copy194_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid195_In0_c0 <= "" & bh7_w35_1_c0 & bh7_w35_2_c0 & bh7_w35_3_c0 & bh7_w35_4_c0 & bh7_w35_5_c0 & bh7_w35_6_c0;
   bh7_w35_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid195_Out0_c0(0);
   bh7_w36_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid195_Out0_c0(1);
   bh7_w37_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid195_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid195: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid195_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid195_Out0_copy196_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid195_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid195_Out0_copy196_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid197_In0_c0 <= "" & bh7_w36_1_c0 & bh7_w36_2_c0 & bh7_w36_3_c0 & bh7_w36_4_c0 & bh7_w36_5_c0 & bh7_w36_6_c0;
   bh7_w36_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid197_Out0_c0(0);
   bh7_w37_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid197_Out0_c0(1);
   bh7_w38_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid197_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid197: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid197_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid197_Out0_copy198_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid197_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid197_Out0_copy198_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid199_In0_c0 <= "" & bh7_w37_1_c0 & bh7_w37_2_c0 & bh7_w37_3_c0 & bh7_w37_4_c0 & bh7_w37_5_c0 & bh7_w37_6_c0;
   bh7_w37_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid199_Out0_c0(0);
   bh7_w38_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid199_Out0_c0(1);
   bh7_w39_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid199_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid199: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid199_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid199_Out0_copy200_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid199_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid199_Out0_copy200_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid201_In0_c0 <= "" & bh7_w38_1_c0 & bh7_w38_2_c0 & bh7_w38_3_c0 & bh7_w38_4_c0 & bh7_w38_5_c0 & bh7_w38_6_c0;
   bh7_w38_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid201_Out0_c0(0);
   bh7_w39_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid201_Out0_c0(1);
   bh7_w40_7_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid201_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid201: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid201_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid201_Out0_copy202_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid201_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid201_Out0_copy202_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid203_In0_c0 <= "" & bh7_w39_1_c0 & bh7_w39_2_c0 & bh7_w39_3_c0 & bh7_w39_4_c0 & bh7_w39_5_c0 & bh7_w39_6_c0;
   bh7_w39_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid203_Out0_c0(0);
   bh7_w40_8_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid203_Out0_c0(1);
   bh7_w41_5_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid203_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid203: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid203_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid203_Out0_copy204_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid203_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid203_Out0_copy204_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid170_bh7_uid205_In0_c0 <= "" & bh7_w40_1_c0 & bh7_w40_2_c0 & bh7_w40_3_c0 & bh7_w40_4_c0 & bh7_w40_5_c0 & bh7_w40_6_c0;
   bh7_w40_9_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid205_Out0_c0(0);
   bh7_w41_6_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid205_Out0_c0(1);
   bh7_w42_5_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid205_Out0_c0(2);
   Compressor_6_3_Freq500_uid170_uid205: Compressor_6_3_Freq500_uid170
      port map ( X0 => Compressor_6_3_Freq500_uid170_bh7_uid205_In0_c0,
                 R => Compressor_6_3_Freq500_uid170_bh7_uid205_Out0_copy206_c0);
   Compressor_6_3_Freq500_uid170_bh7_uid205_Out0_c0 <= Compressor_6_3_Freq500_uid170_bh7_uid205_Out0_copy206_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid207_In0_c0 <= "" & bh7_w41_0_c0 & bh7_w41_1_c0 & bh7_w41_2_c0 & bh7_w41_3_c0;
   Compressor_14_3_Freq500_uid164_bh7_uid207_In1_c0 <= "" & bh7_w42_0_c0;
   bh7_w41_7_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid207_Out0_c0(0);
   bh7_w42_6_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid207_Out0_c0(1);
   bh7_w43_4_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid207_Out0_c0(2);
   Compressor_14_3_Freq500_uid164_uid207: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid207_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid207_In1_c0,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid207_Out0_copy208_c0);
   Compressor_14_3_Freq500_uid164_bh7_uid207_Out0_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid207_Out0_copy208_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid209_In0_c0 <= "" & bh7_w42_1_c0 & bh7_w42_2_c0 & bh7_w42_3_c0 & bh7_w42_4_c0;
   Compressor_14_3_Freq500_uid164_bh7_uid209_In1_c0 <= "" & bh7_w43_0_c0;
   bh7_w42_7_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid209_Out0_c0(0);
   bh7_w43_5_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid209_Out0_c0(1);
   bh7_w44_3_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid209_Out0_c0(2);
   Compressor_14_3_Freq500_uid164_uid209: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid209_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid209_In1_c0,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid209_Out0_copy210_c0);
   Compressor_14_3_Freq500_uid164_bh7_uid209_Out0_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid209_Out0_copy210_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid211_In0_c0 <= "" & bh7_w43_1_c0 & bh7_w43_2_c0 & bh7_w43_3_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid211_In1_c0 <= "" & bh7_w44_0_c0 & bh7_w44_1_c0;
   bh7_w43_6_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid211_Out0_c0(0);
   bh7_w44_4_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid211_Out0_c0(1);
   bh7_w45_2_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid211_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid211: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid211_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid211_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid211_Out0_copy212_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid211_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid211_Out0_copy212_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid213_In0_c0 <= "" & bh7_w45_0_c0 & bh7_w45_1_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid213_In1_c0 <= "" & bh7_w46_0_c0 & bh7_w46_1_c0;
   bh7_w45_3_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid213_Out0_c0(0);
   bh7_w46_2_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid213_Out0_c0(1);
   bh7_w47_0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid213_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid213: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid213_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid213_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid213_Out0_copy214_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid213_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid213_Out0_copy214_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid215_In0_c0 <= "" & bh7_w20_5_c0 & bh7_w20_4_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid215_In1_c0 <= "" & bh7_w21_6_c0 & bh7_w21_5_c0;
   bh7_w20_6_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid215_Out0_c0(0);
   bh7_w21_7_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid215_Out0_c0(1);
   bh7_w22_7_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid215_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid215: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid215_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid215_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid215_Out0_copy216_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid215_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid215_Out0_copy216_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid160_bh7_uid217_In0_c0 <= "" & bh7_w22_6_c0 & bh7_w22_5_c0 & "0";
   bh7_w22_8_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid217_Out0_c0(0);
   bh7_w23_10_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid217_Out0_c0(1);
   Compressor_3_2_Freq500_uid160_uid217: Compressor_3_2_Freq500_uid160
      port map ( X0 => Compressor_3_2_Freq500_uid160_bh7_uid217_In0_c0,
                 R => Compressor_3_2_Freq500_uid160_bh7_uid217_Out0_copy218_c0);
   Compressor_3_2_Freq500_uid160_bh7_uid217_Out0_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid217_Out0_copy218_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid219_In0_c0 <= "" & bh7_w23_8_c0 & bh7_w23_7_c0 & bh7_w23_9_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid219_In1_c0 <= "" & bh7_w24_8_c0 & bh7_w24_7_c0;
   bh7_w23_11_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid219_Out0_c0(0);
   bh7_w24_9_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid219_Out0_c0(1);
   bh7_w25_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid219_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid219: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid219_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid219_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid219_Out0_copy220_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid219_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid219_Out0_copy220_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid221_In0_c0 <= "" & bh7_w25_9_c0 & bh7_w25_8_c0 & bh7_w25_7_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid221_In1_c0 <= "" & bh7_w26_9_c0 & bh7_w26_8_c0;
   bh7_w25_11_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid221_Out0_c0(0);
   bh7_w26_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid221_Out0_c0(1);
   bh7_w27_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid221_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid221: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid221_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid221_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid221_Out0_copy222_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid221_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid221_Out0_copy222_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid223_In0_c0 <= "" & bh7_w27_9_c0 & bh7_w27_8_c0 & bh7_w27_7_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid223_In1_c0 <= "" & bh7_w28_9_c0 & bh7_w28_8_c0;
   bh7_w27_11_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid223_Out0_c0(0);
   bh7_w28_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid223_Out0_c0(1);
   bh7_w29_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid223_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid223: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid223_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid223_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid223_Out0_copy224_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid223_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid223_Out0_copy224_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid225_In0_c0 <= "" & bh7_w29_9_c0 & bh7_w29_8_c0 & bh7_w29_7_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid225_In1_c0 <= "" & bh7_w30_9_c0 & bh7_w30_8_c0;
   bh7_w29_11_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid225_Out0_c0(0);
   bh7_w30_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid225_Out0_c0(1);
   bh7_w31_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid225_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid225: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid225_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid225_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid225_Out0_copy226_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid225_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid225_Out0_copy226_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid227_In0_c0 <= "" & bh7_w31_9_c0 & bh7_w31_8_c0 & bh7_w31_7_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid227_In1_c0 <= "" & bh7_w32_9_c0 & bh7_w32_8_c0;
   bh7_w31_11_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid227_Out0_c0(0);
   bh7_w32_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid227_Out0_c0(1);
   bh7_w33_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid227_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid227: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid227_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid227_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid227_Out0_copy228_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid227_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid227_Out0_copy228_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid229_In0_c0 <= "" & bh7_w33_9_c0 & bh7_w33_8_c0 & bh7_w33_7_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid229_In1_c0 <= "" & bh7_w34_9_c0 & bh7_w34_8_c0;
   bh7_w33_11_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid229_Out0_c0(0);
   bh7_w34_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid229_Out0_c0(1);
   bh7_w35_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid229_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid229: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid229_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid229_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid229_Out0_copy230_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid229_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid229_Out0_copy230_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid231_In0_c0 <= "" & bh7_w35_9_c0 & bh7_w35_8_c0 & bh7_w35_7_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid231_In1_c0 <= "" & bh7_w36_9_c0 & bh7_w36_8_c0;
   bh7_w35_11_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid231_Out0_c0(0);
   bh7_w36_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid231_Out0_c0(1);
   bh7_w37_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid231_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid231: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid231_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid231_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid231_Out0_copy232_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid231_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid231_Out0_copy232_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid233_In0_c0 <= "" & bh7_w37_9_c0 & bh7_w37_8_c0 & bh7_w37_7_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid233_In1_c0 <= "" & bh7_w38_9_c0 & bh7_w38_8_c0;
   bh7_w37_11_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid233_Out0_c0(0);
   bh7_w38_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid233_Out0_c0(1);
   bh7_w39_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid233_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid233: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid233_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid233_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid233_Out0_copy234_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid233_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid233_Out0_copy234_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid235_In0_c0 <= "" & bh7_w39_9_c0 & bh7_w39_8_c0 & bh7_w39_7_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid235_In1_c0 <= "" & bh7_w40_9_c0 & bh7_w40_8_c0;
   bh7_w39_11_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid235_Out0_c0(0);
   bh7_w40_10_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid235_Out0_c0(1);
   bh7_w41_8_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid235_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid235: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid235_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid235_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid235_Out0_copy236_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid235_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid235_Out0_copy236_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid237_In0_c0 <= "" & bh7_w41_4_c0 & bh7_w41_7_c0 & bh7_w41_6_c0 & bh7_w41_5_c0;
   Compressor_14_3_Freq500_uid164_bh7_uid237_In1_c0 <= "" & "0";
   bh7_w41_9_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid237_Out0_c0(0);
   bh7_w42_8_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid237_Out0_c0(1);
   bh7_w43_7_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid237_Out0_c0(2);
   Compressor_14_3_Freq500_uid164_uid237: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid237_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid237_In1_c0,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid237_Out0_copy238_c0);
   Compressor_14_3_Freq500_uid164_bh7_uid237_Out0_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid237_Out0_copy238_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid160_bh7_uid239_In0_c0 <= "" & bh7_w42_7_c0 & bh7_w42_6_c0 & bh7_w42_5_c0;
   bh7_w42_9_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid239_Out0_c0(0);
   bh7_w43_8_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid239_Out0_c0(1);
   Compressor_3_2_Freq500_uid160_uid239: Compressor_3_2_Freq500_uid160
      port map ( X0 => Compressor_3_2_Freq500_uid160_bh7_uid239_In0_c0,
                 R => Compressor_3_2_Freq500_uid160_bh7_uid239_Out0_copy240_c0);
   Compressor_3_2_Freq500_uid160_bh7_uid239_Out0_c0 <= Compressor_3_2_Freq500_uid160_bh7_uid239_Out0_copy240_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid241_In0_c0 <= "" & bh7_w43_6_c0 & bh7_w43_5_c0 & bh7_w43_4_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid241_In1_c0 <= "" & bh7_w44_2_c0 & bh7_w44_4_c0;
   bh7_w43_9_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid241_Out0_c0(0);
   bh7_w44_5_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid241_Out0_c0(1);
   bh7_w45_4_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid241_Out0_c0(2);
   Compressor_23_3_Freq500_uid156_uid241: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid241_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid241_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid241_Out0_copy242_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid241_Out0_c0 <= Compressor_23_3_Freq500_uid156_bh7_uid241_Out0_copy242_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid243_In0_c0 <= "" & bh7_w45_3_c0 & bh7_w45_2_c0 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid243_In1_c0 <= "" & bh7_w46_2_c0;
   bh7_w45_5_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid243_Out0_c0(0);
   bh7_w46_3_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid243_Out0_c0(1);
   bh7_w47_1_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid243_Out0_c0(2);
   Compressor_14_3_Freq500_uid164_uid243: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid243_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid243_In1_c0,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid243_Out0_copy244_c0);
   Compressor_14_3_Freq500_uid164_bh7_uid243_Out0_c0 <= Compressor_14_3_Freq500_uid164_bh7_uid243_Out0_copy244_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid245_In0_c0 <= "" & bh7_w22_8_c0 & bh7_w22_7_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid245_In1_c0 <= "" & bh7_w23_10_c0 & bh7_w23_11_c0;
   bh7_w22_9_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_c1(0);
   bh7_w23_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_c1(1);
   bh7_w24_10_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid245: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid245_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid245_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_copy246_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid245_Out0_copy246_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid247_In0_c0 <= "" & bh7_w25_11_c0 & bh7_w25_10_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid247_In1_c0 <= "" & bh7_w26_7_c0 & bh7_w26_10_c0;
   bh7_w25_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_c1(0);
   bh7_w26_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_c1(1);
   bh7_w27_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid247: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid247_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid247_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_copy248_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid247_Out0_copy248_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid249_In0_c0 <= "" & bh7_w27_11_c0 & bh7_w27_10_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid249_In1_c0 <= "" & bh7_w28_7_c0 & bh7_w28_10_c0;
   bh7_w27_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_c1(0);
   bh7_w28_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_c1(1);
   bh7_w29_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid249: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid249_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid249_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_copy250_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid249_Out0_copy250_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid251_In0_c0 <= "" & bh7_w29_11_c0 & bh7_w29_10_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid251_In1_c0 <= "" & bh7_w30_7_c0 & bh7_w30_10_c0;
   bh7_w29_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_c1(0);
   bh7_w30_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_c1(1);
   bh7_w31_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid251: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid251_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid251_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_copy252_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid251_Out0_copy252_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid253_In0_c0 <= "" & bh7_w31_11_c0 & bh7_w31_10_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid253_In1_c0 <= "" & bh7_w32_7_c0 & bh7_w32_10_c0;
   bh7_w31_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_c1(0);
   bh7_w32_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_c1(1);
   bh7_w33_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid253: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid253_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid253_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_copy254_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid253_Out0_copy254_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid255_In0_c0 <= "" & bh7_w33_11_c0 & bh7_w33_10_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid255_In1_c0 <= "" & bh7_w34_7_c0 & bh7_w34_10_c0;
   bh7_w33_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_c1(0);
   bh7_w34_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_c1(1);
   bh7_w35_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid255: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid255_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid255_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_copy256_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid255_Out0_copy256_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid257_In0_c0 <= "" & bh7_w35_11_c0 & bh7_w35_10_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid257_In1_c0 <= "" & bh7_w36_7_c0 & bh7_w36_10_c0;
   bh7_w35_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_c1(0);
   bh7_w36_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_c1(1);
   bh7_w37_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid257: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid257_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid257_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_copy258_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid257_Out0_copy258_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid259_In0_c0 <= "" & bh7_w37_11_c0 & bh7_w37_10_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid259_In1_c0 <= "" & bh7_w38_7_c0 & bh7_w38_10_c0;
   bh7_w37_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_c1(0);
   bh7_w38_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_c1(1);
   bh7_w39_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid259: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid259_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid259_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_copy260_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid259_Out0_copy260_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid261_In0_c0 <= "" & bh7_w39_11_c0 & bh7_w39_10_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid261_In1_c0 <= "" & bh7_w40_7_c0 & bh7_w40_10_c0;
   bh7_w39_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_c1(0);
   bh7_w40_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_c1(1);
   bh7_w41_10_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid261: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid261_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid261_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_copy262_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid261_Out0_copy262_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid263_In0_c0 <= "" & bh7_w41_9_c0 & bh7_w41_8_c0 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid263_In1_c0 <= "" & bh7_w42_8_c0 & bh7_w42_9_c0;
   bh7_w41_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_c1(0);
   bh7_w42_10_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_c1(1);
   bh7_w43_10_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid263: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid263_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid263_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_copy264_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid263_Out0_copy264_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid265_In0_c0 <= "" & bh7_w43_7_c0 & bh7_w43_9_c0 & bh7_w43_8_c0;
   Compressor_23_3_Freq500_uid156_bh7_uid265_In1_c0 <= "" & bh7_w44_3_c0 & bh7_w44_5_c0;
   bh7_w43_11_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_c1(0);
   bh7_w44_6_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_c1(1);
   bh7_w45_6_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid265: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid265_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid265_In1_c0,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_copy266_c0);
   Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid265_Out0_copy266_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid267_In0_c0 <= "" & bh7_w45_5_c0 & bh7_w45_4_c0 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid267_In1_c0 <= "" & bh7_w46_3_c0;
   bh7_w45_7_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_c1(0);
   bh7_w46_4_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_c1(1);
   bh7_w47_2_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid267: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid267_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid267_In1_c0,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_copy268_c0);
   Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid267_Out0_copy268_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid160_bh7_uid269_In0_c0 <= "" & bh7_w47_0_c0 & bh7_w47_1_c0 & "0";
   bh7_w47_3_c1 <= Compressor_3_2_Freq500_uid160_bh7_uid269_Out0_c1(0);
   Compressor_3_2_Freq500_uid160_uid269: Compressor_3_2_Freq500_uid160
      port map ( X0 => Compressor_3_2_Freq500_uid160_bh7_uid269_In0_c0,
                 R => Compressor_3_2_Freq500_uid160_bh7_uid269_Out0_copy270_c0);
   Compressor_3_2_Freq500_uid160_bh7_uid269_Out0_c1 <= Compressor_3_2_Freq500_uid160_bh7_uid269_Out0_copy270_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid271_In0_c1 <= "" & bh7_w24_9_c1 & bh7_w24_10_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid271_In1_c1 <= "" & bh7_w25_12_c1;
   bh7_w24_11_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid271_Out0_c1(0);
   bh7_w25_13_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid271_Out0_c1(1);
   bh7_w26_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid271_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid271: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid271_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid271_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid271_Out0_copy272_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid271_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid271_Out0_copy272_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid273_In0_c1 <= "" & bh7_w27_13_c1 & bh7_w27_12_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid273_In1_c1 <= "" & bh7_w28_11_c1;
   bh7_w27_14_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid273_Out0_c1(0);
   bh7_w28_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid273_Out0_c1(1);
   bh7_w29_14_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid273_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid273: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid273_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid273_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid273_Out0_copy274_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid273_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid273_Out0_copy274_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid275_In0_c1 <= "" & bh7_w29_13_c1 & bh7_w29_12_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid275_In1_c1 <= "" & bh7_w30_11_c1;
   bh7_w29_15_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid275_Out0_c1(0);
   bh7_w30_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid275_Out0_c1(1);
   bh7_w31_14_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid275_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid275: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid275_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid275_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid275_Out0_copy276_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid275_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid275_Out0_copy276_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid277_In0_c1 <= "" & bh7_w31_13_c1 & bh7_w31_12_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid277_In1_c1 <= "" & bh7_w32_11_c1;
   bh7_w31_15_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid277_Out0_c1(0);
   bh7_w32_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid277_Out0_c1(1);
   bh7_w33_14_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid277_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid277: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid277_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid277_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid277_Out0_copy278_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid277_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid277_Out0_copy278_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid279_In0_c1 <= "" & bh7_w33_13_c1 & bh7_w33_12_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid279_In1_c1 <= "" & bh7_w34_11_c1;
   bh7_w33_15_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid279_Out0_c1(0);
   bh7_w34_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid279_Out0_c1(1);
   bh7_w35_14_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid279_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid279: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid279_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid279_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid279_Out0_copy280_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid279_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid279_Out0_copy280_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid281_In0_c1 <= "" & bh7_w35_13_c1 & bh7_w35_12_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid281_In1_c1 <= "" & bh7_w36_11_c1;
   bh7_w35_15_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid281_Out0_c1(0);
   bh7_w36_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid281_Out0_c1(1);
   bh7_w37_14_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid281_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid281: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid281_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid281_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid281_Out0_copy282_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid281_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid281_Out0_copy282_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid283_In0_c1 <= "" & bh7_w37_13_c1 & bh7_w37_12_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid283_In1_c1 <= "" & bh7_w38_11_c1;
   bh7_w37_15_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid283_Out0_c1(0);
   bh7_w38_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid283_Out0_c1(1);
   bh7_w39_14_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid283_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid283: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid283_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid283_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid283_Out0_copy284_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid283_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid283_Out0_copy284_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid285_In0_c1 <= "" & bh7_w39_13_c1 & bh7_w39_12_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid285_In1_c1 <= "" & bh7_w40_11_c1;
   bh7_w39_15_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid285_Out0_c1(0);
   bh7_w40_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid285_Out0_c1(1);
   bh7_w41_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid285_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid285: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid285_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid285_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid285_Out0_copy286_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid285_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid285_Out0_copy286_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid287_In0_c1 <= "" & bh7_w41_11_c1 & bh7_w41_10_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid287_In1_c1 <= "" & bh7_w42_10_c1;
   bh7_w41_13_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid287_Out0_c1(0);
   bh7_w42_11_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid287_Out0_c1(1);
   bh7_w43_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid287_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid287: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid287_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid287_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid287_Out0_copy288_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid287_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid287_Out0_copy288_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid289_In0_c1 <= "" & bh7_w43_10_c1 & bh7_w43_11_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid289_In1_c1 <= "" & bh7_w44_6_c1;
   bh7_w43_13_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid289_Out0_c1(0);
   bh7_w44_7_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid289_Out0_c1(1);
   bh7_w45_8_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid289_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid289: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid289_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid289_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid289_Out0_copy290_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid289_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid289_Out0_copy290_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid291_In0_c1 <= "" & bh7_w45_6_c1 & bh7_w45_7_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid291_In1_c1 <= "" & bh7_w46_4_c1;
   bh7_w45_9_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid291_Out0_c1(0);
   bh7_w46_5_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid291_Out0_c1(1);
   bh7_w47_4_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid291_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid291: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid291_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid291_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid291_Out0_copy292_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid291_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid291_Out0_copy292_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid293_In0_c1 <= "" & bh7_w47_3_c1 & bh7_w47_2_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid293_In1_c0 <= "" & "0";
   bh7_w47_5_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid293_Out0_c1(0);
   Compressor_14_3_Freq500_uid164_uid293: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid293_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid293_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid293_Out0_copy294_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid293_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid293_Out0_copy294_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid295_In0_c1 <= "" & bh7_w17_1_c1 & bh7_w17_0_c1 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid295_In1_c1 <= "" & bh7_w18_2_c1 & bh7_w18_0_c1;
   bh7_w17_2_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid295_Out0_c1(0);
   bh7_w18_3_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid295_Out0_c1(1);
   bh7_w19_4_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid295_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid295: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid295_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid295_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid295_Out0_copy296_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid295_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid295_Out0_copy296_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid297_In0_c1 <= "" & bh7_w19_3_c1 & bh7_w19_0_c1 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid297_In1_c1 <= "" & bh7_w20_6_c1 & bh7_w20_0_c1;
   bh7_w19_5_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid297_Out0_c1(0);
   bh7_w20_7_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid297_Out0_c1(1);
   bh7_w21_8_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid297_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid297: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid297_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid297_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid297_Out0_copy298_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid297_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid297_Out0_copy298_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid299_In0_c1 <= "" & bh7_w21_7_c1 & bh7_w21_0_c1 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid299_In1_c1 <= "" & bh7_w22_9_c1 & bh7_w22_0_c1;
   bh7_w21_9_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid299_Out0_c1(0);
   bh7_w22_10_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid299_Out0_c1(1);
   bh7_w23_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid299_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid299: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid299_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid299_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid299_Out0_copy300_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid299_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid299_Out0_copy300_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid301_In0_c1 <= "" & bh7_w23_12_c1 & bh7_w23_0_c1 & "0";
   Compressor_23_3_Freq500_uid156_bh7_uid301_In1_c1 <= "" & bh7_w24_11_c1 & bh7_w24_0_c1;
   bh7_w23_14_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid301_Out0_c1(0);
   bh7_w24_12_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid301_Out0_c1(1);
   bh7_w25_14_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid301_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid301: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid301_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid301_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid301_Out0_copy302_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid301_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid301_Out0_copy302_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid160_bh7_uid303_In0_c1 <= "" & bh7_w25_13_c1 & bh7_w25_0_c1 & "0";
   bh7_w25_15_c1 <= Compressor_3_2_Freq500_uid160_bh7_uid303_Out0_c1(0);
   bh7_w26_13_c1 <= Compressor_3_2_Freq500_uid160_bh7_uid303_Out0_c1(1);
   Compressor_3_2_Freq500_uid160_uid303: Compressor_3_2_Freq500_uid160
      port map ( X0 => Compressor_3_2_Freq500_uid160_bh7_uid303_In0_c1,
                 R => Compressor_3_2_Freq500_uid160_bh7_uid303_Out0_copy304_c1);
   Compressor_3_2_Freq500_uid160_bh7_uid303_Out0_c1 <= Compressor_3_2_Freq500_uid160_bh7_uid303_Out0_copy304_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid305_In0_c1 <= "" & bh7_w26_11_c1 & bh7_w26_12_c1 & bh7_w26_0_c1;
   Compressor_23_3_Freq500_uid156_bh7_uid305_In1_c1 <= "" & bh7_w27_14_c1 & bh7_w27_0_c1;
   bh7_w26_14_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid305_Out0_c1(0);
   bh7_w27_15_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid305_Out0_c1(1);
   bh7_w28_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid305_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid305: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid305_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid305_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid305_Out0_copy306_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid305_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid305_Out0_copy306_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid160_bh7_uid307_In0_c1 <= "" & bh7_w28_12_c1 & bh7_w28_0_c1 & "0";
   bh7_w28_14_c1 <= Compressor_3_2_Freq500_uid160_bh7_uid307_Out0_c1(0);
   bh7_w29_16_c1 <= Compressor_3_2_Freq500_uid160_bh7_uid307_Out0_c1(1);
   Compressor_3_2_Freq500_uid160_uid307: Compressor_3_2_Freq500_uid160
      port map ( X0 => Compressor_3_2_Freq500_uid160_bh7_uid307_In0_c1,
                 R => Compressor_3_2_Freq500_uid160_bh7_uid307_Out0_copy308_c1);
   Compressor_3_2_Freq500_uid160_bh7_uid307_Out0_c1 <= Compressor_3_2_Freq500_uid160_bh7_uid307_Out0_copy308_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid309_In0_c1 <= "" & bh7_w29_15_c1 & bh7_w29_14_c1 & bh7_w29_0_c1;
   Compressor_23_3_Freq500_uid156_bh7_uid309_In1_c1 <= "" & bh7_w30_12_c1 & bh7_w30_0_c1;
   bh7_w29_17_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid309_Out0_c1(0);
   bh7_w30_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid309_Out0_c1(1);
   bh7_w31_16_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid309_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid309: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid309_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid309_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid309_Out0_copy310_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid309_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid309_Out0_copy310_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid311_In0_c1 <= "" & bh7_w31_15_c1 & bh7_w31_14_c1 & bh7_w31_0_c1;
   Compressor_23_3_Freq500_uid156_bh7_uid311_In1_c1 <= "" & bh7_w32_12_c1 & bh7_w32_0_c1;
   bh7_w31_17_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid311_Out0_c1(0);
   bh7_w32_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid311_Out0_c1(1);
   bh7_w33_16_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid311_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid311: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid311_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid311_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid311_Out0_copy312_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid311_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid311_Out0_copy312_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid313_In0_c1 <= "" & bh7_w33_15_c1 & bh7_w33_14_c1 & bh7_w33_0_c1;
   Compressor_23_3_Freq500_uid156_bh7_uid313_In1_c1 <= "" & bh7_w34_12_c1 & bh7_w34_0_c1;
   bh7_w33_17_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid313_Out0_c1(0);
   bh7_w34_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid313_Out0_c1(1);
   bh7_w35_16_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid313_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid313: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid313_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid313_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid313_Out0_copy314_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid313_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid313_Out0_copy314_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid315_In0_c1 <= "" & bh7_w35_15_c1 & bh7_w35_14_c1 & bh7_w35_0_c1;
   Compressor_23_3_Freq500_uid156_bh7_uid315_In1_c1 <= "" & bh7_w36_12_c1 & bh7_w36_0_c1;
   bh7_w35_17_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid315_Out0_c1(0);
   bh7_w36_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid315_Out0_c1(1);
   bh7_w37_16_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid315_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid315: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid315_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid315_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid315_Out0_copy316_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid315_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid315_Out0_copy316_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid317_In0_c1 <= "" & bh7_w37_15_c1 & bh7_w37_14_c1 & bh7_w37_0_c1;
   Compressor_23_3_Freq500_uid156_bh7_uid317_In1_c1 <= "" & bh7_w38_12_c1 & bh7_w38_0_c1;
   bh7_w37_17_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid317_Out0_c1(0);
   bh7_w38_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid317_Out0_c1(1);
   bh7_w39_16_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid317_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid317: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid317_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid317_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid317_Out0_copy318_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid317_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid317_Out0_copy318_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid156_bh7_uid319_In0_c1 <= "" & bh7_w39_15_c1 & bh7_w39_14_c1 & bh7_w39_0_c1;
   Compressor_23_3_Freq500_uid156_bh7_uid319_In1_c1 <= "" & bh7_w40_12_c1 & bh7_w40_0_c1;
   bh7_w39_17_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid319_Out0_c1(0);
   bh7_w40_13_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid319_Out0_c1(1);
   bh7_w41_14_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid319_Out0_c1(2);
   Compressor_23_3_Freq500_uid156_uid319: Compressor_23_3_Freq500_uid156
      port map ( X0 => Compressor_23_3_Freq500_uid156_bh7_uid319_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid156_bh7_uid319_In1_c1,
                 R => Compressor_23_3_Freq500_uid156_bh7_uid319_Out0_copy320_c1);
   Compressor_23_3_Freq500_uid156_bh7_uid319_Out0_c1 <= Compressor_23_3_Freq500_uid156_bh7_uid319_Out0_copy320_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid321_In0_c1 <= "" & bh7_w41_13_c1 & bh7_w41_12_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid321_In1_c1 <= "" & bh7_w42_11_c1;
   bh7_w41_15_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid321_Out0_c1(0);
   bh7_w42_12_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid321_Out0_c1(1);
   bh7_w43_14_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid321_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid321: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid321_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid321_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid321_Out0_copy322_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid321_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid321_Out0_copy322_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid323_In0_c1 <= "" & bh7_w43_12_c1 & bh7_w43_13_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid323_In1_c1 <= "" & bh7_w44_7_c1;
   bh7_w43_15_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid323_Out0_c1(0);
   bh7_w44_8_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid323_Out0_c1(1);
   bh7_w45_10_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid323_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid323: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid323_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid323_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid323_Out0_copy324_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid323_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid323_Out0_copy324_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid325_In0_c1 <= "" & bh7_w45_8_c1 & bh7_w45_9_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid325_In1_c1 <= "" & bh7_w46_5_c1;
   bh7_w45_11_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid325_Out0_c1(0);
   bh7_w46_6_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid325_Out0_c1(1);
   bh7_w47_6_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid325_Out0_c1(2);
   Compressor_14_3_Freq500_uid164_uid325: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid325_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid325_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid325_Out0_copy326_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid325_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid325_Out0_copy326_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid164_bh7_uid327_In0_c1 <= "" & bh7_w47_4_c1 & bh7_w47_5_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid164_bh7_uid327_In1_c0 <= "" & "0";
   bh7_w47_7_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid327_Out0_c1(0);
   Compressor_14_3_Freq500_uid164_uid327: Compressor_14_3_Freq500_uid164
      port map ( X0 => Compressor_14_3_Freq500_uid164_bh7_uid327_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid164_bh7_uid327_In1_c1,
                 R => Compressor_14_3_Freq500_uid164_bh7_uid327_Out0_copy328_c1);
   Compressor_14_3_Freq500_uid164_bh7_uid327_Out0_c1 <= Compressor_14_3_Freq500_uid164_bh7_uid327_Out0_copy328_c1; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh7_18_c1 <= bh7_w18_3_c1 & bh7_w17_2_c1 & bh7_w16_0_c1 & bh7_w15_0_c1 & bh7_w14_0_c1 & bh7_w13_0_c1 & bh7_w12_0_c1 & bh7_w11_0_c1 & bh7_w10_0_c1 & bh7_w9_0_c1 & bh7_w8_0_c1 & bh7_w7_0_c1 & bh7_w6_0_c1 & bh7_w5_0_c1 & bh7_w4_0_c1 & bh7_w3_0_c1 & bh7_w2_0_c1 & bh7_w1_0_c1 & bh7_w0_0_c1;

   bitheapFinalAdd_bh7_In0_c1 <= "0" & bh7_w47_6_c1 & bh7_w46_6_c1 & bh7_w45_10_c1 & bh7_w44_8_c1 & bh7_w43_14_c1 & bh7_w42_12_c1 & bh7_w41_15_c1 & bh7_w40_13_c1 & bh7_w39_17_c1 & bh7_w38_13_c1 & bh7_w37_17_c1 & bh7_w36_13_c1 & bh7_w35_17_c1 & bh7_w34_13_c1 & bh7_w33_17_c1 & bh7_w32_13_c1 & bh7_w31_17_c1 & bh7_w30_13_c1 & bh7_w29_17_c1 & bh7_w28_14_c1 & bh7_w27_15_c1 & bh7_w26_14_c1 & bh7_w25_15_c1 & bh7_w24_12_c1 & bh7_w23_14_c1 & bh7_w22_10_c1 & bh7_w21_9_c1 & bh7_w20_7_c1 & bh7_w19_5_c1;
   bitheapFinalAdd_bh7_In1_c1 <= "0" & bh7_w47_7_c1 & "0" & bh7_w45_11_c1 & "0" & bh7_w43_15_c1 & "0" & bh7_w41_14_c1 & "0" & bh7_w39_16_c1 & "0" & bh7_w37_16_c1 & "0" & bh7_w35_16_c1 & "0" & bh7_w33_16_c1 & "0" & bh7_w31_16_c1 & "0" & bh7_w29_16_c1 & bh7_w28_13_c1 & "0" & bh7_w26_13_c1 & bh7_w25_14_c1 & "0" & bh7_w23_13_c1 & "0" & bh7_w21_8_c1 & "0" & bh7_w19_4_c1;
   bitheapFinalAdd_bh7_Cin_c0 <= '0';

   bitheapFinalAdd_bh7: IntAdder_30_Freq500_uid330
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 Cin => bitheapFinalAdd_bh7_Cin_c0,
                 X => bitheapFinalAdd_bh7_In0_c1,
                 Y => bitheapFinalAdd_bh7_In1_c1,
                 R => bitheapFinalAdd_bh7_Out_c2);
   bitheapResult_bh7_c2 <= bitheapFinalAdd_bh7_Out_c2(28 downto 0) & tmp_bitheapResult_bh7_18_c2;
   R <= bitheapResult_bh7_c2(47 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_Freq500_uid333
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_Freq500_uid333 is
    port (clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(32 downto 0);
          Y : in  std_logic_vector(32 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_Freq500_uid333 is
signal Cin_1_c3, Cin_1_c4 :  std_logic;
signal X_1_c2, X_1_c3, X_1_c4 :  std_logic_vector(33 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3, Y_1_c4 :  std_logic_vector(33 downto 0);
signal S_1_c4 :  std_logic_vector(33 downto 0);
signal R_1_c4 :  std_logic_vector(32 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_1_c1 <= Y_1_c0;
            end if;
            if ce_2 = '1' then
               Y_1_c2 <= Y_1_c1;
            end if;
            if ce_3 = '1' then
               X_1_c3 <= X_1_c2;
               Y_1_c3 <= Y_1_c2;
            end if;
            if ce_4 = '1' then
               Cin_1_c4 <= Cin_1_c3;
               X_1_c4 <= X_1_c3;
               Y_1_c4 <= Y_1_c3;
            end if;
         end if;
      end process;
   Cin_1_c3 <= Cin;
   X_1_c2 <= '0' & X(32 downto 0);
   Y_1_c0 <= '0' & Y(32 downto 0);
   S_1_c4 <= X_1_c4 + Y_1_c4 + Cin_1_c4;
   R_1_c4 <= S_1_c4(32 downto 0);
   R <= R_1_c4 ;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointMultiplier
--                      (FPMult_8_23_uid2_Freq500_uid3)
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointMultiplier_32_2_783000 is
    port (clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointMultiplier_32_2_783000 is
   component IntMultiplier_24x24_48_Freq500_uid5 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_Freq500_uid333 is
      port ( clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
             X : in  std_logic_vector(32 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(32 downto 0)   );
   end component;

signal sign_c0, sign_c1, sign_c2, sign_c3, sign_c4 :  std_logic;
signal expX_c0 :  std_logic_vector(7 downto 0);
signal expY_c0 :  std_logic_vector(7 downto 0);
signal expSumPreSub_c0, expSumPreSub_c1 :  std_logic_vector(9 downto 0);
signal bias_c0, bias_c1 :  std_logic_vector(9 downto 0);
signal expSum_c1, expSum_c2 :  std_logic_vector(9 downto 0);
signal sigX_c0 :  std_logic_vector(23 downto 0);
signal sigY_c0 :  std_logic_vector(23 downto 0);
signal sigProd_c2 :  std_logic_vector(47 downto 0);
signal excSel_c0 :  std_logic_vector(3 downto 0);
signal exc_c0, exc_c1, exc_c2, exc_c3, exc_c4 :  std_logic_vector(1 downto 0);
signal norm_c2 :  std_logic;
signal expPostNorm_c2 :  std_logic_vector(9 downto 0);
signal sigProdExt_c2, sigProdExt_c3 :  std_logic_vector(47 downto 0);
signal expSig_c2 :  std_logic_vector(32 downto 0);
signal sticky_c2, sticky_c3 :  std_logic;
signal guard_c3 :  std_logic;
signal round_c3 :  std_logic;
signal expSigPostRound_c4 :  std_logic_vector(32 downto 0);
signal excPostNorm_c4 :  std_logic_vector(1 downto 0);
signal finalExc_c4 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               sign_c1 <= sign_c0;
               expSumPreSub_c1 <= expSumPreSub_c0;
               bias_c1 <= bias_c0;
               exc_c1 <= exc_c0;
            end if;
            if ce_2 = '1' then
               sign_c2 <= sign_c1;
               expSum_c2 <= expSum_c1;
               exc_c2 <= exc_c1;
            end if;
            if ce_3 = '1' then
               sign_c3 <= sign_c2;
               exc_c3 <= exc_c2;
               sigProdExt_c3 <= sigProdExt_c2;
               sticky_c3 <= sticky_c2;
            end if;
            if ce_4 = '1' then
               sign_c4 <= sign_c3;
               exc_c4 <= exc_c3;
            end if;
         end if;
      end process;
   sign_c0 <= X(31) xor Y(31);
   expX_c0 <= X(30 downto 23);
   expY_c0 <= Y(30 downto 23);
   expSumPreSub_c0 <= ("00" & expX_c0) + ("00" & expY_c0);
   bias_c0 <= CONV_STD_LOGIC_VECTOR(127,10);
   expSum_c1 <= expSumPreSub_c1 - bias_c1;
   sigX_c0 <= "1" & X(22 downto 0);
   sigY_c0 <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_24x24_48_Freq500_uid5
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => sigX_c0,
                 Y => sigY_c0,
                 R => sigProd_c2);
   excSel_c0 <= X(33 downto 32) & Y(33 downto 32);
   with excSel_c0  select  
   exc_c0 <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm_c2 <= sigProd_c2(47);
   -- exponent update
   expPostNorm_c2 <= expSum_c2 + ("000000000" & norm_c2);
   -- significand normalization shift
   sigProdExt_c2 <= sigProd_c2(46 downto 0) & "0" when norm_c2='1' else
                         sigProd_c2(45 downto 0) & "00";
   expSig_c2 <= expPostNorm_c2 & sigProdExt_c2(47 downto 25);
   sticky_c2 <= sigProdExt_c2(24);
   guard_c3 <= '0' when sigProdExt_c3(23 downto 0)="000000000000000000000000" else '1';
   round_c3 <= sticky_c3 and ( (guard_c3 and not(sigProdExt_c3(25))) or (sigProdExt_c3(25) ))  ;
   RoundingAdder: IntAdder_33_Freq500_uid333
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 Cin => round_c3,
                 X => expSig_c2,
                 Y => "000000000000000000000000000000000",
                 R => expSigPostRound_c4);
   with expSigPostRound_c4(32 downto 31)  select 
   excPostNorm_c4 <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_c4  select  
   finalExc_c4 <= exc_c4 when  "11"|"10"|"00",
                       excPostNorm_c4 when others; 
   R <= finalExc_c4 & sign_c4 & expSigPostRound_c4(30 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid15
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid15 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid15 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid20
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid20 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid20 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid27
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid27 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid27 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid32
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid32 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid32 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid39
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid39 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid39 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid44
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid44 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid44 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid51
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid51 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid51 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid56
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid56 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid56 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid63
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid63 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid63 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid68
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid68 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid68 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid75
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid75 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid75 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid80
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid80 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid80 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid87
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid87 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid87 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid92
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid92 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid92 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid99
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid99 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid99 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid104
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid104 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid104 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid111
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid111 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid111 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid116
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid116 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid116 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid123
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid128
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid128 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid128 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid135
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid135 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid135 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid140
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid140 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid140 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid147
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid147 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid147 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid152
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid152 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid152 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq300_uid156
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid156 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid156 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid160
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid160 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid160 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq300_uid164
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid164 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid164 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid170
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid170 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid170 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid9
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid9 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid9 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq300_uid11
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid11 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid11 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid13
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid13 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid13 is
   component MultTable_Freq300_uid15 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy16_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid15
      port map ( X => Xtable_c0,
                 Y => Y1_copy16_c0);
   Y1_c0 <= Y1_copy16_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid18
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid18 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid18 is
   component MultTable_Freq300_uid20 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy21_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid20
      port map ( X => Xtable_c0,
                 Y => Y1_copy21_c0);
   Y1_c0 <= Y1_copy21_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq300_uid23
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid23 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid23 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid25
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid25 is
   component MultTable_Freq300_uid27 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy28_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid27
      port map ( X => Xtable_c0,
                 Y => Y1_copy28_c0);
   Y1_c0 <= Y1_copy28_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid30
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid30 is
   component MultTable_Freq300_uid32 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy33_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid32
      port map ( X => Xtable_c0,
                 Y => Y1_copy33_c0);
   Y1_c0 <= Y1_copy33_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq300_uid35
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid35 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid35 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid37
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid37 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid37 is
   component MultTable_Freq300_uid39 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy40_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid39
      port map ( X => Xtable_c0,
                 Y => Y1_copy40_c0);
   Y1_c0 <= Y1_copy40_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid42
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid42 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid42 is
   component MultTable_Freq300_uid44 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy45_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid44
      port map ( X => Xtable_c0,
                 Y => Y1_copy45_c0);
   Y1_c0 <= Y1_copy45_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq300_uid47
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid47 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid47 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid49
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid49 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid49 is
   component MultTable_Freq300_uid51 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy52_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid51
      port map ( X => Xtable_c0,
                 Y => Y1_copy52_c0);
   Y1_c0 <= Y1_copy52_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid54
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid54 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid54 is
   component MultTable_Freq300_uid56 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy57_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid56
      port map ( X => Xtable_c0,
                 Y => Y1_copy57_c0);
   Y1_c0 <= Y1_copy57_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq300_uid59
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid59 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid59 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid61
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid61 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid61 is
   component MultTable_Freq300_uid63 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy64_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid63
      port map ( X => Xtable_c0,
                 Y => Y1_copy64_c0);
   Y1_c0 <= Y1_copy64_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid66
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid66 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid66 is
   component MultTable_Freq300_uid68 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy69_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid68
      port map ( X => Xtable_c0,
                 Y => Y1_copy69_c0);
   Y1_c0 <= Y1_copy69_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq300_uid71
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid71 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid73
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid73 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid73 is
   component MultTable_Freq300_uid75 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy76_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid75
      port map ( X => Xtable_c0,
                 Y => Y1_copy76_c0);
   Y1_c0 <= Y1_copy76_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid78
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid78 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid78 is
   component MultTable_Freq300_uid80 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy81_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid80
      port map ( X => Xtable_c0,
                 Y => Y1_copy81_c0);
   Y1_c0 <= Y1_copy81_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq300_uid83
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid83 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid83 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid85
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid85 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid85 is
   component MultTable_Freq300_uid87 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy88_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid87
      port map ( X => Xtable_c0,
                 Y => Y1_copy88_c0);
   Y1_c0 <= Y1_copy88_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid90
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid90 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid90 is
   component MultTable_Freq300_uid92 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy93_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid92
      port map ( X => Xtable_c0,
                 Y => Y1_copy93_c0);
   Y1_c0 <= Y1_copy93_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_1x2_Freq300_uid95
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid95 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid95 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_3x2_Freq300_uid97
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid97 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid97 is
   component MultTable_Freq300_uid99 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy100_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid99
      port map ( X => Xtable_c0,
                 Y => Y1_copy100_c0);
   Y1_c0 <= Y1_copy100_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid102
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid102 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid102 is
   component MultTable_Freq300_uid104 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy105_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid104
      port map ( X => Xtable_c0,
                 Y => Y1_copy105_c0);
   Y1_c0 <= Y1_copy105_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq300_uid107
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid107 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid107 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid109
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid109 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid109 is
   component MultTable_Freq300_uid111 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy112_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid111
      port map ( X => Xtable_c0,
                 Y => Y1_copy112_c0);
   Y1_c0 <= Y1_copy112_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid114
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid114 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid114 is
   component MultTable_Freq300_uid116 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy117_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid116
      port map ( X => Xtable_c0,
                 Y => Y1_copy117_c0);
   Y1_c0 <= Y1_copy117_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq300_uid119
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid119 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid119 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid121
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid121 is
   component MultTable_Freq300_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy124_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid123
      port map ( X => Xtable_c0,
                 Y => Y1_copy124_c0);
   Y1_c0 <= Y1_copy124_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid126
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid126 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid126 is
   component MultTable_Freq300_uid128 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy129_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid128
      port map ( X => Xtable_c0,
                 Y => Y1_copy129_c0);
   Y1_c0 <= Y1_copy129_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq300_uid131
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid131 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid131 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid133
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid133 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid133 is
   component MultTable_Freq300_uid135 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy136_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid135
      port map ( X => Xtable_c0,
                 Y => Y1_copy136_c0);
   Y1_c0 <= Y1_copy136_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid138
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid138 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid138 is
   component MultTable_Freq300_uid140 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy141_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid140
      port map ( X => Xtable_c0,
                 Y => Y1_copy141_c0);
   Y1_c0 <= Y1_copy141_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x2_Freq300_uid143
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x2_Freq300_uid143 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x2_Freq300_uid143 is
signal replicated_c0 :  std_logic_vector(1 downto 0);
signal prod_c0 :  std_logic_vector(1 downto 0);
begin
   replicated_c0 <= (1 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid145
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid145 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid145 is
   component MultTable_Freq300_uid147 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy148_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid147
      port map ( X => Xtable_c0,
                 Y => Y1_copy148_c0);
   Y1_c0 <= Y1_copy148_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid150
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid150 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid150 is
   component MultTable_Freq300_uid152 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy153_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid152
      port map ( X => Xtable_c0,
                 Y => Y1_copy153_c0);
   Y1_c0 <= Y1_copy153_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_30_Freq300_uid352
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_30_Freq300_uid352 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(29 downto 0);
          Y : in  std_logic_vector(29 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of IntAdder_30_Freq300_uid352 is
signal Rtmp_c1 :  std_logic_vector(29 downto 0);
signal Cin_c1 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
         end if;
      end process;
   Rtmp_c1 <= X + Y + Cin_c1;
   R <= Rtmp_c1;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_24x24_48_Freq300_uid5
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_24x24_48_Freq300_uid5 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of IntMultiplier_24x24_48_Freq300_uid5 is
   component DSPBlock_17x24_Freq300_uid9 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid11 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid13 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid18 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid23 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid35 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid37 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid42 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid47 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid49 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid54 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid59 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid61 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid66 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid73 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid78 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid83 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid85 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid90 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid95 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid97 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid102 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid107 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid109 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid114 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid119 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid126 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid131 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid133 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid138 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x2_Freq300_uid143 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid145 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid150 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid156 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid160 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid164 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid170 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_30_Freq300_uid352 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(29 downto 0);
             Y : in  std_logic_vector(29 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(29 downto 0)   );
   end component;

signal XX_m6_c0 :  std_logic_vector(23 downto 0);
signal YY_m6_c0 :  std_logic_vector(23 downto 0);
signal tile_0_X_c0 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_0_output_c0 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w0_0_c0, bh7_w0_0_c1 :  std_logic;
signal bh7_w1_0_c0, bh7_w1_0_c1 :  std_logic;
signal bh7_w2_0_c0, bh7_w2_0_c1 :  std_logic;
signal bh7_w3_0_c0, bh7_w3_0_c1 :  std_logic;
signal bh7_w4_0_c0, bh7_w4_0_c1 :  std_logic;
signal bh7_w5_0_c0, bh7_w5_0_c1 :  std_logic;
signal bh7_w6_0_c0, bh7_w6_0_c1 :  std_logic;
signal bh7_w7_0_c0, bh7_w7_0_c1 :  std_logic;
signal bh7_w8_0_c0, bh7_w8_0_c1 :  std_logic;
signal bh7_w9_0_c0, bh7_w9_0_c1 :  std_logic;
signal bh7_w10_0_c0, bh7_w10_0_c1 :  std_logic;
signal bh7_w11_0_c0, bh7_w11_0_c1 :  std_logic;
signal bh7_w12_0_c0, bh7_w12_0_c1 :  std_logic;
signal bh7_w13_0_c0, bh7_w13_0_c1 :  std_logic;
signal bh7_w14_0_c0, bh7_w14_0_c1 :  std_logic;
signal bh7_w15_0_c0, bh7_w15_0_c1 :  std_logic;
signal bh7_w16_0_c0, bh7_w16_0_c1 :  std_logic;
signal bh7_w17_0_c0 :  std_logic;
signal bh7_w18_0_c0 :  std_logic;
signal bh7_w19_0_c0 :  std_logic;
signal bh7_w20_0_c0 :  std_logic;
signal bh7_w21_0_c0 :  std_logic;
signal bh7_w22_0_c0 :  std_logic;
signal bh7_w23_0_c0 :  std_logic;
signal bh7_w24_0_c0 :  std_logic;
signal bh7_w25_0_c0 :  std_logic;
signal bh7_w26_0_c0, bh7_w26_0_c1 :  std_logic;
signal bh7_w27_0_c0, bh7_w27_0_c1 :  std_logic;
signal bh7_w28_0_c0, bh7_w28_0_c1 :  std_logic;
signal bh7_w29_0_c0, bh7_w29_0_c1 :  std_logic;
signal bh7_w30_0_c0, bh7_w30_0_c1 :  std_logic;
signal bh7_w31_0_c0, bh7_w31_0_c1 :  std_logic;
signal bh7_w32_0_c0, bh7_w32_0_c1 :  std_logic;
signal bh7_w33_0_c0, bh7_w33_0_c1 :  std_logic;
signal bh7_w34_0_c0, bh7_w34_0_c1 :  std_logic;
signal bh7_w35_0_c0, bh7_w35_0_c1 :  std_logic;
signal bh7_w36_0_c0, bh7_w36_0_c1 :  std_logic;
signal bh7_w37_0_c0, bh7_w37_0_c1 :  std_logic;
signal bh7_w38_0_c0, bh7_w38_0_c1 :  std_logic;
signal bh7_w39_0_c0, bh7_w39_0_c1 :  std_logic;
signal bh7_w40_0_c0, bh7_w40_0_c1 :  std_logic;
signal tile_1_X_c0 :  std_logic_vector(0 downto 0);
signal tile_1_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_1_output_c0 :  std_logic_vector(1 downto 0);
signal tile_1_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w45_0_c0 :  std_logic;
signal bh7_w46_0_c0 :  std_logic;
signal tile_2_X_c0 :  std_logic_vector(2 downto 0);
signal tile_2_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_2_output_c0 :  std_logic_vector(4 downto 0);
signal tile_2_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w42_0_c0 :  std_logic;
signal bh7_w43_0_c0 :  std_logic;
signal bh7_w44_0_c0 :  std_logic;
signal bh7_w45_1_c0 :  std_logic;
signal bh7_w46_1_c0 :  std_logic;
signal tile_3_X_c0 :  std_logic_vector(2 downto 0);
signal tile_3_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_3_output_c0 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w39_1_c0 :  std_logic;
signal bh7_w40_1_c0 :  std_logic;
signal bh7_w41_0_c0 :  std_logic;
signal bh7_w42_1_c0 :  std_logic;
signal bh7_w43_1_c0 :  std_logic;
signal tile_4_X_c0 :  std_logic_vector(0 downto 0);
signal tile_4_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_4_output_c0 :  std_logic_vector(1 downto 0);
signal tile_4_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w43_2_c0 :  std_logic;
signal bh7_w44_1_c0 :  std_logic;
signal tile_5_X_c0 :  std_logic_vector(2 downto 0);
signal tile_5_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_5_output_c0 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w40_2_c0 :  std_logic;
signal bh7_w41_1_c0 :  std_logic;
signal bh7_w42_2_c0 :  std_logic;
signal bh7_w43_3_c0 :  std_logic;
signal bh7_w44_2_c0 :  std_logic;
signal tile_6_X_c0 :  std_logic_vector(2 downto 0);
signal tile_6_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_6_output_c0 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w37_1_c0 :  std_logic;
signal bh7_w38_1_c0 :  std_logic;
signal bh7_w39_2_c0 :  std_logic;
signal bh7_w40_3_c0 :  std_logic;
signal bh7_w41_2_c0 :  std_logic;
signal tile_7_X_c0 :  std_logic_vector(0 downto 0);
signal tile_7_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_7_output_c0 :  std_logic_vector(1 downto 0);
signal tile_7_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w41_3_c0 :  std_logic;
signal bh7_w42_3_c0 :  std_logic;
signal tile_8_X_c0 :  std_logic_vector(2 downto 0);
signal tile_8_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_8_output_c0 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w38_2_c0 :  std_logic;
signal bh7_w39_3_c0 :  std_logic;
signal bh7_w40_4_c0 :  std_logic;
signal bh7_w41_4_c0 :  std_logic;
signal bh7_w42_4_c0 :  std_logic;
signal tile_9_X_c0 :  std_logic_vector(2 downto 0);
signal tile_9_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_9_output_c0 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w35_1_c0 :  std_logic;
signal bh7_w36_1_c0 :  std_logic;
signal bh7_w37_2_c0 :  std_logic;
signal bh7_w38_3_c0 :  std_logic;
signal bh7_w39_4_c0 :  std_logic;
signal tile_10_X_c0 :  std_logic_vector(0 downto 0);
signal tile_10_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_10_output_c0 :  std_logic_vector(1 downto 0);
signal tile_10_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w39_5_c0 :  std_logic;
signal bh7_w40_5_c0 :  std_logic;
signal tile_11_X_c0 :  std_logic_vector(2 downto 0);
signal tile_11_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_11_output_c0 :  std_logic_vector(4 downto 0);
signal tile_11_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w36_2_c0 :  std_logic;
signal bh7_w37_3_c0 :  std_logic;
signal bh7_w38_4_c0 :  std_logic;
signal bh7_w39_6_c0 :  std_logic;
signal bh7_w40_6_c0 :  std_logic;
signal tile_12_X_c0 :  std_logic_vector(2 downto 0);
signal tile_12_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_12_output_c0 :  std_logic_vector(4 downto 0);
signal tile_12_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w33_1_c0 :  std_logic;
signal bh7_w34_1_c0 :  std_logic;
signal bh7_w35_2_c0 :  std_logic;
signal bh7_w36_3_c0 :  std_logic;
signal bh7_w37_4_c0 :  std_logic;
signal tile_13_X_c0 :  std_logic_vector(0 downto 0);
signal tile_13_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_13_output_c0 :  std_logic_vector(1 downto 0);
signal tile_13_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w37_5_c0 :  std_logic;
signal bh7_w38_5_c0 :  std_logic;
signal tile_14_X_c0 :  std_logic_vector(2 downto 0);
signal tile_14_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_14_output_c0 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w34_2_c0 :  std_logic;
signal bh7_w35_3_c0 :  std_logic;
signal bh7_w36_4_c0 :  std_logic;
signal bh7_w37_6_c0 :  std_logic;
signal bh7_w38_6_c0 :  std_logic;
signal tile_15_X_c0 :  std_logic_vector(2 downto 0);
signal tile_15_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_15_output_c0 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w31_1_c0 :  std_logic;
signal bh7_w32_1_c0 :  std_logic;
signal bh7_w33_2_c0 :  std_logic;
signal bh7_w34_3_c0 :  std_logic;
signal bh7_w35_4_c0 :  std_logic;
signal tile_16_X_c0 :  std_logic_vector(0 downto 0);
signal tile_16_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_16_output_c0 :  std_logic_vector(1 downto 0);
signal tile_16_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w35_5_c0 :  std_logic;
signal bh7_w36_5_c0 :  std_logic;
signal tile_17_X_c0 :  std_logic_vector(2 downto 0);
signal tile_17_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_17_output_c0 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w32_2_c0 :  std_logic;
signal bh7_w33_3_c0 :  std_logic;
signal bh7_w34_4_c0 :  std_logic;
signal bh7_w35_6_c0 :  std_logic;
signal bh7_w36_6_c0 :  std_logic;
signal tile_18_X_c0 :  std_logic_vector(2 downto 0);
signal tile_18_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_18_output_c0 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w29_1_c0 :  std_logic;
signal bh7_w30_1_c0 :  std_logic;
signal bh7_w31_2_c0 :  std_logic;
signal bh7_w32_3_c0 :  std_logic;
signal bh7_w33_4_c0 :  std_logic;
signal tile_19_X_c0 :  std_logic_vector(0 downto 0);
signal tile_19_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_19_output_c0 :  std_logic_vector(1 downto 0);
signal tile_19_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w33_5_c0 :  std_logic;
signal bh7_w34_5_c0 :  std_logic;
signal tile_20_X_c0 :  std_logic_vector(2 downto 0);
signal tile_20_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_20_output_c0 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w30_2_c0 :  std_logic;
signal bh7_w31_3_c0 :  std_logic;
signal bh7_w32_4_c0 :  std_logic;
signal bh7_w33_6_c0 :  std_logic;
signal bh7_w34_6_c0 :  std_logic;
signal tile_21_X_c0 :  std_logic_vector(2 downto 0);
signal tile_21_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_21_output_c0 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w27_1_c0 :  std_logic;
signal bh7_w28_1_c0 :  std_logic;
signal bh7_w29_2_c0 :  std_logic;
signal bh7_w30_3_c0 :  std_logic;
signal bh7_w31_4_c0 :  std_logic;
signal tile_22_X_c0 :  std_logic_vector(0 downto 0);
signal tile_22_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_22_output_c0 :  std_logic_vector(1 downto 0);
signal tile_22_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w31_5_c0 :  std_logic;
signal bh7_w32_5_c0 :  std_logic;
signal tile_23_X_c0 :  std_logic_vector(2 downto 0);
signal tile_23_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_23_output_c0 :  std_logic_vector(4 downto 0);
signal tile_23_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w28_2_c0 :  std_logic;
signal bh7_w29_3_c0 :  std_logic;
signal bh7_w30_4_c0 :  std_logic;
signal bh7_w31_6_c0 :  std_logic;
signal bh7_w32_6_c0 :  std_logic;
signal tile_24_X_c0 :  std_logic_vector(2 downto 0);
signal tile_24_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_24_output_c0 :  std_logic_vector(4 downto 0);
signal tile_24_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w25_1_c0 :  std_logic;
signal bh7_w26_1_c0 :  std_logic;
signal bh7_w27_2_c0 :  std_logic;
signal bh7_w28_3_c0 :  std_logic;
signal bh7_w29_4_c0 :  std_logic;
signal tile_25_X_c0 :  std_logic_vector(0 downto 0);
signal tile_25_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_25_output_c0 :  std_logic_vector(1 downto 0);
signal tile_25_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w29_5_c0 :  std_logic;
signal bh7_w30_5_c0 :  std_logic;
signal tile_26_X_c0 :  std_logic_vector(2 downto 0);
signal tile_26_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_26_output_c0 :  std_logic_vector(4 downto 0);
signal tile_26_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w26_2_c0 :  std_logic;
signal bh7_w27_3_c0 :  std_logic;
signal bh7_w28_4_c0 :  std_logic;
signal bh7_w29_6_c0 :  std_logic;
signal bh7_w30_6_c0 :  std_logic;
signal tile_27_X_c0 :  std_logic_vector(2 downto 0);
signal tile_27_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_27_output_c0 :  std_logic_vector(4 downto 0);
signal tile_27_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w23_1_c0 :  std_logic;
signal bh7_w24_1_c0 :  std_logic;
signal bh7_w25_2_c0 :  std_logic;
signal bh7_w26_3_c0 :  std_logic;
signal bh7_w27_4_c0 :  std_logic;
signal tile_28_X_c0 :  std_logic_vector(0 downto 0);
signal tile_28_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_28_output_c0 :  std_logic_vector(1 downto 0);
signal tile_28_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w27_5_c0 :  std_logic;
signal bh7_w28_5_c0 :  std_logic;
signal tile_29_X_c0 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_29_output_c0 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w24_2_c0 :  std_logic;
signal bh7_w25_3_c0 :  std_logic;
signal bh7_w26_4_c0 :  std_logic;
signal bh7_w27_6_c0 :  std_logic;
signal bh7_w28_6_c0 :  std_logic;
signal tile_30_X_c0 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_30_output_c0 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w21_1_c0 :  std_logic;
signal bh7_w22_1_c0 :  std_logic;
signal bh7_w23_2_c0 :  std_logic;
signal bh7_w24_3_c0 :  std_logic;
signal bh7_w25_4_c0 :  std_logic;
signal tile_31_X_c0 :  std_logic_vector(0 downto 0);
signal tile_31_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_31_output_c0 :  std_logic_vector(1 downto 0);
signal tile_31_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w25_5_c0 :  std_logic;
signal bh7_w26_5_c0 :  std_logic;
signal tile_32_X_c0 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_32_output_c0 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w22_2_c0 :  std_logic;
signal bh7_w23_3_c0 :  std_logic;
signal bh7_w24_4_c0 :  std_logic;
signal bh7_w25_6_c0 :  std_logic;
signal bh7_w26_6_c0 :  std_logic;
signal tile_33_X_c0 :  std_logic_vector(2 downto 0);
signal tile_33_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_33_output_c0 :  std_logic_vector(4 downto 0);
signal tile_33_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w19_1_c0 :  std_logic;
signal bh7_w20_1_c0 :  std_logic;
signal bh7_w21_2_c0 :  std_logic;
signal bh7_w22_3_c0 :  std_logic;
signal bh7_w23_4_c0 :  std_logic;
signal tile_34_X_c0 :  std_logic_vector(0 downto 0);
signal tile_34_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_34_output_c0 :  std_logic_vector(1 downto 0);
signal tile_34_filtered_output_c0 :  unsigned(1-0 downto 0);
signal bh7_w23_5_c0 :  std_logic;
signal bh7_w24_5_c0 :  std_logic;
signal tile_35_X_c0 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_35_output_c0 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w20_2_c0 :  std_logic;
signal bh7_w21_3_c0 :  std_logic;
signal bh7_w22_4_c0 :  std_logic;
signal bh7_w23_6_c0 :  std_logic;
signal bh7_w24_6_c0 :  std_logic;
signal tile_36_X_c0 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_36_output_c0 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w17_1_c0 :  std_logic;
signal bh7_w18_1_c0 :  std_logic;
signal bh7_w19_2_c0 :  std_logic;
signal bh7_w20_3_c0 :  std_logic;
signal bh7_w21_4_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid157_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid157_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid157_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w18_2_c0 :  std_logic;
signal bh7_w19_3_c0 :  std_logic;
signal bh7_w20_4_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid157_Out0_copy158_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid161_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid161_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w20_5_c0 :  std_logic;
signal bh7_w21_5_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid160_bh7_uid161_Out0_copy162_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid165_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid165_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid165_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w21_6_c0 :  std_logic;
signal bh7_w22_5_c0 :  std_logic;
signal bh7_w23_7_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid165_Out0_copy166_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid167_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid167_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w22_6_c0 :  std_logic;
signal bh7_w23_8_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid160_bh7_uid167_Out0_copy168_c0 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid171_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid171_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w23_9_c0 :  std_logic;
signal bh7_w24_7_c0 :  std_logic;
signal bh7_w25_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid171_Out0_copy172_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid173_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid173_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w24_8_c0 :  std_logic;
signal bh7_w25_8_c0 :  std_logic;
signal bh7_w26_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid173_Out0_copy174_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid175_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid175_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w25_9_c0 :  std_logic;
signal bh7_w26_8_c0 :  std_logic;
signal bh7_w27_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid175_Out0_copy176_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid177_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid177_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w26_9_c0 :  std_logic;
signal bh7_w27_8_c0 :  std_logic;
signal bh7_w28_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid177_Out0_copy178_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid179_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid179_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w27_9_c0 :  std_logic;
signal bh7_w28_8_c0 :  std_logic;
signal bh7_w29_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid179_Out0_copy180_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid181_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid181_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w28_9_c0 :  std_logic;
signal bh7_w29_8_c0 :  std_logic;
signal bh7_w30_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid181_Out0_copy182_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid183_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid183_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w29_9_c0 :  std_logic;
signal bh7_w30_8_c0 :  std_logic;
signal bh7_w31_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid183_Out0_copy184_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid185_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid185_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w30_9_c0 :  std_logic;
signal bh7_w31_8_c0 :  std_logic;
signal bh7_w32_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid185_Out0_copy186_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid187_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid187_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w31_9_c0 :  std_logic;
signal bh7_w32_8_c0 :  std_logic;
signal bh7_w33_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid187_Out0_copy188_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid189_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid189_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w32_9_c0 :  std_logic;
signal bh7_w33_8_c0 :  std_logic;
signal bh7_w34_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid189_Out0_copy190_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid191_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid191_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w33_9_c0 :  std_logic;
signal bh7_w34_8_c0 :  std_logic;
signal bh7_w35_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid191_Out0_copy192_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid193_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid193_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w34_9_c0 :  std_logic;
signal bh7_w35_8_c0 :  std_logic;
signal bh7_w36_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid193_Out0_copy194_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid195_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid195_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w35_9_c0 :  std_logic;
signal bh7_w36_8_c0 :  std_logic;
signal bh7_w37_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid195_Out0_copy196_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid197_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid197_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w36_9_c0 :  std_logic;
signal bh7_w37_8_c0 :  std_logic;
signal bh7_w38_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid197_Out0_copy198_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid199_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid199_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w37_9_c0 :  std_logic;
signal bh7_w38_8_c0 :  std_logic;
signal bh7_w39_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid199_Out0_copy200_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid201_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid201_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w38_9_c0 :  std_logic;
signal bh7_w39_8_c0 :  std_logic;
signal bh7_w40_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid201_Out0_copy202_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid203_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid203_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w39_9_c0 :  std_logic;
signal bh7_w40_8_c0 :  std_logic;
signal bh7_w41_5_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid203_Out0_copy204_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid205_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid170_bh7_uid205_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w40_9_c0 :  std_logic;
signal bh7_w41_6_c0 :  std_logic;
signal bh7_w42_5_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid170_bh7_uid205_Out0_copy206_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid207_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid207_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid207_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w41_7_c0 :  std_logic;
signal bh7_w42_6_c0 :  std_logic;
signal bh7_w43_4_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid207_Out0_copy208_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid209_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid209_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid209_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w42_7_c0 :  std_logic;
signal bh7_w43_5_c0 :  std_logic;
signal bh7_w44_3_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid209_Out0_copy210_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid211_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid211_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid211_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w43_6_c0 :  std_logic;
signal bh7_w44_4_c0 :  std_logic;
signal bh7_w45_2_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid211_Out0_copy212_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid213_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid213_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid213_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w45_3_c0 :  std_logic;
signal bh7_w46_2_c0 :  std_logic;
signal bh7_w47_0_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid213_Out0_copy214_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid215_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid215_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid215_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w20_6_c0 :  std_logic;
signal bh7_w21_7_c0 :  std_logic;
signal bh7_w22_7_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid215_Out0_copy216_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid217_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid217_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w22_8_c0 :  std_logic;
signal bh7_w23_10_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid160_bh7_uid217_Out0_copy218_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid219_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid219_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid219_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w23_11_c0 :  std_logic;
signal bh7_w24_9_c0 :  std_logic;
signal bh7_w25_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid219_Out0_copy220_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid221_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid221_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid221_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w25_11_c0 :  std_logic;
signal bh7_w26_10_c0 :  std_logic;
signal bh7_w27_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid221_Out0_copy222_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid223_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid223_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid223_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w27_11_c0 :  std_logic;
signal bh7_w28_10_c0 :  std_logic;
signal bh7_w29_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid223_Out0_copy224_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid225_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid225_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid225_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w29_11_c0 :  std_logic;
signal bh7_w30_10_c0 :  std_logic;
signal bh7_w31_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid225_Out0_copy226_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid227_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid227_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid227_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w31_11_c0 :  std_logic;
signal bh7_w32_10_c0 :  std_logic;
signal bh7_w33_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid227_Out0_copy228_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid229_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid229_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid229_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w33_11_c0 :  std_logic;
signal bh7_w34_10_c0 :  std_logic;
signal bh7_w35_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid229_Out0_copy230_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid231_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid231_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid231_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w35_11_c0 :  std_logic;
signal bh7_w36_10_c0 :  std_logic;
signal bh7_w37_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid231_Out0_copy232_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid233_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid233_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid233_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w37_11_c0 :  std_logic;
signal bh7_w38_10_c0 :  std_logic;
signal bh7_w39_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid233_Out0_copy234_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid235_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid235_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid235_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w39_11_c0 :  std_logic;
signal bh7_w40_10_c0 :  std_logic;
signal bh7_w41_8_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid235_Out0_copy236_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid237_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid237_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid237_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w41_9_c0 :  std_logic;
signal bh7_w42_8_c0 :  std_logic;
signal bh7_w43_7_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid237_Out0_copy238_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid239_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid239_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w42_9_c0 :  std_logic;
signal bh7_w43_8_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid160_bh7_uid239_Out0_copy240_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid241_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid241_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid241_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w43_9_c0 :  std_logic;
signal bh7_w44_5_c0 :  std_logic;
signal bh7_w45_4_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid241_Out0_copy242_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid243_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid243_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid243_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w45_5_c0 :  std_logic;
signal bh7_w46_3_c0 :  std_logic;
signal bh7_w47_1_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid243_Out0_copy244_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid245_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid245_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid245_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w22_9_c0 :  std_logic;
signal bh7_w23_12_c0 :  std_logic;
signal bh7_w24_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid245_Out0_copy246_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid247_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid247_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid247_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w25_12_c0 :  std_logic;
signal bh7_w26_11_c0 :  std_logic;
signal bh7_w27_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid247_Out0_copy248_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid249_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid249_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid249_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w27_13_c0 :  std_logic;
signal bh7_w28_11_c0 :  std_logic;
signal bh7_w29_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid249_Out0_copy250_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid251_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid251_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid251_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w29_13_c0 :  std_logic;
signal bh7_w30_11_c0 :  std_logic;
signal bh7_w31_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid251_Out0_copy252_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid253_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid253_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid253_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w31_13_c0 :  std_logic;
signal bh7_w32_11_c0 :  std_logic;
signal bh7_w33_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid253_Out0_copy254_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid255_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid255_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid255_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w33_13_c0 :  std_logic;
signal bh7_w34_11_c0 :  std_logic;
signal bh7_w35_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid255_Out0_copy256_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid257_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid257_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid257_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w35_13_c0 :  std_logic;
signal bh7_w36_11_c0 :  std_logic;
signal bh7_w37_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid257_Out0_copy258_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid259_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid259_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid259_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w37_13_c0 :  std_logic;
signal bh7_w38_11_c0 :  std_logic;
signal bh7_w39_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid259_Out0_copy260_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid261_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid261_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid261_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w39_13_c0 :  std_logic;
signal bh7_w40_11_c0 :  std_logic;
signal bh7_w41_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid261_Out0_copy262_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid263_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid263_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid263_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w41_11_c0 :  std_logic;
signal bh7_w42_10_c0 :  std_logic;
signal bh7_w43_10_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid263_Out0_copy264_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid265_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid265_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid265_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w43_11_c0 :  std_logic;
signal bh7_w44_6_c0 :  std_logic;
signal bh7_w45_6_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid265_Out0_copy266_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid267_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid267_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid267_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w45_7_c0 :  std_logic;
signal bh7_w46_4_c0 :  std_logic;
signal bh7_w47_2_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid267_Out0_copy268_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid269_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid269_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w47_3_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid160_bh7_uid269_Out0_copy270_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid271_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid271_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid271_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w24_11_c0 :  std_logic;
signal bh7_w25_13_c0 :  std_logic;
signal bh7_w26_12_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid271_Out0_copy272_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid273_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid273_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid273_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w27_14_c0 :  std_logic;
signal bh7_w28_12_c0, bh7_w28_12_c1 :  std_logic;
signal bh7_w29_14_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid273_Out0_copy274_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid275_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid275_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid275_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w29_15_c0 :  std_logic;
signal bh7_w30_12_c0 :  std_logic;
signal bh7_w31_14_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid275_Out0_copy276_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid277_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid277_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid277_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w31_15_c0 :  std_logic;
signal bh7_w32_12_c0 :  std_logic;
signal bh7_w33_14_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid277_Out0_copy278_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid279_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid279_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid279_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w33_15_c0 :  std_logic;
signal bh7_w34_12_c0 :  std_logic;
signal bh7_w35_14_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid279_Out0_copy280_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid281_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid281_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid281_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w35_15_c0 :  std_logic;
signal bh7_w36_12_c0 :  std_logic;
signal bh7_w37_14_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid281_Out0_copy282_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid283_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid283_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid283_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w37_15_c0 :  std_logic;
signal bh7_w38_12_c0 :  std_logic;
signal bh7_w39_14_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid283_Out0_copy284_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid285_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid285_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid285_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w39_15_c0 :  std_logic;
signal bh7_w40_12_c0 :  std_logic;
signal bh7_w41_12_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid285_Out0_copy286_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid287_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid287_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid287_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w41_13_c0 :  std_logic;
signal bh7_w42_11_c0 :  std_logic;
signal bh7_w43_12_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid287_Out0_copy288_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid289_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid289_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid289_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w43_13_c0 :  std_logic;
signal bh7_w44_7_c0 :  std_logic;
signal bh7_w45_8_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid289_Out0_copy290_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid291_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid291_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid291_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w45_9_c0 :  std_logic;
signal bh7_w46_5_c0 :  std_logic;
signal bh7_w47_4_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid291_Out0_copy292_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid293_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid293_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid293_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w47_5_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid293_Out0_copy294_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid295_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid295_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w26_13_c1 :  std_logic;
signal bh7_w27_15_c1 :  std_logic;
signal bh7_w28_13_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_copy296_c0, Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_copy296_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid297_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid297_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_16_c1 :  std_logic;
signal bh7_w30_13_c1 :  std_logic;
signal bh7_w31_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_copy298_c0, Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_copy298_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid299_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid299_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_17_c1 :  std_logic;
signal bh7_w32_13_c1 :  std_logic;
signal bh7_w33_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_copy300_c0, Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_copy300_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid301_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid301_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_17_c1 :  std_logic;
signal bh7_w34_13_c1 :  std_logic;
signal bh7_w35_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_copy302_c0, Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_copy302_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid303_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid303_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w35_17_c1 :  std_logic;
signal bh7_w36_13_c1 :  std_logic;
signal bh7_w37_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_copy304_c0, Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_copy304_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid305_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid305_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w37_17_c1 :  std_logic;
signal bh7_w38_13_c1 :  std_logic;
signal bh7_w39_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_copy306_c0, Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_copy306_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid307_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid307_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w39_17_c1 :  std_logic;
signal bh7_w40_13_c1 :  std_logic;
signal bh7_w41_14_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_copy308_c0, Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_copy308_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid309_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid309_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w41_15_c1 :  std_logic;
signal bh7_w42_12_c1 :  std_logic;
signal bh7_w43_14_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_copy310_c0, Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_copy310_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid311_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid311_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w43_15_c1 :  std_logic;
signal bh7_w44_8_c1 :  std_logic;
signal bh7_w45_10_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_copy312_c0, Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_copy312_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid313_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid313_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w45_11_c1 :  std_logic;
signal bh7_w46_6_c1 :  std_logic;
signal bh7_w47_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_copy314_c0, Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_copy314_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid315_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid315_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid315_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w47_7_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid315_Out0_copy316_c0, Compressor_14_3_Freq300_uid164_bh7_uid315_Out0_copy316_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid317_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid317_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w17_2_c1 :  std_logic;
signal bh7_w18_3_c1 :  std_logic;
signal bh7_w19_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_copy318_c0, Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_copy318_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid319_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid319_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w19_5_c1 :  std_logic;
signal bh7_w20_7_c1 :  std_logic;
signal bh7_w21_8_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_copy320_c0, Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_copy320_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid321_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid321_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_9_c1 :  std_logic;
signal bh7_w22_10_c1 :  std_logic;
signal bh7_w23_13_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_copy322_c0, Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_copy322_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid323_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid323_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w23_14_c1 :  std_logic;
signal bh7_w24_12_c1 :  std_logic;
signal bh7_w25_14_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_copy324_c0, Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_copy324_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid325_In0_c0, Compressor_23_3_Freq300_uid156_bh7_uid325_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid325_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid325_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w25_15_c1 :  std_logic;
signal bh7_w26_14_c1 :  std_logic;
signal bh7_w27_16_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid325_Out0_copy326_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid327_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid327_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w27_17_c1 :  std_logic;
signal bh7_w28_14_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid160_bh7_uid327_Out0_copy328_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid329_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid329_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid329_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w28_15_c1 :  std_logic;
signal bh7_w29_17_c1 :  std_logic;
signal bh7_w30_14_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid329_Out0_copy330_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid331_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid160_bh7_uid331_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w30_15_c1 :  std_logic;
signal bh7_w31_18_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid160_bh7_uid331_Out0_copy332_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid333_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid333_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid333_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_19_c1 :  std_logic;
signal bh7_w32_14_c1 :  std_logic;
signal bh7_w33_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid333_Out0_copy334_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid335_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid335_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid335_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_19_c1 :  std_logic;
signal bh7_w34_14_c1 :  std_logic;
signal bh7_w35_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid335_Out0_copy336_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid337_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid337_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid337_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w35_19_c1 :  std_logic;
signal bh7_w36_14_c1 :  std_logic;
signal bh7_w37_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid337_Out0_copy338_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid339_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid339_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid339_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w37_19_c1 :  std_logic;
signal bh7_w38_14_c1 :  std_logic;
signal bh7_w39_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid339_Out0_copy340_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid341_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid341_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid156_bh7_uid341_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w39_19_c1 :  std_logic;
signal bh7_w40_14_c1 :  std_logic;
signal bh7_w41_16_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid156_bh7_uid341_Out0_copy342_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid343_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid343_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid343_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w41_17_c1 :  std_logic;
signal bh7_w42_13_c1 :  std_logic;
signal bh7_w43_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid343_Out0_copy344_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid345_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid345_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid345_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w43_17_c1 :  std_logic;
signal bh7_w44_9_c1 :  std_logic;
signal bh7_w45_12_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid345_Out0_copy346_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid347_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid347_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid347_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w45_13_c1 :  std_logic;
signal bh7_w46_7_c1 :  std_logic;
signal bh7_w47_8_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid347_Out0_copy348_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid349_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid349_In1_c0, Compressor_14_3_Freq300_uid164_bh7_uid349_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid164_bh7_uid349_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w47_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid164_bh7_uid349_Out0_copy350_c1 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh7_18_c1 :  std_logic_vector(18 downto 0);
signal bitheapFinalAdd_bh7_In0_c1 :  std_logic_vector(29 downto 0);
signal bitheapFinalAdd_bh7_In1_c1 :  std_logic_vector(29 downto 0);
signal bitheapFinalAdd_bh7_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh7_Out_c1 :  std_logic_vector(29 downto 0);
signal bitheapResult_bh7_c1 :  std_logic_vector(47 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               bh7_w0_0_c1 <= bh7_w0_0_c0;
               bh7_w1_0_c1 <= bh7_w1_0_c0;
               bh7_w2_0_c1 <= bh7_w2_0_c0;
               bh7_w3_0_c1 <= bh7_w3_0_c0;
               bh7_w4_0_c1 <= bh7_w4_0_c0;
               bh7_w5_0_c1 <= bh7_w5_0_c0;
               bh7_w6_0_c1 <= bh7_w6_0_c0;
               bh7_w7_0_c1 <= bh7_w7_0_c0;
               bh7_w8_0_c1 <= bh7_w8_0_c0;
               bh7_w9_0_c1 <= bh7_w9_0_c0;
               bh7_w10_0_c1 <= bh7_w10_0_c0;
               bh7_w11_0_c1 <= bh7_w11_0_c0;
               bh7_w12_0_c1 <= bh7_w12_0_c0;
               bh7_w13_0_c1 <= bh7_w13_0_c0;
               bh7_w14_0_c1 <= bh7_w14_0_c0;
               bh7_w15_0_c1 <= bh7_w15_0_c0;
               bh7_w16_0_c1 <= bh7_w16_0_c0;
               bh7_w26_0_c1 <= bh7_w26_0_c0;
               bh7_w27_0_c1 <= bh7_w27_0_c0;
               bh7_w28_0_c1 <= bh7_w28_0_c0;
               bh7_w29_0_c1 <= bh7_w29_0_c0;
               bh7_w30_0_c1 <= bh7_w30_0_c0;
               bh7_w31_0_c1 <= bh7_w31_0_c0;
               bh7_w32_0_c1 <= bh7_w32_0_c0;
               bh7_w33_0_c1 <= bh7_w33_0_c0;
               bh7_w34_0_c1 <= bh7_w34_0_c0;
               bh7_w35_0_c1 <= bh7_w35_0_c0;
               bh7_w36_0_c1 <= bh7_w36_0_c0;
               bh7_w37_0_c1 <= bh7_w37_0_c0;
               bh7_w38_0_c1 <= bh7_w38_0_c0;
               bh7_w39_0_c1 <= bh7_w39_0_c0;
               bh7_w40_0_c1 <= bh7_w40_0_c0;
               bh7_w28_12_c1 <= bh7_w28_12_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_copy296_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_copy296_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_copy298_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_copy298_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_copy300_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_copy300_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_copy302_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_copy302_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_copy304_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_copy304_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_copy306_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_copy306_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_copy308_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_copy308_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_copy310_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_copy310_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_copy312_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_copy312_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_copy314_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_copy314_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid315_Out0_copy316_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid315_Out0_copy316_c0;
               Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_copy318_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_copy318_c0;
               Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_copy320_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_copy320_c0;
               Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_copy322_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_copy322_c0;
               Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_copy324_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_copy324_c0;
               Compressor_23_3_Freq300_uid156_bh7_uid325_In0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid325_In0_c0;
               Compressor_14_3_Freq300_uid164_bh7_uid349_In1_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid349_In1_c0;
            end if;
         end if;
      end process;
   XX_m6_c0 <= X ;
   YY_m6_c0 <= Y ;
   tile_0_X_c0 <= X(16 downto 0);
   tile_0_Y_c0 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid9
      port map ( clk  => clk,
                 X => tile_0_X_c0,
                 Y => tile_0_Y_c0,
                 R => tile_0_output_c0);

   tile_0_filtered_output_c0 <= unsigned(tile_0_output_c0(40 downto 0));
   bh7_w0_0_c0 <= tile_0_filtered_output_c0(0);
   bh7_w1_0_c0 <= tile_0_filtered_output_c0(1);
   bh7_w2_0_c0 <= tile_0_filtered_output_c0(2);
   bh7_w3_0_c0 <= tile_0_filtered_output_c0(3);
   bh7_w4_0_c0 <= tile_0_filtered_output_c0(4);
   bh7_w5_0_c0 <= tile_0_filtered_output_c0(5);
   bh7_w6_0_c0 <= tile_0_filtered_output_c0(6);
   bh7_w7_0_c0 <= tile_0_filtered_output_c0(7);
   bh7_w8_0_c0 <= tile_0_filtered_output_c0(8);
   bh7_w9_0_c0 <= tile_0_filtered_output_c0(9);
   bh7_w10_0_c0 <= tile_0_filtered_output_c0(10);
   bh7_w11_0_c0 <= tile_0_filtered_output_c0(11);
   bh7_w12_0_c0 <= tile_0_filtered_output_c0(12);
   bh7_w13_0_c0 <= tile_0_filtered_output_c0(13);
   bh7_w14_0_c0 <= tile_0_filtered_output_c0(14);
   bh7_w15_0_c0 <= tile_0_filtered_output_c0(15);
   bh7_w16_0_c0 <= tile_0_filtered_output_c0(16);
   bh7_w17_0_c0 <= tile_0_filtered_output_c0(17);
   bh7_w18_0_c0 <= tile_0_filtered_output_c0(18);
   bh7_w19_0_c0 <= tile_0_filtered_output_c0(19);
   bh7_w20_0_c0 <= tile_0_filtered_output_c0(20);
   bh7_w21_0_c0 <= tile_0_filtered_output_c0(21);
   bh7_w22_0_c0 <= tile_0_filtered_output_c0(22);
   bh7_w23_0_c0 <= tile_0_filtered_output_c0(23);
   bh7_w24_0_c0 <= tile_0_filtered_output_c0(24);
   bh7_w25_0_c0 <= tile_0_filtered_output_c0(25);
   bh7_w26_0_c0 <= tile_0_filtered_output_c0(26);
   bh7_w27_0_c0 <= tile_0_filtered_output_c0(27);
   bh7_w28_0_c0 <= tile_0_filtered_output_c0(28);
   bh7_w29_0_c0 <= tile_0_filtered_output_c0(29);
   bh7_w30_0_c0 <= tile_0_filtered_output_c0(30);
   bh7_w31_0_c0 <= tile_0_filtered_output_c0(31);
   bh7_w32_0_c0 <= tile_0_filtered_output_c0(32);
   bh7_w33_0_c0 <= tile_0_filtered_output_c0(33);
   bh7_w34_0_c0 <= tile_0_filtered_output_c0(34);
   bh7_w35_0_c0 <= tile_0_filtered_output_c0(35);
   bh7_w36_0_c0 <= tile_0_filtered_output_c0(36);
   bh7_w37_0_c0 <= tile_0_filtered_output_c0(37);
   bh7_w38_0_c0 <= tile_0_filtered_output_c0(38);
   bh7_w39_0_c0 <= tile_0_filtered_output_c0(39);
   bh7_w40_0_c0 <= tile_0_filtered_output_c0(40);
   tile_1_X_c0 <= X(23 downto 23);
   tile_1_Y_c0 <= Y(23 downto 22);
   tile_1_mult: IntMultiplierLUT_1x2_Freq300_uid11
      port map ( clk  => clk,
                 X => tile_1_X_c0,
                 Y => tile_1_Y_c0,
                 R => tile_1_output_c0);

   tile_1_filtered_output_c0 <= unsigned(tile_1_output_c0(1 downto 0));
   bh7_w45_0_c0 <= tile_1_filtered_output_c0(0);
   bh7_w46_0_c0 <= tile_1_filtered_output_c0(1);
   tile_2_X_c0 <= X(22 downto 20);
   tile_2_Y_c0 <= Y(23 downto 22);
   tile_2_mult: IntMultiplierLUT_3x2_Freq300_uid13
      port map ( clk  => clk,
                 X => tile_2_X_c0,
                 Y => tile_2_Y_c0,
                 R => tile_2_output_c0);

   tile_2_filtered_output_c0 <= unsigned(tile_2_output_c0(4 downto 0));
   bh7_w42_0_c0 <= tile_2_filtered_output_c0(0);
   bh7_w43_0_c0 <= tile_2_filtered_output_c0(1);
   bh7_w44_0_c0 <= tile_2_filtered_output_c0(2);
   bh7_w45_1_c0 <= tile_2_filtered_output_c0(3);
   bh7_w46_1_c0 <= tile_2_filtered_output_c0(4);
   tile_3_X_c0 <= X(19 downto 17);
   tile_3_Y_c0 <= Y(23 downto 22);
   tile_3_mult: IntMultiplierLUT_3x2_Freq300_uid18
      port map ( clk  => clk,
                 X => tile_3_X_c0,
                 Y => tile_3_Y_c0,
                 R => tile_3_output_c0);

   tile_3_filtered_output_c0 <= unsigned(tile_3_output_c0(4 downto 0));
   bh7_w39_1_c0 <= tile_3_filtered_output_c0(0);
   bh7_w40_1_c0 <= tile_3_filtered_output_c0(1);
   bh7_w41_0_c0 <= tile_3_filtered_output_c0(2);
   bh7_w42_1_c0 <= tile_3_filtered_output_c0(3);
   bh7_w43_1_c0 <= tile_3_filtered_output_c0(4);
   tile_4_X_c0 <= X(23 downto 23);
   tile_4_Y_c0 <= Y(21 downto 20);
   tile_4_mult: IntMultiplierLUT_1x2_Freq300_uid23
      port map ( clk  => clk,
                 X => tile_4_X_c0,
                 Y => tile_4_Y_c0,
                 R => tile_4_output_c0);

   tile_4_filtered_output_c0 <= unsigned(tile_4_output_c0(1 downto 0));
   bh7_w43_2_c0 <= tile_4_filtered_output_c0(0);
   bh7_w44_1_c0 <= tile_4_filtered_output_c0(1);
   tile_5_X_c0 <= X(22 downto 20);
   tile_5_Y_c0 <= Y(21 downto 20);
   tile_5_mult: IntMultiplierLUT_3x2_Freq300_uid25
      port map ( clk  => clk,
                 X => tile_5_X_c0,
                 Y => tile_5_Y_c0,
                 R => tile_5_output_c0);

   tile_5_filtered_output_c0 <= unsigned(tile_5_output_c0(4 downto 0));
   bh7_w40_2_c0 <= tile_5_filtered_output_c0(0);
   bh7_w41_1_c0 <= tile_5_filtered_output_c0(1);
   bh7_w42_2_c0 <= tile_5_filtered_output_c0(2);
   bh7_w43_3_c0 <= tile_5_filtered_output_c0(3);
   bh7_w44_2_c0 <= tile_5_filtered_output_c0(4);
   tile_6_X_c0 <= X(19 downto 17);
   tile_6_Y_c0 <= Y(21 downto 20);
   tile_6_mult: IntMultiplierLUT_3x2_Freq300_uid30
      port map ( clk  => clk,
                 X => tile_6_X_c0,
                 Y => tile_6_Y_c0,
                 R => tile_6_output_c0);

   tile_6_filtered_output_c0 <= unsigned(tile_6_output_c0(4 downto 0));
   bh7_w37_1_c0 <= tile_6_filtered_output_c0(0);
   bh7_w38_1_c0 <= tile_6_filtered_output_c0(1);
   bh7_w39_2_c0 <= tile_6_filtered_output_c0(2);
   bh7_w40_3_c0 <= tile_6_filtered_output_c0(3);
   bh7_w41_2_c0 <= tile_6_filtered_output_c0(4);
   tile_7_X_c0 <= X(23 downto 23);
   tile_7_Y_c0 <= Y(19 downto 18);
   tile_7_mult: IntMultiplierLUT_1x2_Freq300_uid35
      port map ( clk  => clk,
                 X => tile_7_X_c0,
                 Y => tile_7_Y_c0,
                 R => tile_7_output_c0);

   tile_7_filtered_output_c0 <= unsigned(tile_7_output_c0(1 downto 0));
   bh7_w41_3_c0 <= tile_7_filtered_output_c0(0);
   bh7_w42_3_c0 <= tile_7_filtered_output_c0(1);
   tile_8_X_c0 <= X(22 downto 20);
   tile_8_Y_c0 <= Y(19 downto 18);
   tile_8_mult: IntMultiplierLUT_3x2_Freq300_uid37
      port map ( clk  => clk,
                 X => tile_8_X_c0,
                 Y => tile_8_Y_c0,
                 R => tile_8_output_c0);

   tile_8_filtered_output_c0 <= unsigned(tile_8_output_c0(4 downto 0));
   bh7_w38_2_c0 <= tile_8_filtered_output_c0(0);
   bh7_w39_3_c0 <= tile_8_filtered_output_c0(1);
   bh7_w40_4_c0 <= tile_8_filtered_output_c0(2);
   bh7_w41_4_c0 <= tile_8_filtered_output_c0(3);
   bh7_w42_4_c0 <= tile_8_filtered_output_c0(4);
   tile_9_X_c0 <= X(19 downto 17);
   tile_9_Y_c0 <= Y(19 downto 18);
   tile_9_mult: IntMultiplierLUT_3x2_Freq300_uid42
      port map ( clk  => clk,
                 X => tile_9_X_c0,
                 Y => tile_9_Y_c0,
                 R => tile_9_output_c0);

   tile_9_filtered_output_c0 <= unsigned(tile_9_output_c0(4 downto 0));
   bh7_w35_1_c0 <= tile_9_filtered_output_c0(0);
   bh7_w36_1_c0 <= tile_9_filtered_output_c0(1);
   bh7_w37_2_c0 <= tile_9_filtered_output_c0(2);
   bh7_w38_3_c0 <= tile_9_filtered_output_c0(3);
   bh7_w39_4_c0 <= tile_9_filtered_output_c0(4);
   tile_10_X_c0 <= X(23 downto 23);
   tile_10_Y_c0 <= Y(17 downto 16);
   tile_10_mult: IntMultiplierLUT_1x2_Freq300_uid47
      port map ( clk  => clk,
                 X => tile_10_X_c0,
                 Y => tile_10_Y_c0,
                 R => tile_10_output_c0);

   tile_10_filtered_output_c0 <= unsigned(tile_10_output_c0(1 downto 0));
   bh7_w39_5_c0 <= tile_10_filtered_output_c0(0);
   bh7_w40_5_c0 <= tile_10_filtered_output_c0(1);
   tile_11_X_c0 <= X(22 downto 20);
   tile_11_Y_c0 <= Y(17 downto 16);
   tile_11_mult: IntMultiplierLUT_3x2_Freq300_uid49
      port map ( clk  => clk,
                 X => tile_11_X_c0,
                 Y => tile_11_Y_c0,
                 R => tile_11_output_c0);

   tile_11_filtered_output_c0 <= unsigned(tile_11_output_c0(4 downto 0));
   bh7_w36_2_c0 <= tile_11_filtered_output_c0(0);
   bh7_w37_3_c0 <= tile_11_filtered_output_c0(1);
   bh7_w38_4_c0 <= tile_11_filtered_output_c0(2);
   bh7_w39_6_c0 <= tile_11_filtered_output_c0(3);
   bh7_w40_6_c0 <= tile_11_filtered_output_c0(4);
   tile_12_X_c0 <= X(19 downto 17);
   tile_12_Y_c0 <= Y(17 downto 16);
   tile_12_mult: IntMultiplierLUT_3x2_Freq300_uid54
      port map ( clk  => clk,
                 X => tile_12_X_c0,
                 Y => tile_12_Y_c0,
                 R => tile_12_output_c0);

   tile_12_filtered_output_c0 <= unsigned(tile_12_output_c0(4 downto 0));
   bh7_w33_1_c0 <= tile_12_filtered_output_c0(0);
   bh7_w34_1_c0 <= tile_12_filtered_output_c0(1);
   bh7_w35_2_c0 <= tile_12_filtered_output_c0(2);
   bh7_w36_3_c0 <= tile_12_filtered_output_c0(3);
   bh7_w37_4_c0 <= tile_12_filtered_output_c0(4);
   tile_13_X_c0 <= X(23 downto 23);
   tile_13_Y_c0 <= Y(15 downto 14);
   tile_13_mult: IntMultiplierLUT_1x2_Freq300_uid59
      port map ( clk  => clk,
                 X => tile_13_X_c0,
                 Y => tile_13_Y_c0,
                 R => tile_13_output_c0);

   tile_13_filtered_output_c0 <= unsigned(tile_13_output_c0(1 downto 0));
   bh7_w37_5_c0 <= tile_13_filtered_output_c0(0);
   bh7_w38_5_c0 <= tile_13_filtered_output_c0(1);
   tile_14_X_c0 <= X(22 downto 20);
   tile_14_Y_c0 <= Y(15 downto 14);
   tile_14_mult: IntMultiplierLUT_3x2_Freq300_uid61
      port map ( clk  => clk,
                 X => tile_14_X_c0,
                 Y => tile_14_Y_c0,
                 R => tile_14_output_c0);

   tile_14_filtered_output_c0 <= unsigned(tile_14_output_c0(4 downto 0));
   bh7_w34_2_c0 <= tile_14_filtered_output_c0(0);
   bh7_w35_3_c0 <= tile_14_filtered_output_c0(1);
   bh7_w36_4_c0 <= tile_14_filtered_output_c0(2);
   bh7_w37_6_c0 <= tile_14_filtered_output_c0(3);
   bh7_w38_6_c0 <= tile_14_filtered_output_c0(4);
   tile_15_X_c0 <= X(19 downto 17);
   tile_15_Y_c0 <= Y(15 downto 14);
   tile_15_mult: IntMultiplierLUT_3x2_Freq300_uid66
      port map ( clk  => clk,
                 X => tile_15_X_c0,
                 Y => tile_15_Y_c0,
                 R => tile_15_output_c0);

   tile_15_filtered_output_c0 <= unsigned(tile_15_output_c0(4 downto 0));
   bh7_w31_1_c0 <= tile_15_filtered_output_c0(0);
   bh7_w32_1_c0 <= tile_15_filtered_output_c0(1);
   bh7_w33_2_c0 <= tile_15_filtered_output_c0(2);
   bh7_w34_3_c0 <= tile_15_filtered_output_c0(3);
   bh7_w35_4_c0 <= tile_15_filtered_output_c0(4);
   tile_16_X_c0 <= X(23 downto 23);
   tile_16_Y_c0 <= Y(13 downto 12);
   tile_16_mult: IntMultiplierLUT_1x2_Freq300_uid71
      port map ( clk  => clk,
                 X => tile_16_X_c0,
                 Y => tile_16_Y_c0,
                 R => tile_16_output_c0);

   tile_16_filtered_output_c0 <= unsigned(tile_16_output_c0(1 downto 0));
   bh7_w35_5_c0 <= tile_16_filtered_output_c0(0);
   bh7_w36_5_c0 <= tile_16_filtered_output_c0(1);
   tile_17_X_c0 <= X(22 downto 20);
   tile_17_Y_c0 <= Y(13 downto 12);
   tile_17_mult: IntMultiplierLUT_3x2_Freq300_uid73
      port map ( clk  => clk,
                 X => tile_17_X_c0,
                 Y => tile_17_Y_c0,
                 R => tile_17_output_c0);

   tile_17_filtered_output_c0 <= unsigned(tile_17_output_c0(4 downto 0));
   bh7_w32_2_c0 <= tile_17_filtered_output_c0(0);
   bh7_w33_3_c0 <= tile_17_filtered_output_c0(1);
   bh7_w34_4_c0 <= tile_17_filtered_output_c0(2);
   bh7_w35_6_c0 <= tile_17_filtered_output_c0(3);
   bh7_w36_6_c0 <= tile_17_filtered_output_c0(4);
   tile_18_X_c0 <= X(19 downto 17);
   tile_18_Y_c0 <= Y(13 downto 12);
   tile_18_mult: IntMultiplierLUT_3x2_Freq300_uid78
      port map ( clk  => clk,
                 X => tile_18_X_c0,
                 Y => tile_18_Y_c0,
                 R => tile_18_output_c0);

   tile_18_filtered_output_c0 <= unsigned(tile_18_output_c0(4 downto 0));
   bh7_w29_1_c0 <= tile_18_filtered_output_c0(0);
   bh7_w30_1_c0 <= tile_18_filtered_output_c0(1);
   bh7_w31_2_c0 <= tile_18_filtered_output_c0(2);
   bh7_w32_3_c0 <= tile_18_filtered_output_c0(3);
   bh7_w33_4_c0 <= tile_18_filtered_output_c0(4);
   tile_19_X_c0 <= X(23 downto 23);
   tile_19_Y_c0 <= Y(11 downto 10);
   tile_19_mult: IntMultiplierLUT_1x2_Freq300_uid83
      port map ( clk  => clk,
                 X => tile_19_X_c0,
                 Y => tile_19_Y_c0,
                 R => tile_19_output_c0);

   tile_19_filtered_output_c0 <= unsigned(tile_19_output_c0(1 downto 0));
   bh7_w33_5_c0 <= tile_19_filtered_output_c0(0);
   bh7_w34_5_c0 <= tile_19_filtered_output_c0(1);
   tile_20_X_c0 <= X(22 downto 20);
   tile_20_Y_c0 <= Y(11 downto 10);
   tile_20_mult: IntMultiplierLUT_3x2_Freq300_uid85
      port map ( clk  => clk,
                 X => tile_20_X_c0,
                 Y => tile_20_Y_c0,
                 R => tile_20_output_c0);

   tile_20_filtered_output_c0 <= unsigned(tile_20_output_c0(4 downto 0));
   bh7_w30_2_c0 <= tile_20_filtered_output_c0(0);
   bh7_w31_3_c0 <= tile_20_filtered_output_c0(1);
   bh7_w32_4_c0 <= tile_20_filtered_output_c0(2);
   bh7_w33_6_c0 <= tile_20_filtered_output_c0(3);
   bh7_w34_6_c0 <= tile_20_filtered_output_c0(4);
   tile_21_X_c0 <= X(19 downto 17);
   tile_21_Y_c0 <= Y(11 downto 10);
   tile_21_mult: IntMultiplierLUT_3x2_Freq300_uid90
      port map ( clk  => clk,
                 X => tile_21_X_c0,
                 Y => tile_21_Y_c0,
                 R => tile_21_output_c0);

   tile_21_filtered_output_c0 <= unsigned(tile_21_output_c0(4 downto 0));
   bh7_w27_1_c0 <= tile_21_filtered_output_c0(0);
   bh7_w28_1_c0 <= tile_21_filtered_output_c0(1);
   bh7_w29_2_c0 <= tile_21_filtered_output_c0(2);
   bh7_w30_3_c0 <= tile_21_filtered_output_c0(3);
   bh7_w31_4_c0 <= tile_21_filtered_output_c0(4);
   tile_22_X_c0 <= X(23 downto 23);
   tile_22_Y_c0 <= Y(9 downto 8);
   tile_22_mult: IntMultiplierLUT_1x2_Freq300_uid95
      port map ( clk  => clk,
                 X => tile_22_X_c0,
                 Y => tile_22_Y_c0,
                 R => tile_22_output_c0);

   tile_22_filtered_output_c0 <= unsigned(tile_22_output_c0(1 downto 0));
   bh7_w31_5_c0 <= tile_22_filtered_output_c0(0);
   bh7_w32_5_c0 <= tile_22_filtered_output_c0(1);
   tile_23_X_c0 <= X(22 downto 20);
   tile_23_Y_c0 <= Y(9 downto 8);
   tile_23_mult: IntMultiplierLUT_3x2_Freq300_uid97
      port map ( clk  => clk,
                 X => tile_23_X_c0,
                 Y => tile_23_Y_c0,
                 R => tile_23_output_c0);

   tile_23_filtered_output_c0 <= unsigned(tile_23_output_c0(4 downto 0));
   bh7_w28_2_c0 <= tile_23_filtered_output_c0(0);
   bh7_w29_3_c0 <= tile_23_filtered_output_c0(1);
   bh7_w30_4_c0 <= tile_23_filtered_output_c0(2);
   bh7_w31_6_c0 <= tile_23_filtered_output_c0(3);
   bh7_w32_6_c0 <= tile_23_filtered_output_c0(4);
   tile_24_X_c0 <= X(19 downto 17);
   tile_24_Y_c0 <= Y(9 downto 8);
   tile_24_mult: IntMultiplierLUT_3x2_Freq300_uid102
      port map ( clk  => clk,
                 X => tile_24_X_c0,
                 Y => tile_24_Y_c0,
                 R => tile_24_output_c0);

   tile_24_filtered_output_c0 <= unsigned(tile_24_output_c0(4 downto 0));
   bh7_w25_1_c0 <= tile_24_filtered_output_c0(0);
   bh7_w26_1_c0 <= tile_24_filtered_output_c0(1);
   bh7_w27_2_c0 <= tile_24_filtered_output_c0(2);
   bh7_w28_3_c0 <= tile_24_filtered_output_c0(3);
   bh7_w29_4_c0 <= tile_24_filtered_output_c0(4);
   tile_25_X_c0 <= X(23 downto 23);
   tile_25_Y_c0 <= Y(7 downto 6);
   tile_25_mult: IntMultiplierLUT_1x2_Freq300_uid107
      port map ( clk  => clk,
                 X => tile_25_X_c0,
                 Y => tile_25_Y_c0,
                 R => tile_25_output_c0);

   tile_25_filtered_output_c0 <= unsigned(tile_25_output_c0(1 downto 0));
   bh7_w29_5_c0 <= tile_25_filtered_output_c0(0);
   bh7_w30_5_c0 <= tile_25_filtered_output_c0(1);
   tile_26_X_c0 <= X(22 downto 20);
   tile_26_Y_c0 <= Y(7 downto 6);
   tile_26_mult: IntMultiplierLUT_3x2_Freq300_uid109
      port map ( clk  => clk,
                 X => tile_26_X_c0,
                 Y => tile_26_Y_c0,
                 R => tile_26_output_c0);

   tile_26_filtered_output_c0 <= unsigned(tile_26_output_c0(4 downto 0));
   bh7_w26_2_c0 <= tile_26_filtered_output_c0(0);
   bh7_w27_3_c0 <= tile_26_filtered_output_c0(1);
   bh7_w28_4_c0 <= tile_26_filtered_output_c0(2);
   bh7_w29_6_c0 <= tile_26_filtered_output_c0(3);
   bh7_w30_6_c0 <= tile_26_filtered_output_c0(4);
   tile_27_X_c0 <= X(19 downto 17);
   tile_27_Y_c0 <= Y(7 downto 6);
   tile_27_mult: IntMultiplierLUT_3x2_Freq300_uid114
      port map ( clk  => clk,
                 X => tile_27_X_c0,
                 Y => tile_27_Y_c0,
                 R => tile_27_output_c0);

   tile_27_filtered_output_c0 <= unsigned(tile_27_output_c0(4 downto 0));
   bh7_w23_1_c0 <= tile_27_filtered_output_c0(0);
   bh7_w24_1_c0 <= tile_27_filtered_output_c0(1);
   bh7_w25_2_c0 <= tile_27_filtered_output_c0(2);
   bh7_w26_3_c0 <= tile_27_filtered_output_c0(3);
   bh7_w27_4_c0 <= tile_27_filtered_output_c0(4);
   tile_28_X_c0 <= X(23 downto 23);
   tile_28_Y_c0 <= Y(5 downto 4);
   tile_28_mult: IntMultiplierLUT_1x2_Freq300_uid119
      port map ( clk  => clk,
                 X => tile_28_X_c0,
                 Y => tile_28_Y_c0,
                 R => tile_28_output_c0);

   tile_28_filtered_output_c0 <= unsigned(tile_28_output_c0(1 downto 0));
   bh7_w27_5_c0 <= tile_28_filtered_output_c0(0);
   bh7_w28_5_c0 <= tile_28_filtered_output_c0(1);
   tile_29_X_c0 <= X(22 downto 20);
   tile_29_Y_c0 <= Y(5 downto 4);
   tile_29_mult: IntMultiplierLUT_3x2_Freq300_uid121
      port map ( clk  => clk,
                 X => tile_29_X_c0,
                 Y => tile_29_Y_c0,
                 R => tile_29_output_c0);

   tile_29_filtered_output_c0 <= unsigned(tile_29_output_c0(4 downto 0));
   bh7_w24_2_c0 <= tile_29_filtered_output_c0(0);
   bh7_w25_3_c0 <= tile_29_filtered_output_c0(1);
   bh7_w26_4_c0 <= tile_29_filtered_output_c0(2);
   bh7_w27_6_c0 <= tile_29_filtered_output_c0(3);
   bh7_w28_6_c0 <= tile_29_filtered_output_c0(4);
   tile_30_X_c0 <= X(19 downto 17);
   tile_30_Y_c0 <= Y(5 downto 4);
   tile_30_mult: IntMultiplierLUT_3x2_Freq300_uid126
      port map ( clk  => clk,
                 X => tile_30_X_c0,
                 Y => tile_30_Y_c0,
                 R => tile_30_output_c0);

   tile_30_filtered_output_c0 <= unsigned(tile_30_output_c0(4 downto 0));
   bh7_w21_1_c0 <= tile_30_filtered_output_c0(0);
   bh7_w22_1_c0 <= tile_30_filtered_output_c0(1);
   bh7_w23_2_c0 <= tile_30_filtered_output_c0(2);
   bh7_w24_3_c0 <= tile_30_filtered_output_c0(3);
   bh7_w25_4_c0 <= tile_30_filtered_output_c0(4);
   tile_31_X_c0 <= X(23 downto 23);
   tile_31_Y_c0 <= Y(3 downto 2);
   tile_31_mult: IntMultiplierLUT_1x2_Freq300_uid131
      port map ( clk  => clk,
                 X => tile_31_X_c0,
                 Y => tile_31_Y_c0,
                 R => tile_31_output_c0);

   tile_31_filtered_output_c0 <= unsigned(tile_31_output_c0(1 downto 0));
   bh7_w25_5_c0 <= tile_31_filtered_output_c0(0);
   bh7_w26_5_c0 <= tile_31_filtered_output_c0(1);
   tile_32_X_c0 <= X(22 downto 20);
   tile_32_Y_c0 <= Y(3 downto 2);
   tile_32_mult: IntMultiplierLUT_3x2_Freq300_uid133
      port map ( clk  => clk,
                 X => tile_32_X_c0,
                 Y => tile_32_Y_c0,
                 R => tile_32_output_c0);

   tile_32_filtered_output_c0 <= unsigned(tile_32_output_c0(4 downto 0));
   bh7_w22_2_c0 <= tile_32_filtered_output_c0(0);
   bh7_w23_3_c0 <= tile_32_filtered_output_c0(1);
   bh7_w24_4_c0 <= tile_32_filtered_output_c0(2);
   bh7_w25_6_c0 <= tile_32_filtered_output_c0(3);
   bh7_w26_6_c0 <= tile_32_filtered_output_c0(4);
   tile_33_X_c0 <= X(19 downto 17);
   tile_33_Y_c0 <= Y(3 downto 2);
   tile_33_mult: IntMultiplierLUT_3x2_Freq300_uid138
      port map ( clk  => clk,
                 X => tile_33_X_c0,
                 Y => tile_33_Y_c0,
                 R => tile_33_output_c0);

   tile_33_filtered_output_c0 <= unsigned(tile_33_output_c0(4 downto 0));
   bh7_w19_1_c0 <= tile_33_filtered_output_c0(0);
   bh7_w20_1_c0 <= tile_33_filtered_output_c0(1);
   bh7_w21_2_c0 <= tile_33_filtered_output_c0(2);
   bh7_w22_3_c0 <= tile_33_filtered_output_c0(3);
   bh7_w23_4_c0 <= tile_33_filtered_output_c0(4);
   tile_34_X_c0 <= X(23 downto 23);
   tile_34_Y_c0 <= Y(1 downto 0);
   tile_34_mult: IntMultiplierLUT_1x2_Freq300_uid143
      port map ( clk  => clk,
                 X => tile_34_X_c0,
                 Y => tile_34_Y_c0,
                 R => tile_34_output_c0);

   tile_34_filtered_output_c0 <= unsigned(tile_34_output_c0(1 downto 0));
   bh7_w23_5_c0 <= tile_34_filtered_output_c0(0);
   bh7_w24_5_c0 <= tile_34_filtered_output_c0(1);
   tile_35_X_c0 <= X(22 downto 20);
   tile_35_Y_c0 <= Y(1 downto 0);
   tile_35_mult: IntMultiplierLUT_3x2_Freq300_uid145
      port map ( clk  => clk,
                 X => tile_35_X_c0,
                 Y => tile_35_Y_c0,
                 R => tile_35_output_c0);

   tile_35_filtered_output_c0 <= unsigned(tile_35_output_c0(4 downto 0));
   bh7_w20_2_c0 <= tile_35_filtered_output_c0(0);
   bh7_w21_3_c0 <= tile_35_filtered_output_c0(1);
   bh7_w22_4_c0 <= tile_35_filtered_output_c0(2);
   bh7_w23_6_c0 <= tile_35_filtered_output_c0(3);
   bh7_w24_6_c0 <= tile_35_filtered_output_c0(4);
   tile_36_X_c0 <= X(19 downto 17);
   tile_36_Y_c0 <= Y(1 downto 0);
   tile_36_mult: IntMultiplierLUT_3x2_Freq300_uid150
      port map ( clk  => clk,
                 X => tile_36_X_c0,
                 Y => tile_36_Y_c0,
                 R => tile_36_output_c0);

   tile_36_filtered_output_c0 <= unsigned(tile_36_output_c0(4 downto 0));
   bh7_w17_1_c0 <= tile_36_filtered_output_c0(0);
   bh7_w18_1_c0 <= tile_36_filtered_output_c0(1);
   bh7_w19_2_c0 <= tile_36_filtered_output_c0(2);
   bh7_w20_3_c0 <= tile_36_filtered_output_c0(3);
   bh7_w21_4_c0 <= tile_36_filtered_output_c0(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq300_uid156_bh7_uid157_In0_c0 <= "" & bh7_w18_1_c0 & "0" & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid157_In1_c0 <= "" & bh7_w19_1_c0 & bh7_w19_2_c0;
   bh7_w18_2_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid157_Out0_c0(0);
   bh7_w19_3_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid157_Out0_c0(1);
   bh7_w20_4_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid157_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid157: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid157_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid157_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid157_Out0_copy158_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid157_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid157_Out0_copy158_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid160_bh7_uid161_In0_c0 <= "" & bh7_w20_1_c0 & bh7_w20_2_c0 & bh7_w20_3_c0;
   bh7_w20_5_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid161_Out0_c0(0);
   bh7_w21_5_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid161_Out0_c0(1);
   Compressor_3_2_Freq300_uid160_uid161: Compressor_3_2_Freq300_uid160
      port map ( X0 => Compressor_3_2_Freq300_uid160_bh7_uid161_In0_c0,
                 R => Compressor_3_2_Freq300_uid160_bh7_uid161_Out0_copy162_c0);
   Compressor_3_2_Freq300_uid160_bh7_uid161_Out0_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid161_Out0_copy162_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid165_In0_c0 <= "" & bh7_w21_1_c0 & bh7_w21_2_c0 & bh7_w21_3_c0 & bh7_w21_4_c0;
   Compressor_14_3_Freq300_uid164_bh7_uid165_In1_c0 <= "" & bh7_w22_1_c0;
   bh7_w21_6_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid165_Out0_c0(0);
   bh7_w22_5_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid165_Out0_c0(1);
   bh7_w23_7_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid165_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid165: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid165_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid165_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid165_Out0_copy166_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid165_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid165_Out0_copy166_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid160_bh7_uid167_In0_c0 <= "" & bh7_w22_2_c0 & bh7_w22_3_c0 & bh7_w22_4_c0;
   bh7_w22_6_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid167_Out0_c0(0);
   bh7_w23_8_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid167_Out0_c0(1);
   Compressor_3_2_Freq300_uid160_uid167: Compressor_3_2_Freq300_uid160
      port map ( X0 => Compressor_3_2_Freq300_uid160_bh7_uid167_In0_c0,
                 R => Compressor_3_2_Freq300_uid160_bh7_uid167_Out0_copy168_c0);
   Compressor_3_2_Freq300_uid160_bh7_uid167_Out0_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid167_Out0_copy168_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid171_In0_c0 <= "" & bh7_w23_1_c0 & bh7_w23_2_c0 & bh7_w23_3_c0 & bh7_w23_4_c0 & bh7_w23_5_c0 & bh7_w23_6_c0;
   bh7_w23_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid171_Out0_c0(0);
   bh7_w24_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid171_Out0_c0(1);
   bh7_w25_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid171_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid171: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid171_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid171_Out0_copy172_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid171_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid171_Out0_copy172_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid173_In0_c0 <= "" & bh7_w24_1_c0 & bh7_w24_2_c0 & bh7_w24_3_c0 & bh7_w24_4_c0 & bh7_w24_5_c0 & bh7_w24_6_c0;
   bh7_w24_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid173_Out0_c0(0);
   bh7_w25_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid173_Out0_c0(1);
   bh7_w26_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid173_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid173: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid173_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid173_Out0_copy174_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid173_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid173_Out0_copy174_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid175_In0_c0 <= "" & bh7_w25_1_c0 & bh7_w25_2_c0 & bh7_w25_3_c0 & bh7_w25_4_c0 & bh7_w25_5_c0 & bh7_w25_6_c0;
   bh7_w25_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid175_Out0_c0(0);
   bh7_w26_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid175_Out0_c0(1);
   bh7_w27_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid175_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid175: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid175_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid175_Out0_copy176_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid175_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid175_Out0_copy176_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid177_In0_c0 <= "" & bh7_w26_1_c0 & bh7_w26_2_c0 & bh7_w26_3_c0 & bh7_w26_4_c0 & bh7_w26_5_c0 & bh7_w26_6_c0;
   bh7_w26_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid177_Out0_c0(0);
   bh7_w27_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid177_Out0_c0(1);
   bh7_w28_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid177_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid177: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid177_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid177_Out0_copy178_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid177_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid177_Out0_copy178_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid179_In0_c0 <= "" & bh7_w27_1_c0 & bh7_w27_2_c0 & bh7_w27_3_c0 & bh7_w27_4_c0 & bh7_w27_5_c0 & bh7_w27_6_c0;
   bh7_w27_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid179_Out0_c0(0);
   bh7_w28_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid179_Out0_c0(1);
   bh7_w29_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid179_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid179: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid179_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid179_Out0_copy180_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid179_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid179_Out0_copy180_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid181_In0_c0 <= "" & bh7_w28_1_c0 & bh7_w28_2_c0 & bh7_w28_3_c0 & bh7_w28_4_c0 & bh7_w28_5_c0 & bh7_w28_6_c0;
   bh7_w28_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid181_Out0_c0(0);
   bh7_w29_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid181_Out0_c0(1);
   bh7_w30_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid181_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid181: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid181_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid181_Out0_copy182_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid181_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid181_Out0_copy182_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid183_In0_c0 <= "" & bh7_w29_1_c0 & bh7_w29_2_c0 & bh7_w29_3_c0 & bh7_w29_4_c0 & bh7_w29_5_c0 & bh7_w29_6_c0;
   bh7_w29_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid183_Out0_c0(0);
   bh7_w30_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid183_Out0_c0(1);
   bh7_w31_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid183_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid183: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid183_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid183_Out0_copy184_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid183_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid183_Out0_copy184_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid185_In0_c0 <= "" & bh7_w30_1_c0 & bh7_w30_2_c0 & bh7_w30_3_c0 & bh7_w30_4_c0 & bh7_w30_5_c0 & bh7_w30_6_c0;
   bh7_w30_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid185_Out0_c0(0);
   bh7_w31_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid185_Out0_c0(1);
   bh7_w32_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid185_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid185: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid185_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid185_Out0_copy186_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid185_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid185_Out0_copy186_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid187_In0_c0 <= "" & bh7_w31_1_c0 & bh7_w31_2_c0 & bh7_w31_3_c0 & bh7_w31_4_c0 & bh7_w31_5_c0 & bh7_w31_6_c0;
   bh7_w31_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid187_Out0_c0(0);
   bh7_w32_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid187_Out0_c0(1);
   bh7_w33_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid187_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid187: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid187_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid187_Out0_copy188_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid187_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid187_Out0_copy188_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid189_In0_c0 <= "" & bh7_w32_1_c0 & bh7_w32_2_c0 & bh7_w32_3_c0 & bh7_w32_4_c0 & bh7_w32_5_c0 & bh7_w32_6_c0;
   bh7_w32_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid189_Out0_c0(0);
   bh7_w33_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid189_Out0_c0(1);
   bh7_w34_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid189_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid189: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid189_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid189_Out0_copy190_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid189_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid189_Out0_copy190_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid191_In0_c0 <= "" & bh7_w33_1_c0 & bh7_w33_2_c0 & bh7_w33_3_c0 & bh7_w33_4_c0 & bh7_w33_5_c0 & bh7_w33_6_c0;
   bh7_w33_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid191_Out0_c0(0);
   bh7_w34_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid191_Out0_c0(1);
   bh7_w35_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid191_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid191: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid191_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid191_Out0_copy192_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid191_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid191_Out0_copy192_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid193_In0_c0 <= "" & bh7_w34_1_c0 & bh7_w34_2_c0 & bh7_w34_3_c0 & bh7_w34_4_c0 & bh7_w34_5_c0 & bh7_w34_6_c0;
   bh7_w34_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid193_Out0_c0(0);
   bh7_w35_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid193_Out0_c0(1);
   bh7_w36_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid193_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid193: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid193_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid193_Out0_copy194_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid193_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid193_Out0_copy194_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid195_In0_c0 <= "" & bh7_w35_1_c0 & bh7_w35_2_c0 & bh7_w35_3_c0 & bh7_w35_4_c0 & bh7_w35_5_c0 & bh7_w35_6_c0;
   bh7_w35_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid195_Out0_c0(0);
   bh7_w36_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid195_Out0_c0(1);
   bh7_w37_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid195_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid195: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid195_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid195_Out0_copy196_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid195_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid195_Out0_copy196_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid197_In0_c0 <= "" & bh7_w36_1_c0 & bh7_w36_2_c0 & bh7_w36_3_c0 & bh7_w36_4_c0 & bh7_w36_5_c0 & bh7_w36_6_c0;
   bh7_w36_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid197_Out0_c0(0);
   bh7_w37_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid197_Out0_c0(1);
   bh7_w38_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid197_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid197: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid197_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid197_Out0_copy198_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid197_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid197_Out0_copy198_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid199_In0_c0 <= "" & bh7_w37_1_c0 & bh7_w37_2_c0 & bh7_w37_3_c0 & bh7_w37_4_c0 & bh7_w37_5_c0 & bh7_w37_6_c0;
   bh7_w37_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid199_Out0_c0(0);
   bh7_w38_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid199_Out0_c0(1);
   bh7_w39_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid199_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid199: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid199_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid199_Out0_copy200_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid199_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid199_Out0_copy200_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid201_In0_c0 <= "" & bh7_w38_1_c0 & bh7_w38_2_c0 & bh7_w38_3_c0 & bh7_w38_4_c0 & bh7_w38_5_c0 & bh7_w38_6_c0;
   bh7_w38_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid201_Out0_c0(0);
   bh7_w39_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid201_Out0_c0(1);
   bh7_w40_7_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid201_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid201: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid201_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid201_Out0_copy202_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid201_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid201_Out0_copy202_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid203_In0_c0 <= "" & bh7_w39_1_c0 & bh7_w39_2_c0 & bh7_w39_3_c0 & bh7_w39_4_c0 & bh7_w39_5_c0 & bh7_w39_6_c0;
   bh7_w39_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid203_Out0_c0(0);
   bh7_w40_8_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid203_Out0_c0(1);
   bh7_w41_5_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid203_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid203: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid203_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid203_Out0_copy204_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid203_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid203_Out0_copy204_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid170_bh7_uid205_In0_c0 <= "" & bh7_w40_1_c0 & bh7_w40_2_c0 & bh7_w40_3_c0 & bh7_w40_4_c0 & bh7_w40_5_c0 & bh7_w40_6_c0;
   bh7_w40_9_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid205_Out0_c0(0);
   bh7_w41_6_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid205_Out0_c0(1);
   bh7_w42_5_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid205_Out0_c0(2);
   Compressor_6_3_Freq300_uid170_uid205: Compressor_6_3_Freq300_uid170
      port map ( X0 => Compressor_6_3_Freq300_uid170_bh7_uid205_In0_c0,
                 R => Compressor_6_3_Freq300_uid170_bh7_uid205_Out0_copy206_c0);
   Compressor_6_3_Freq300_uid170_bh7_uid205_Out0_c0 <= Compressor_6_3_Freq300_uid170_bh7_uid205_Out0_copy206_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid207_In0_c0 <= "" & bh7_w41_0_c0 & bh7_w41_1_c0 & bh7_w41_2_c0 & bh7_w41_3_c0;
   Compressor_14_3_Freq300_uid164_bh7_uid207_In1_c0 <= "" & bh7_w42_0_c0;
   bh7_w41_7_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid207_Out0_c0(0);
   bh7_w42_6_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid207_Out0_c0(1);
   bh7_w43_4_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid207_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid207: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid207_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid207_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid207_Out0_copy208_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid207_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid207_Out0_copy208_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid209_In0_c0 <= "" & bh7_w42_1_c0 & bh7_w42_2_c0 & bh7_w42_3_c0 & bh7_w42_4_c0;
   Compressor_14_3_Freq300_uid164_bh7_uid209_In1_c0 <= "" & bh7_w43_0_c0;
   bh7_w42_7_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid209_Out0_c0(0);
   bh7_w43_5_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid209_Out0_c0(1);
   bh7_w44_3_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid209_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid209: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid209_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid209_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid209_Out0_copy210_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid209_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid209_Out0_copy210_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid211_In0_c0 <= "" & bh7_w43_1_c0 & bh7_w43_2_c0 & bh7_w43_3_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid211_In1_c0 <= "" & bh7_w44_0_c0 & bh7_w44_1_c0;
   bh7_w43_6_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid211_Out0_c0(0);
   bh7_w44_4_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid211_Out0_c0(1);
   bh7_w45_2_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid211_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid211: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid211_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid211_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid211_Out0_copy212_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid211_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid211_Out0_copy212_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid213_In0_c0 <= "" & bh7_w45_0_c0 & bh7_w45_1_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid213_In1_c0 <= "" & bh7_w46_0_c0 & bh7_w46_1_c0;
   bh7_w45_3_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid213_Out0_c0(0);
   bh7_w46_2_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid213_Out0_c0(1);
   bh7_w47_0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid213_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid213: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid213_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid213_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid213_Out0_copy214_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid213_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid213_Out0_copy214_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid215_In0_c0 <= "" & bh7_w20_5_c0 & bh7_w20_4_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid215_In1_c0 <= "" & bh7_w21_6_c0 & bh7_w21_5_c0;
   bh7_w20_6_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid215_Out0_c0(0);
   bh7_w21_7_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid215_Out0_c0(1);
   bh7_w22_7_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid215_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid215: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid215_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid215_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid215_Out0_copy216_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid215_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid215_Out0_copy216_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid160_bh7_uid217_In0_c0 <= "" & bh7_w22_6_c0 & bh7_w22_5_c0 & "0";
   bh7_w22_8_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid217_Out0_c0(0);
   bh7_w23_10_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid217_Out0_c0(1);
   Compressor_3_2_Freq300_uid160_uid217: Compressor_3_2_Freq300_uid160
      port map ( X0 => Compressor_3_2_Freq300_uid160_bh7_uid217_In0_c0,
                 R => Compressor_3_2_Freq300_uid160_bh7_uid217_Out0_copy218_c0);
   Compressor_3_2_Freq300_uid160_bh7_uid217_Out0_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid217_Out0_copy218_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid219_In0_c0 <= "" & bh7_w23_8_c0 & bh7_w23_7_c0 & bh7_w23_9_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid219_In1_c0 <= "" & bh7_w24_8_c0 & bh7_w24_7_c0;
   bh7_w23_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid219_Out0_c0(0);
   bh7_w24_9_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid219_Out0_c0(1);
   bh7_w25_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid219_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid219: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid219_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid219_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid219_Out0_copy220_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid219_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid219_Out0_copy220_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid221_In0_c0 <= "" & bh7_w25_9_c0 & bh7_w25_8_c0 & bh7_w25_7_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid221_In1_c0 <= "" & bh7_w26_9_c0 & bh7_w26_8_c0;
   bh7_w25_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid221_Out0_c0(0);
   bh7_w26_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid221_Out0_c0(1);
   bh7_w27_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid221_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid221: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid221_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid221_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid221_Out0_copy222_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid221_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid221_Out0_copy222_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid223_In0_c0 <= "" & bh7_w27_9_c0 & bh7_w27_8_c0 & bh7_w27_7_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid223_In1_c0 <= "" & bh7_w28_9_c0 & bh7_w28_8_c0;
   bh7_w27_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid223_Out0_c0(0);
   bh7_w28_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid223_Out0_c0(1);
   bh7_w29_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid223_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid223: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid223_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid223_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid223_Out0_copy224_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid223_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid223_Out0_copy224_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid225_In0_c0 <= "" & bh7_w29_9_c0 & bh7_w29_8_c0 & bh7_w29_7_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid225_In1_c0 <= "" & bh7_w30_9_c0 & bh7_w30_8_c0;
   bh7_w29_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid225_Out0_c0(0);
   bh7_w30_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid225_Out0_c0(1);
   bh7_w31_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid225_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid225: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid225_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid225_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid225_Out0_copy226_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid225_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid225_Out0_copy226_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid227_In0_c0 <= "" & bh7_w31_9_c0 & bh7_w31_8_c0 & bh7_w31_7_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid227_In1_c0 <= "" & bh7_w32_9_c0 & bh7_w32_8_c0;
   bh7_w31_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid227_Out0_c0(0);
   bh7_w32_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid227_Out0_c0(1);
   bh7_w33_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid227_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid227: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid227_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid227_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid227_Out0_copy228_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid227_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid227_Out0_copy228_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid229_In0_c0 <= "" & bh7_w33_9_c0 & bh7_w33_8_c0 & bh7_w33_7_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid229_In1_c0 <= "" & bh7_w34_9_c0 & bh7_w34_8_c0;
   bh7_w33_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid229_Out0_c0(0);
   bh7_w34_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid229_Out0_c0(1);
   bh7_w35_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid229_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid229: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid229_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid229_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid229_Out0_copy230_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid229_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid229_Out0_copy230_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid231_In0_c0 <= "" & bh7_w35_9_c0 & bh7_w35_8_c0 & bh7_w35_7_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid231_In1_c0 <= "" & bh7_w36_9_c0 & bh7_w36_8_c0;
   bh7_w35_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid231_Out0_c0(0);
   bh7_w36_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid231_Out0_c0(1);
   bh7_w37_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid231_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid231: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid231_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid231_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid231_Out0_copy232_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid231_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid231_Out0_copy232_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid233_In0_c0 <= "" & bh7_w37_9_c0 & bh7_w37_8_c0 & bh7_w37_7_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid233_In1_c0 <= "" & bh7_w38_9_c0 & bh7_w38_8_c0;
   bh7_w37_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid233_Out0_c0(0);
   bh7_w38_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid233_Out0_c0(1);
   bh7_w39_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid233_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid233: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid233_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid233_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid233_Out0_copy234_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid233_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid233_Out0_copy234_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid235_In0_c0 <= "" & bh7_w39_9_c0 & bh7_w39_8_c0 & bh7_w39_7_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid235_In1_c0 <= "" & bh7_w40_9_c0 & bh7_w40_8_c0;
   bh7_w39_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid235_Out0_c0(0);
   bh7_w40_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid235_Out0_c0(1);
   bh7_w41_8_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid235_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid235: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid235_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid235_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid235_Out0_copy236_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid235_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid235_Out0_copy236_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid237_In0_c0 <= "" & bh7_w41_4_c0 & bh7_w41_7_c0 & bh7_w41_6_c0 & bh7_w41_5_c0;
   Compressor_14_3_Freq300_uid164_bh7_uid237_In1_c0 <= "" & "0";
   bh7_w41_9_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid237_Out0_c0(0);
   bh7_w42_8_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid237_Out0_c0(1);
   bh7_w43_7_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid237_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid237: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid237_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid237_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid237_Out0_copy238_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid237_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid237_Out0_copy238_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid160_bh7_uid239_In0_c0 <= "" & bh7_w42_7_c0 & bh7_w42_6_c0 & bh7_w42_5_c0;
   bh7_w42_9_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid239_Out0_c0(0);
   bh7_w43_8_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid239_Out0_c0(1);
   Compressor_3_2_Freq300_uid160_uid239: Compressor_3_2_Freq300_uid160
      port map ( X0 => Compressor_3_2_Freq300_uid160_bh7_uid239_In0_c0,
                 R => Compressor_3_2_Freq300_uid160_bh7_uid239_Out0_copy240_c0);
   Compressor_3_2_Freq300_uid160_bh7_uid239_Out0_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid239_Out0_copy240_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid241_In0_c0 <= "" & bh7_w43_6_c0 & bh7_w43_5_c0 & bh7_w43_4_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid241_In1_c0 <= "" & bh7_w44_2_c0 & bh7_w44_4_c0;
   bh7_w43_9_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid241_Out0_c0(0);
   bh7_w44_5_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid241_Out0_c0(1);
   bh7_w45_4_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid241_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid241: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid241_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid241_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid241_Out0_copy242_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid241_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid241_Out0_copy242_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid243_In0_c0 <= "" & bh7_w45_3_c0 & bh7_w45_2_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid243_In1_c0 <= "" & bh7_w46_2_c0;
   bh7_w45_5_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid243_Out0_c0(0);
   bh7_w46_3_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid243_Out0_c0(1);
   bh7_w47_1_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid243_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid243: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid243_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid243_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid243_Out0_copy244_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid243_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid243_Out0_copy244_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid245_In0_c0 <= "" & bh7_w22_8_c0 & bh7_w22_7_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid245_In1_c0 <= "" & bh7_w23_10_c0 & bh7_w23_11_c0;
   bh7_w22_9_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid245_Out0_c0(0);
   bh7_w23_12_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid245_Out0_c0(1);
   bh7_w24_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid245_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid245: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid245_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid245_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid245_Out0_copy246_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid245_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid245_Out0_copy246_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid247_In0_c0 <= "" & bh7_w25_11_c0 & bh7_w25_10_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid247_In1_c0 <= "" & bh7_w26_7_c0 & bh7_w26_10_c0;
   bh7_w25_12_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid247_Out0_c0(0);
   bh7_w26_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid247_Out0_c0(1);
   bh7_w27_12_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid247_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid247: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid247_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid247_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid247_Out0_copy248_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid247_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid247_Out0_copy248_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid249_In0_c0 <= "" & bh7_w27_11_c0 & bh7_w27_10_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid249_In1_c0 <= "" & bh7_w28_7_c0 & bh7_w28_10_c0;
   bh7_w27_13_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid249_Out0_c0(0);
   bh7_w28_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid249_Out0_c0(1);
   bh7_w29_12_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid249_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid249: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid249_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid249_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid249_Out0_copy250_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid249_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid249_Out0_copy250_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid251_In0_c0 <= "" & bh7_w29_11_c0 & bh7_w29_10_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid251_In1_c0 <= "" & bh7_w30_7_c0 & bh7_w30_10_c0;
   bh7_w29_13_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid251_Out0_c0(0);
   bh7_w30_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid251_Out0_c0(1);
   bh7_w31_12_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid251_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid251: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid251_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid251_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid251_Out0_copy252_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid251_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid251_Out0_copy252_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid253_In0_c0 <= "" & bh7_w31_11_c0 & bh7_w31_10_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid253_In1_c0 <= "" & bh7_w32_7_c0 & bh7_w32_10_c0;
   bh7_w31_13_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid253_Out0_c0(0);
   bh7_w32_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid253_Out0_c0(1);
   bh7_w33_12_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid253_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid253: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid253_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid253_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid253_Out0_copy254_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid253_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid253_Out0_copy254_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid255_In0_c0 <= "" & bh7_w33_11_c0 & bh7_w33_10_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid255_In1_c0 <= "" & bh7_w34_7_c0 & bh7_w34_10_c0;
   bh7_w33_13_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid255_Out0_c0(0);
   bh7_w34_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid255_Out0_c0(1);
   bh7_w35_12_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid255_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid255: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid255_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid255_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid255_Out0_copy256_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid255_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid255_Out0_copy256_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid257_In0_c0 <= "" & bh7_w35_11_c0 & bh7_w35_10_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid257_In1_c0 <= "" & bh7_w36_7_c0 & bh7_w36_10_c0;
   bh7_w35_13_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid257_Out0_c0(0);
   bh7_w36_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid257_Out0_c0(1);
   bh7_w37_12_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid257_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid257: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid257_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid257_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid257_Out0_copy258_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid257_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid257_Out0_copy258_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid259_In0_c0 <= "" & bh7_w37_11_c0 & bh7_w37_10_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid259_In1_c0 <= "" & bh7_w38_7_c0 & bh7_w38_10_c0;
   bh7_w37_13_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid259_Out0_c0(0);
   bh7_w38_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid259_Out0_c0(1);
   bh7_w39_12_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid259_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid259: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid259_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid259_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid259_Out0_copy260_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid259_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid259_Out0_copy260_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid261_In0_c0 <= "" & bh7_w39_11_c0 & bh7_w39_10_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid261_In1_c0 <= "" & bh7_w40_7_c0 & bh7_w40_10_c0;
   bh7_w39_13_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid261_Out0_c0(0);
   bh7_w40_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid261_Out0_c0(1);
   bh7_w41_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid261_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid261: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid261_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid261_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid261_Out0_copy262_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid261_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid261_Out0_copy262_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid263_In0_c0 <= "" & bh7_w41_9_c0 & bh7_w41_8_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid263_In1_c0 <= "" & bh7_w42_8_c0 & bh7_w42_9_c0;
   bh7_w41_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid263_Out0_c0(0);
   bh7_w42_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid263_Out0_c0(1);
   bh7_w43_10_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid263_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid263: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid263_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid263_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid263_Out0_copy264_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid263_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid263_Out0_copy264_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid265_In0_c0 <= "" & bh7_w43_7_c0 & bh7_w43_9_c0 & bh7_w43_8_c0;
   Compressor_23_3_Freq300_uid156_bh7_uid265_In1_c0 <= "" & bh7_w44_3_c0 & bh7_w44_5_c0;
   bh7_w43_11_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid265_Out0_c0(0);
   bh7_w44_6_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid265_Out0_c0(1);
   bh7_w45_6_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid265_Out0_c0(2);
   Compressor_23_3_Freq300_uid156_uid265: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid265_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid265_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid265_Out0_copy266_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid265_Out0_c0 <= Compressor_23_3_Freq300_uid156_bh7_uid265_Out0_copy266_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid267_In0_c0 <= "" & bh7_w45_5_c0 & bh7_w45_4_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid267_In1_c0 <= "" & bh7_w46_3_c0;
   bh7_w45_7_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid267_Out0_c0(0);
   bh7_w46_4_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid267_Out0_c0(1);
   bh7_w47_2_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid267_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid267: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid267_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid267_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid267_Out0_copy268_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid267_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid267_Out0_copy268_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid160_bh7_uid269_In0_c0 <= "" & bh7_w47_0_c0 & bh7_w47_1_c0 & "0";
   bh7_w47_3_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid269_Out0_c0(0);
   Compressor_3_2_Freq300_uid160_uid269: Compressor_3_2_Freq300_uid160
      port map ( X0 => Compressor_3_2_Freq300_uid160_bh7_uid269_In0_c0,
                 R => Compressor_3_2_Freq300_uid160_bh7_uid269_Out0_copy270_c0);
   Compressor_3_2_Freq300_uid160_bh7_uid269_Out0_c0 <= Compressor_3_2_Freq300_uid160_bh7_uid269_Out0_copy270_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid271_In0_c0 <= "" & bh7_w24_9_c0 & bh7_w24_10_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid271_In1_c0 <= "" & bh7_w25_12_c0;
   bh7_w24_11_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid271_Out0_c0(0);
   bh7_w25_13_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid271_Out0_c0(1);
   bh7_w26_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid271_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid271: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid271_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid271_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid271_Out0_copy272_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid271_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid271_Out0_copy272_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid273_In0_c0 <= "" & bh7_w27_13_c0 & bh7_w27_12_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid273_In1_c0 <= "" & bh7_w28_11_c0;
   bh7_w27_14_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid273_Out0_c0(0);
   bh7_w28_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid273_Out0_c0(1);
   bh7_w29_14_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid273_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid273: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid273_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid273_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid273_Out0_copy274_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid273_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid273_Out0_copy274_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid275_In0_c0 <= "" & bh7_w29_13_c0 & bh7_w29_12_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid275_In1_c0 <= "" & bh7_w30_11_c0;
   bh7_w29_15_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid275_Out0_c0(0);
   bh7_w30_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid275_Out0_c0(1);
   bh7_w31_14_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid275_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid275: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid275_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid275_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid275_Out0_copy276_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid275_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid275_Out0_copy276_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid277_In0_c0 <= "" & bh7_w31_13_c0 & bh7_w31_12_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid277_In1_c0 <= "" & bh7_w32_11_c0;
   bh7_w31_15_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid277_Out0_c0(0);
   bh7_w32_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid277_Out0_c0(1);
   bh7_w33_14_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid277_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid277: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid277_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid277_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid277_Out0_copy278_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid277_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid277_Out0_copy278_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid279_In0_c0 <= "" & bh7_w33_13_c0 & bh7_w33_12_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid279_In1_c0 <= "" & bh7_w34_11_c0;
   bh7_w33_15_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid279_Out0_c0(0);
   bh7_w34_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid279_Out0_c0(1);
   bh7_w35_14_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid279_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid279: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid279_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid279_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid279_Out0_copy280_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid279_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid279_Out0_copy280_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid281_In0_c0 <= "" & bh7_w35_13_c0 & bh7_w35_12_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid281_In1_c0 <= "" & bh7_w36_11_c0;
   bh7_w35_15_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid281_Out0_c0(0);
   bh7_w36_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid281_Out0_c0(1);
   bh7_w37_14_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid281_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid281: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid281_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid281_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid281_Out0_copy282_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid281_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid281_Out0_copy282_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid283_In0_c0 <= "" & bh7_w37_13_c0 & bh7_w37_12_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid283_In1_c0 <= "" & bh7_w38_11_c0;
   bh7_w37_15_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid283_Out0_c0(0);
   bh7_w38_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid283_Out0_c0(1);
   bh7_w39_14_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid283_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid283: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid283_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid283_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid283_Out0_copy284_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid283_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid283_Out0_copy284_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid285_In0_c0 <= "" & bh7_w39_13_c0 & bh7_w39_12_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid285_In1_c0 <= "" & bh7_w40_11_c0;
   bh7_w39_15_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid285_Out0_c0(0);
   bh7_w40_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid285_Out0_c0(1);
   bh7_w41_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid285_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid285: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid285_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid285_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid285_Out0_copy286_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid285_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid285_Out0_copy286_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid287_In0_c0 <= "" & bh7_w41_11_c0 & bh7_w41_10_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid287_In1_c0 <= "" & bh7_w42_10_c0;
   bh7_w41_13_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid287_Out0_c0(0);
   bh7_w42_11_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid287_Out0_c0(1);
   bh7_w43_12_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid287_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid287: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid287_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid287_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid287_Out0_copy288_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid287_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid287_Out0_copy288_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid289_In0_c0 <= "" & bh7_w43_10_c0 & bh7_w43_11_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid289_In1_c0 <= "" & bh7_w44_6_c0;
   bh7_w43_13_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid289_Out0_c0(0);
   bh7_w44_7_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid289_Out0_c0(1);
   bh7_w45_8_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid289_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid289: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid289_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid289_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid289_Out0_copy290_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid289_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid289_Out0_copy290_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid291_In0_c0 <= "" & bh7_w45_6_c0 & bh7_w45_7_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid291_In1_c0 <= "" & bh7_w46_4_c0;
   bh7_w45_9_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid291_Out0_c0(0);
   bh7_w46_5_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid291_Out0_c0(1);
   bh7_w47_4_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid291_Out0_c0(2);
   Compressor_14_3_Freq300_uid164_uid291: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid291_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid291_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid291_Out0_copy292_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid291_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid291_Out0_copy292_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid293_In0_c0 <= "" & bh7_w47_3_c0 & bh7_w47_2_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid293_In1_c0 <= "" & "0";
   bh7_w47_5_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid293_Out0_c0(0);
   Compressor_14_3_Freq300_uid164_uid293: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid293_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid293_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid293_Out0_copy294_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid293_Out0_c0 <= Compressor_14_3_Freq300_uid164_bh7_uid293_Out0_copy294_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid295_In0_c0 <= "" & bh7_w26_11_c0 & bh7_w26_12_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid295_In1_c0 <= "" & bh7_w27_14_c0;
   bh7_w26_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_c1(0);
   bh7_w27_15_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_c1(1);
   bh7_w28_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid295: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid295_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid295_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_copy296_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid295_Out0_copy296_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid297_In0_c0 <= "" & bh7_w29_15_c0 & bh7_w29_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid297_In1_c0 <= "" & bh7_w30_12_c0;
   bh7_w29_16_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_c1(0);
   bh7_w30_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_c1(1);
   bh7_w31_16_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid297: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid297_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid297_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_copy298_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid297_Out0_copy298_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid299_In0_c0 <= "" & bh7_w31_15_c0 & bh7_w31_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid299_In1_c0 <= "" & bh7_w32_12_c0;
   bh7_w31_17_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_c1(0);
   bh7_w32_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_c1(1);
   bh7_w33_16_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid299: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid299_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid299_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_copy300_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid299_Out0_copy300_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid301_In0_c0 <= "" & bh7_w33_15_c0 & bh7_w33_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid301_In1_c0 <= "" & bh7_w34_12_c0;
   bh7_w33_17_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_c1(0);
   bh7_w34_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_c1(1);
   bh7_w35_16_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid301: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid301_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid301_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_copy302_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid301_Out0_copy302_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid303_In0_c0 <= "" & bh7_w35_15_c0 & bh7_w35_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid303_In1_c0 <= "" & bh7_w36_12_c0;
   bh7_w35_17_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_c1(0);
   bh7_w36_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_c1(1);
   bh7_w37_16_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid303: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid303_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid303_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_copy304_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid303_Out0_copy304_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid305_In0_c0 <= "" & bh7_w37_15_c0 & bh7_w37_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid305_In1_c0 <= "" & bh7_w38_12_c0;
   bh7_w37_17_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_c1(0);
   bh7_w38_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_c1(1);
   bh7_w39_16_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid305: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid305_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid305_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_copy306_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid305_Out0_copy306_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid307_In0_c0 <= "" & bh7_w39_15_c0 & bh7_w39_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid307_In1_c0 <= "" & bh7_w40_12_c0;
   bh7_w39_17_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_c1(0);
   bh7_w40_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_c1(1);
   bh7_w41_14_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid307: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid307_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid307_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_copy308_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid307_Out0_copy308_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid309_In0_c0 <= "" & bh7_w41_13_c0 & bh7_w41_12_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid309_In1_c0 <= "" & bh7_w42_11_c0;
   bh7_w41_15_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_c1(0);
   bh7_w42_12_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_c1(1);
   bh7_w43_14_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid309: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid309_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid309_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_copy310_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid309_Out0_copy310_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid311_In0_c0 <= "" & bh7_w43_12_c0 & bh7_w43_13_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid311_In1_c0 <= "" & bh7_w44_7_c0;
   bh7_w43_15_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_c1(0);
   bh7_w44_8_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_c1(1);
   bh7_w45_10_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid311: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid311_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid311_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_copy312_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid311_Out0_copy312_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid313_In0_c0 <= "" & bh7_w45_8_c0 & bh7_w45_9_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid313_In1_c0 <= "" & bh7_w46_5_c0;
   bh7_w45_11_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_c1(0);
   bh7_w46_6_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_c1(1);
   bh7_w47_6_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid313: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid313_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid313_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_copy314_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid313_Out0_copy314_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid315_In0_c0 <= "" & bh7_w47_4_c0 & bh7_w47_5_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid315_In1_c0 <= "" & "0";
   bh7_w47_7_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid315_Out0_c1(0);
   Compressor_14_3_Freq300_uid164_uid315: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid315_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid315_In1_c0,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid315_Out0_copy316_c0);
   Compressor_14_3_Freq300_uid164_bh7_uid315_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid315_Out0_copy316_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid317_In0_c0 <= "" & bh7_w17_1_c0 & bh7_w17_0_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid317_In1_c0 <= "" & bh7_w18_2_c0 & bh7_w18_0_c0;
   bh7_w17_2_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_c1(0);
   bh7_w18_3_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_c1(1);
   bh7_w19_4_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid317: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid317_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid317_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_copy318_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid317_Out0_copy318_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid319_In0_c0 <= "" & bh7_w19_3_c0 & bh7_w19_0_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid319_In1_c0 <= "" & bh7_w20_6_c0 & bh7_w20_0_c0;
   bh7_w19_5_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_c1(0);
   bh7_w20_7_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_c1(1);
   bh7_w21_8_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid319: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid319_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid319_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_copy320_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid319_Out0_copy320_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid321_In0_c0 <= "" & bh7_w21_7_c0 & bh7_w21_0_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid321_In1_c0 <= "" & bh7_w22_9_c0 & bh7_w22_0_c0;
   bh7_w21_9_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_c1(0);
   bh7_w22_10_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_c1(1);
   bh7_w23_13_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid321: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid321_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid321_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_copy322_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid321_Out0_copy322_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid323_In0_c0 <= "" & bh7_w23_12_c0 & bh7_w23_0_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid323_In1_c0 <= "" & bh7_w24_11_c0 & bh7_w24_0_c0;
   bh7_w23_14_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_c1(0);
   bh7_w24_12_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_c1(1);
   bh7_w25_14_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid323: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid323_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid323_In1_c0,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_copy324_c0);
   Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid323_Out0_copy324_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid325_In0_c0 <= "" & bh7_w25_13_c0 & bh7_w25_0_c0 & "0";
   Compressor_23_3_Freq300_uid156_bh7_uid325_In1_c1 <= "" & bh7_w26_0_c1 & bh7_w26_13_c1;
   bh7_w25_15_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid325_Out0_c1(0);
   bh7_w26_14_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid325_Out0_c1(1);
   bh7_w27_16_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid325_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid325: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid325_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid325_In1_c1,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid325_Out0_copy326_c1);
   Compressor_23_3_Freq300_uid156_bh7_uid325_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid325_Out0_copy326_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid160_bh7_uid327_In0_c1 <= "" & bh7_w27_0_c1 & bh7_w27_15_c1 & "0";
   bh7_w27_17_c1 <= Compressor_3_2_Freq300_uid160_bh7_uid327_Out0_c1(0);
   bh7_w28_14_c1 <= Compressor_3_2_Freq300_uid160_bh7_uid327_Out0_c1(1);
   Compressor_3_2_Freq300_uid160_uid327: Compressor_3_2_Freq300_uid160
      port map ( X0 => Compressor_3_2_Freq300_uid160_bh7_uid327_In0_c1,
                 R => Compressor_3_2_Freq300_uid160_bh7_uid327_Out0_copy328_c1);
   Compressor_3_2_Freq300_uid160_bh7_uid327_Out0_c1 <= Compressor_3_2_Freq300_uid160_bh7_uid327_Out0_copy328_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid329_In0_c1 <= "" & bh7_w28_12_c1 & bh7_w28_0_c1 & bh7_w28_13_c1;
   Compressor_23_3_Freq300_uid156_bh7_uid329_In1_c1 <= "" & bh7_w29_0_c1 & bh7_w29_16_c1;
   bh7_w28_15_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid329_Out0_c1(0);
   bh7_w29_17_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid329_Out0_c1(1);
   bh7_w30_14_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid329_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid329: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid329_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid329_In1_c1,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid329_Out0_copy330_c1);
   Compressor_23_3_Freq300_uid156_bh7_uid329_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid329_Out0_copy330_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid160_bh7_uid331_In0_c1 <= "" & bh7_w30_0_c1 & bh7_w30_13_c1 & "0";
   bh7_w30_15_c1 <= Compressor_3_2_Freq300_uid160_bh7_uid331_Out0_c1(0);
   bh7_w31_18_c1 <= Compressor_3_2_Freq300_uid160_bh7_uid331_Out0_c1(1);
   Compressor_3_2_Freq300_uid160_uid331: Compressor_3_2_Freq300_uid160
      port map ( X0 => Compressor_3_2_Freq300_uid160_bh7_uid331_In0_c1,
                 R => Compressor_3_2_Freq300_uid160_bh7_uid331_Out0_copy332_c1);
   Compressor_3_2_Freq300_uid160_bh7_uid331_Out0_c1 <= Compressor_3_2_Freq300_uid160_bh7_uid331_Out0_copy332_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid333_In0_c1 <= "" & bh7_w31_0_c1 & bh7_w31_17_c1 & bh7_w31_16_c1;
   Compressor_23_3_Freq300_uid156_bh7_uid333_In1_c1 <= "" & bh7_w32_0_c1 & bh7_w32_13_c1;
   bh7_w31_19_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid333_Out0_c1(0);
   bh7_w32_14_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid333_Out0_c1(1);
   bh7_w33_18_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid333_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid333: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid333_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid333_In1_c1,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid333_Out0_copy334_c1);
   Compressor_23_3_Freq300_uid156_bh7_uid333_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid333_Out0_copy334_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid335_In0_c1 <= "" & bh7_w33_0_c1 & bh7_w33_17_c1 & bh7_w33_16_c1;
   Compressor_23_3_Freq300_uid156_bh7_uid335_In1_c1 <= "" & bh7_w34_0_c1 & bh7_w34_13_c1;
   bh7_w33_19_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid335_Out0_c1(0);
   bh7_w34_14_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid335_Out0_c1(1);
   bh7_w35_18_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid335_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid335: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid335_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid335_In1_c1,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid335_Out0_copy336_c1);
   Compressor_23_3_Freq300_uid156_bh7_uid335_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid335_Out0_copy336_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid337_In0_c1 <= "" & bh7_w35_0_c1 & bh7_w35_17_c1 & bh7_w35_16_c1;
   Compressor_23_3_Freq300_uid156_bh7_uid337_In1_c1 <= "" & bh7_w36_0_c1 & bh7_w36_13_c1;
   bh7_w35_19_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid337_Out0_c1(0);
   bh7_w36_14_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid337_Out0_c1(1);
   bh7_w37_18_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid337_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid337: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid337_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid337_In1_c1,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid337_Out0_copy338_c1);
   Compressor_23_3_Freq300_uid156_bh7_uid337_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid337_Out0_copy338_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid339_In0_c1 <= "" & bh7_w37_0_c1 & bh7_w37_17_c1 & bh7_w37_16_c1;
   Compressor_23_3_Freq300_uid156_bh7_uid339_In1_c1 <= "" & bh7_w38_0_c1 & bh7_w38_13_c1;
   bh7_w37_19_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid339_Out0_c1(0);
   bh7_w38_14_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid339_Out0_c1(1);
   bh7_w39_18_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid339_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid339: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid339_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid339_In1_c1,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid339_Out0_copy340_c1);
   Compressor_23_3_Freq300_uid156_bh7_uid339_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid339_Out0_copy340_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid156_bh7_uid341_In0_c1 <= "" & bh7_w39_0_c1 & bh7_w39_17_c1 & bh7_w39_16_c1;
   Compressor_23_3_Freq300_uid156_bh7_uid341_In1_c1 <= "" & bh7_w40_0_c1 & bh7_w40_13_c1;
   bh7_w39_19_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid341_Out0_c1(0);
   bh7_w40_14_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid341_Out0_c1(1);
   bh7_w41_16_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid341_Out0_c1(2);
   Compressor_23_3_Freq300_uid156_uid341: Compressor_23_3_Freq300_uid156
      port map ( X0 => Compressor_23_3_Freq300_uid156_bh7_uid341_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid156_bh7_uid341_In1_c1,
                 R => Compressor_23_3_Freq300_uid156_bh7_uid341_Out0_copy342_c1);
   Compressor_23_3_Freq300_uid156_bh7_uid341_Out0_c1 <= Compressor_23_3_Freq300_uid156_bh7_uid341_Out0_copy342_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid343_In0_c1 <= "" & bh7_w41_15_c1 & bh7_w41_14_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid343_In1_c1 <= "" & bh7_w42_12_c1;
   bh7_w41_17_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid343_Out0_c1(0);
   bh7_w42_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid343_Out0_c1(1);
   bh7_w43_16_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid343_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid343: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid343_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid343_In1_c1,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid343_Out0_copy344_c1);
   Compressor_14_3_Freq300_uid164_bh7_uid343_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid343_Out0_copy344_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid345_In0_c1 <= "" & bh7_w43_14_c1 & bh7_w43_15_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid345_In1_c1 <= "" & bh7_w44_8_c1;
   bh7_w43_17_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid345_Out0_c1(0);
   bh7_w44_9_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid345_Out0_c1(1);
   bh7_w45_12_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid345_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid345: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid345_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid345_In1_c1,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid345_Out0_copy346_c1);
   Compressor_14_3_Freq300_uid164_bh7_uid345_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid345_Out0_copy346_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid347_In0_c1 <= "" & bh7_w45_10_c1 & bh7_w45_11_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid347_In1_c1 <= "" & bh7_w46_6_c1;
   bh7_w45_13_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid347_Out0_c1(0);
   bh7_w46_7_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid347_Out0_c1(1);
   bh7_w47_8_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid347_Out0_c1(2);
   Compressor_14_3_Freq300_uid164_uid347: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid347_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid347_In1_c1,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid347_Out0_copy348_c1);
   Compressor_14_3_Freq300_uid164_bh7_uid347_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid347_Out0_copy348_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid164_bh7_uid349_In0_c1 <= "" & bh7_w47_6_c1 & bh7_w47_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid164_bh7_uid349_In1_c0 <= "" & "0";
   bh7_w47_9_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid349_Out0_c1(0);
   Compressor_14_3_Freq300_uid164_uid349: Compressor_14_3_Freq300_uid164
      port map ( X0 => Compressor_14_3_Freq300_uid164_bh7_uid349_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid164_bh7_uid349_In1_c1,
                 R => Compressor_14_3_Freq300_uid164_bh7_uid349_Out0_copy350_c1);
   Compressor_14_3_Freq300_uid164_bh7_uid349_Out0_c1 <= Compressor_14_3_Freq300_uid164_bh7_uid349_Out0_copy350_c1; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh7_18_c1 <= bh7_w18_3_c1 & bh7_w17_2_c1 & bh7_w16_0_c1 & bh7_w15_0_c1 & bh7_w14_0_c1 & bh7_w13_0_c1 & bh7_w12_0_c1 & bh7_w11_0_c1 & bh7_w10_0_c1 & bh7_w9_0_c1 & bh7_w8_0_c1 & bh7_w7_0_c1 & bh7_w6_0_c1 & bh7_w5_0_c1 & bh7_w4_0_c1 & bh7_w3_0_c1 & bh7_w2_0_c1 & bh7_w1_0_c1 & bh7_w0_0_c1;

   bitheapFinalAdd_bh7_In0_c1 <= "0" & bh7_w47_8_c1 & bh7_w46_7_c1 & bh7_w45_12_c1 & bh7_w44_9_c1 & bh7_w43_16_c1 & bh7_w42_13_c1 & bh7_w41_17_c1 & bh7_w40_14_c1 & bh7_w39_19_c1 & bh7_w38_14_c1 & bh7_w37_19_c1 & bh7_w36_14_c1 & bh7_w35_19_c1 & bh7_w34_14_c1 & bh7_w33_19_c1 & bh7_w32_14_c1 & bh7_w31_19_c1 & bh7_w30_15_c1 & bh7_w29_17_c1 & bh7_w28_15_c1 & bh7_w27_17_c1 & bh7_w26_14_c1 & bh7_w25_14_c1 & bh7_w24_12_c1 & bh7_w23_14_c1 & bh7_w22_10_c1 & bh7_w21_9_c1 & bh7_w20_7_c1 & bh7_w19_5_c1;
   bitheapFinalAdd_bh7_In1_c1 <= "0" & bh7_w47_9_c1 & "0" & bh7_w45_13_c1 & "0" & bh7_w43_17_c1 & "0" & bh7_w41_16_c1 & "0" & bh7_w39_18_c1 & "0" & bh7_w37_18_c1 & "0" & bh7_w35_18_c1 & "0" & bh7_w33_18_c1 & "0" & bh7_w31_18_c1 & bh7_w30_14_c1 & "0" & bh7_w28_14_c1 & bh7_w27_16_c1 & "0" & bh7_w25_15_c1 & "0" & bh7_w23_13_c1 & "0" & bh7_w21_8_c1 & "0" & bh7_w19_4_c1;
   bitheapFinalAdd_bh7_Cin_c0 <= '0';

   bitheapFinalAdd_bh7: IntAdder_30_Freq300_uid352
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 Cin => bitheapFinalAdd_bh7_Cin_c0,
                 X => bitheapFinalAdd_bh7_In0_c1,
                 Y => bitheapFinalAdd_bh7_In1_c1,
                 R => bitheapFinalAdd_bh7_Out_c1);
   bitheapResult_bh7_c1 <= bitheapFinalAdd_bh7_Out_c1(28 downto 0) & tmp_bitheapResult_bh7_18_c1;
   R <= bitheapResult_bh7_c1(47 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_33_Freq300_uid355
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_33_Freq300_uid355 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(32 downto 0);
          Y : in  std_logic_vector(32 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(32 downto 0)   );
end entity;

architecture arch of IntAdder_33_Freq300_uid355 is
signal Rtmp_c2 :  std_logic_vector(32 downto 0);
signal X_c2 :  std_logic_vector(32 downto 0);
signal Y_c1, Y_c2 :  std_logic_vector(32 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_c1 <= Y;
            end if;
            if ce_2 = '1' then
               X_c2 <= X;
               Y_c2 <= Y_c1;
            end if;
         end if;
      end process;
   Rtmp_c2 <= X_c2 + Y_c2 + Cin;
   R <= Rtmp_c2;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointMultiplier
--                      (FPMult_8_23_uid2_Freq300_uid3)
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointMultiplier_32_2_875333 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointMultiplier_32_2_875333 is
   component IntMultiplier_24x24_48_Freq300_uid5 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_Freq300_uid355 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(32 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(32 downto 0)   );
   end component;

signal sign_c0, sign_c1, sign_c2 :  std_logic;
signal expX_c0 :  std_logic_vector(7 downto 0);
signal expY_c0 :  std_logic_vector(7 downto 0);
signal expSumPreSub_c0 :  std_logic_vector(9 downto 0);
signal bias_c0 :  std_logic_vector(9 downto 0);
signal expSum_c0, expSum_c1 :  std_logic_vector(9 downto 0);
signal sigX_c0 :  std_logic_vector(23 downto 0);
signal sigY_c0 :  std_logic_vector(23 downto 0);
signal sigProd_c1 :  std_logic_vector(47 downto 0);
signal excSel_c0 :  std_logic_vector(3 downto 0);
signal exc_c0, exc_c1, exc_c2 :  std_logic_vector(1 downto 0);
signal norm_c1 :  std_logic;
signal expPostNorm_c1 :  std_logic_vector(9 downto 0);
signal sigProdExt_c1, sigProdExt_c2 :  std_logic_vector(47 downto 0);
signal expSig_c1 :  std_logic_vector(32 downto 0);
signal sticky_c1, sticky_c2 :  std_logic;
signal guard_c2 :  std_logic;
signal round_c2 :  std_logic;
signal expSigPostRound_c2 :  std_logic_vector(32 downto 0);
signal excPostNorm_c2 :  std_logic_vector(1 downto 0);
signal finalExc_c2 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               sign_c1 <= sign_c0;
               expSum_c1 <= expSum_c0;
               exc_c1 <= exc_c0;
            end if;
            if ce_2 = '1' then
               sign_c2 <= sign_c1;
               exc_c2 <= exc_c1;
               sigProdExt_c2 <= sigProdExt_c1;
               sticky_c2 <= sticky_c1;
            end if;
         end if;
      end process;
   sign_c0 <= X(31) xor Y(31);
   expX_c0 <= X(30 downto 23);
   expY_c0 <= Y(30 downto 23);
   expSumPreSub_c0 <= ("00" & expX_c0) + ("00" & expY_c0);
   bias_c0 <= CONV_STD_LOGIC_VECTOR(127,10);
   expSum_c0 <= expSumPreSub_c0 - bias_c0;
   sigX_c0 <= "1" & X(22 downto 0);
   sigY_c0 <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_24x24_48_Freq300_uid5
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 X => sigX_c0,
                 Y => sigY_c0,
                 R => sigProd_c1);
   excSel_c0 <= X(33 downto 32) & Y(33 downto 32);
   with excSel_c0  select  
   exc_c0 <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm_c1 <= sigProd_c1(47);
   -- exponent update
   expPostNorm_c1 <= expSum_c1 + ("000000000" & norm_c1);
   -- significand normalization shift
   sigProdExt_c1 <= sigProd_c1(46 downto 0) & "0" when norm_c1='1' else
                         sigProd_c1(45 downto 0) & "00";
   expSig_c1 <= expPostNorm_c1 & sigProdExt_c1(47 downto 25);
   sticky_c1 <= sigProdExt_c1(24);
   guard_c2 <= '0' when sigProdExt_c2(23 downto 0)="000000000000000000000000" else '1';
   round_c2 <= sticky_c2 and ( (guard_c2 and not(sigProdExt_c2(25))) or (sigProdExt_c2(25) ))  ;
   RoundingAdder: IntAdder_33_Freq300_uid355
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 Cin => round_c2,
                 X => expSig_c1,
                 Y => "000000000000000000000000000000000",
                 R => expSigPostRound_c2);
   with expSigPostRound_c2(32 downto 31)  select 
   excPostNorm_c2 <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_c2  select  
   finalExc_c2 <= exc_c2 when  "11"|"10"|"00",
                       excPostNorm_c2 when others; 
   R <= finalExc_c2 & sign_c2 & expSigPostRound_c2(30 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid17
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid17 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid17 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid22
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid22 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid22 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid27
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid27 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid27 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid32
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid32 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid32 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid37
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid37 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid37 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid42
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid42 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid42 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid47
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid47 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid47 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid52
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid52 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid52 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid63
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid63 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid63 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid68
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid68 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid68 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid73
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid73 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid73 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid78
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid78 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid78 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid83
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid83 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid83 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid88
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid88 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid88 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid93
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid93 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid93 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid98
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid98 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid98 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid113
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid113 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid113 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid118
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid118 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid118 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid123
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid128
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid128 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid128 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid133
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid133 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid133 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid138
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid138 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid138 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid143
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid143 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid143 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid148
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid148 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid148 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid153
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid153 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid153 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid158
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid158 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid158 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid163
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid163 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid163 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid168
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid168 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid168 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid183
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid183 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid183 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid188
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid188 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid188 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid193
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid193 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid193 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid198
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid198 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid198 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid203
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid203 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid203 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid208
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid208 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid208 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid213
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid213 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid213 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid218
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid218 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid218 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid223
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid223 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid223 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid228
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid228 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid228 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid233
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid233 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid233 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid238
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid238 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid238 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid253
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid253 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid253 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid258
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid258 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid258 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid263
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid263 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid263 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid268
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid268 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid268 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid273
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid273 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid273 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid278
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid278 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid278 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid283
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid283 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid283 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid288
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid288 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid288 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid293
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid293 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid293 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid298
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid298 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid298 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid303
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid303 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid303 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid308
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid308 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid308 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid313
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid313 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid313 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq800_uid318
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq800_uid318 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq800_uid318 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq800_uid322
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq800_uid322 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq800_uid322 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq800_uid326
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq800_uid326 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq800_uid326 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq800_uid334
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq800_uid334 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq800_uid334 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq800_uid400
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq800_uid400 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq800_uid400 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq800_uid432
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq800_uid432 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq800_uid432 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid9
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid9 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid9 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid11
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid11 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid11 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid13
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid13 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid13 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid15
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid15 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid15 is
   component MultTable_Freq800_uid17 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy18_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid17
      port map ( X => Xtable_c0,
                 Y => Y1_copy18_c0);
   Y1_c0 <= Y1_copy18_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid20
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid20 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid20 is
   component MultTable_Freq800_uid22 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy23_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid22
      port map ( X => Xtable_c0,
                 Y => Y1_copy23_c0);
   Y1_c0 <= Y1_copy23_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid25
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid25 is
   component MultTable_Freq800_uid27 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy28_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid27
      port map ( X => Xtable_c0,
                 Y => Y1_copy28_c0);
   Y1_c0 <= Y1_copy28_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid30
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid30 is
   component MultTable_Freq800_uid32 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy33_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid32
      port map ( X => Xtable_c0,
                 Y => Y1_copy33_c0);
   Y1_c0 <= Y1_copy33_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid35
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid35 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid35 is
   component MultTable_Freq800_uid37 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy38_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid37
      port map ( X => Xtable_c0,
                 Y => Y1_copy38_c0);
   Y1_c0 <= Y1_copy38_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid40
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid40 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid40 is
   component MultTable_Freq800_uid42 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy43_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid42
      port map ( X => Xtable_c0,
                 Y => Y1_copy43_c0);
   Y1_c0 <= Y1_copy43_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid45
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid45 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid45 is
   component MultTable_Freq800_uid47 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy48_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid47
      port map ( X => Xtable_c0,
                 Y => Y1_copy48_c0);
   Y1_c0 <= Y1_copy48_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid50
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid50 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid50 is
   component MultTable_Freq800_uid52 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy53_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid52
      port map ( X => Xtable_c0,
                 Y => Y1_copy53_c0);
   Y1_c0 <= Y1_copy53_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid55
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid55 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid55 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid57
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid57 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid57 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq800_uid59
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq800_uid59 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq800_uid59 is
signal Mfull_c0, Mfull_c1, Mfull_c2 :  std_logic_vector(40 downto 0);
signal M_c2 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
            if ce_2 = '1' then
               Mfull_c2 <= Mfull_c1;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c2 <= Mfull_c2(40 downto 0);
   R <= M_c2;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid61
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid61 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid61 is
   component MultTable_Freq800_uid63 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy64_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid63
      port map ( X => Xtable_c0,
                 Y => Y1_copy64_c0);
   Y1_c0 <= Y1_copy64_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid66
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid66 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid66 is
   component MultTable_Freq800_uid68 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy69_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid68
      port map ( X => Xtable_c0,
                 Y => Y1_copy69_c0);
   Y1_c0 <= Y1_copy69_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid71
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid71 is
   component MultTable_Freq800_uid73 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy74_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid73
      port map ( X => Xtable_c0,
                 Y => Y1_copy74_c0);
   Y1_c0 <= Y1_copy74_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid76
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid76 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid76 is
   component MultTable_Freq800_uid78 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy79_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid78
      port map ( X => Xtable_c0,
                 Y => Y1_copy79_c0);
   Y1_c0 <= Y1_copy79_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid81
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid81 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid81 is
   component MultTable_Freq800_uid83 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy84_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid83
      port map ( X => Xtable_c0,
                 Y => Y1_copy84_c0);
   Y1_c0 <= Y1_copy84_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid86
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid86 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid86 is
   component MultTable_Freq800_uid88 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy89_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid88
      port map ( X => Xtable_c0,
                 Y => Y1_copy89_c0);
   Y1_c0 <= Y1_copy89_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid91
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid91 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid91 is
   component MultTable_Freq800_uid93 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy94_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid93
      port map ( X => Xtable_c0,
                 Y => Y1_copy94_c0);
   Y1_c0 <= Y1_copy94_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq800_uid96
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid96 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid96 is
   component MultTable_Freq800_uid98 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy99_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid98
      port map ( X => Xtable_c0,
                 Y => Y1_copy99_c0);
   Y1_c0 <= Y1_copy99_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq800_uid101
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid101 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid101 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid103
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid103 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid103 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid105
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid105 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid105 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid107
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid107 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid107 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid109
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid109 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid109 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid111
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid111 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid111 is
   component MultTable_Freq800_uid113 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy114_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid113
      port map ( X => Xtable_c0,
                 Y => Y1_copy114_c0);
   Y1_c0 <= Y1_copy114_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid116
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid116 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid116 is
   component MultTable_Freq800_uid118 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy119_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid118
      port map ( X => Xtable_c0,
                 Y => Y1_copy119_c0);
   Y1_c0 <= Y1_copy119_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid121
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid121 is
   component MultTable_Freq800_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy124_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid123
      port map ( X => Xtable_c0,
                 Y => Y1_copy124_c0);
   Y1_c0 <= Y1_copy124_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid126
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid126 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid126 is
   component MultTable_Freq800_uid128 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy129_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid128
      port map ( X => Xtable_c0,
                 Y => Y1_copy129_c0);
   Y1_c0 <= Y1_copy129_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid131
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid131 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid131 is
   component MultTable_Freq800_uid133 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy134_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid133
      port map ( X => Xtable_c0,
                 Y => Y1_copy134_c0);
   Y1_c0 <= Y1_copy134_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid136
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid136 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid136 is
   component MultTable_Freq800_uid138 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy139_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid138
      port map ( X => Xtable_c0,
                 Y => Y1_copy139_c0);
   Y1_c0 <= Y1_copy139_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid141
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid141 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid141 is
   component MultTable_Freq800_uid143 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy144_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid143
      port map ( X => Xtable_c0,
                 Y => Y1_copy144_c0);
   Y1_c0 <= Y1_copy144_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid146
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid146 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid146 is
   component MultTable_Freq800_uid148 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy149_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid148
      port map ( X => Xtable_c0,
                 Y => Y1_copy149_c0);
   Y1_c0 <= Y1_copy149_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid151
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid151 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid151 is
   component MultTable_Freq800_uid153 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy154_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid153
      port map ( X => Xtable_c0,
                 Y => Y1_copy154_c0);
   Y1_c0 <= Y1_copy154_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid156
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid156 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid156 is
   component MultTable_Freq800_uid158 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy159_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid158
      port map ( X => Xtable_c0,
                 Y => Y1_copy159_c0);
   Y1_c0 <= Y1_copy159_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid161
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid161 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid161 is
   component MultTable_Freq800_uid163 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy164_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid163
      port map ( X => Xtable_c0,
                 Y => Y1_copy164_c0);
   Y1_c0 <= Y1_copy164_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid166
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid166 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid166 is
   component MultTable_Freq800_uid168 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy169_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid168
      port map ( X => Xtable_c0,
                 Y => Y1_copy169_c0);
   Y1_c0 <= Y1_copy169_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq800_uid171
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid171 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid171 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid173
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid173 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid173 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid175
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid175 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid175 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid177
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid177 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid177 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid179
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid179 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid179 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid181
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid181 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid181 is
   component MultTable_Freq800_uid183 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy184_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid183
      port map ( X => Xtable_c0,
                 Y => Y1_copy184_c0);
   Y1_c0 <= Y1_copy184_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid186
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid186 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid186 is
   component MultTable_Freq800_uid188 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy189_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid188
      port map ( X => Xtable_c0,
                 Y => Y1_copy189_c0);
   Y1_c0 <= Y1_copy189_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid191
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid191 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid191 is
   component MultTable_Freq800_uid193 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy194_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid193
      port map ( X => Xtable_c0,
                 Y => Y1_copy194_c0);
   Y1_c0 <= Y1_copy194_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid196
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid196 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid196 is
   component MultTable_Freq800_uid198 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy199_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid198
      port map ( X => Xtable_c0,
                 Y => Y1_copy199_c0);
   Y1_c0 <= Y1_copy199_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid201
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid201 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid201 is
   component MultTable_Freq800_uid203 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy204_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid203
      port map ( X => Xtable_c0,
                 Y => Y1_copy204_c0);
   Y1_c0 <= Y1_copy204_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid206
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid206 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid206 is
   component MultTable_Freq800_uid208 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy209_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid208
      port map ( X => Xtable_c0,
                 Y => Y1_copy209_c0);
   Y1_c0 <= Y1_copy209_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid211
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid211 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid211 is
   component MultTable_Freq800_uid213 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy214_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid213
      port map ( X => Xtable_c0,
                 Y => Y1_copy214_c0);
   Y1_c0 <= Y1_copy214_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid216
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid216 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid216 is
   component MultTable_Freq800_uid218 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy219_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid218
      port map ( X => Xtable_c0,
                 Y => Y1_copy219_c0);
   Y1_c0 <= Y1_copy219_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid221
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid221 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid221 is
   component MultTable_Freq800_uid223 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy224_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid223
      port map ( X => Xtable_c0,
                 Y => Y1_copy224_c0);
   Y1_c0 <= Y1_copy224_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid226
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid226 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid226 is
   component MultTable_Freq800_uid228 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy229_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid228
      port map ( X => Xtable_c0,
                 Y => Y1_copy229_c0);
   Y1_c0 <= Y1_copy229_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid231
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid231 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid231 is
   component MultTable_Freq800_uid233 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy234_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid233
      port map ( X => Xtable_c0,
                 Y => Y1_copy234_c0);
   Y1_c0 <= Y1_copy234_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid236
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid236 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid236 is
   component MultTable_Freq800_uid238 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy239_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid238
      port map ( X => Xtable_c0,
                 Y => Y1_copy239_c0);
   Y1_c0 <= Y1_copy239_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq800_uid241
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq800_uid241 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq800_uid241 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid243
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid243 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid243 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid245
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid245 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid245 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid247
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid247 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid247 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq800_uid249
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq800_uid249 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq800_uid249 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid251
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid251 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid251 is
   component MultTable_Freq800_uid253 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy254_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid253
      port map ( X => Xtable_c0,
                 Y => Y1_copy254_c0);
   Y1_c0 <= Y1_copy254_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid256
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid256 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid256 is
   component MultTable_Freq800_uid258 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy259_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid258
      port map ( X => Xtable_c0,
                 Y => Y1_copy259_c0);
   Y1_c0 <= Y1_copy259_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid261
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid261 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid261 is
   component MultTable_Freq800_uid263 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy264_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid263
      port map ( X => Xtable_c0,
                 Y => Y1_copy264_c0);
   Y1_c0 <= Y1_copy264_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid266
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid266 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid266 is
   component MultTable_Freq800_uid268 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy269_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid268
      port map ( X => Xtable_c0,
                 Y => Y1_copy269_c0);
   Y1_c0 <= Y1_copy269_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid271
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid271 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid271 is
   component MultTable_Freq800_uid273 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy274_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid273
      port map ( X => Xtable_c0,
                 Y => Y1_copy274_c0);
   Y1_c0 <= Y1_copy274_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid276
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid276 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid276 is
   component MultTable_Freq800_uid278 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy279_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid278
      port map ( X => Xtable_c0,
                 Y => Y1_copy279_c0);
   Y1_c0 <= Y1_copy279_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid281
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid281 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid281 is
   component MultTable_Freq800_uid283 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy284_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid283
      port map ( X => Xtable_c0,
                 Y => Y1_copy284_c0);
   Y1_c0 <= Y1_copy284_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid286
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid286 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid286 is
   component MultTable_Freq800_uid288 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy289_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid288
      port map ( X => Xtable_c0,
                 Y => Y1_copy289_c0);
   Y1_c0 <= Y1_copy289_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid291
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid291 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid291 is
   component MultTable_Freq800_uid293 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy294_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid293
      port map ( X => Xtable_c0,
                 Y => Y1_copy294_c0);
   Y1_c0 <= Y1_copy294_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid296
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid296 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid296 is
   component MultTable_Freq800_uid298 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy299_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid298
      port map ( X => Xtable_c0,
                 Y => Y1_copy299_c0);
   Y1_c0 <= Y1_copy299_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid301
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid301 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid301 is
   component MultTable_Freq800_uid303 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy304_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid303
      port map ( X => Xtable_c0,
                 Y => Y1_copy304_c0);
   Y1_c0 <= Y1_copy304_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq800_uid306
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq800_uid306 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq800_uid306 is
   component MultTable_Freq800_uid308 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy309_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid308
      port map ( X => Xtable_c0,
                 Y => Y1_copy309_c0);
   Y1_c0 <= Y1_copy309_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq800_uid311
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq800_uid311 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq800_uid311 is
   component MultTable_Freq800_uid313 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy314_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid313
      port map ( X => Xtable_c0,
                 Y => Y1_copy314_c0);
   Y1_c0 <= Y1_copy314_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x3_Freq800_uid316
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq800_uid316 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq800_uid316 is
   component MultTable_Freq800_uid318 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy319_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq800_uid318
      port map ( X => Xtable_c0,
                 Y => Y1_copy319_c0);
   Y1_c0 <= Y1_copy319_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_84_Freq800_uid972
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 33 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_84_Freq800_uid972 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33 : in std_logic;
          X : in  std_logic_vector(83 downto 0);
          Y : in  std_logic_vector(83 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(83 downto 0)   );
end entity;

architecture arch of IntAdder_84_Freq800_uid972 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3, Cin_0_c4, Cin_0_c5 :  std_logic;
signal X_0_c4, X_0_c5 :  std_logic_vector(3 downto 0);
signal Y_0_c4, Y_0_c5 :  std_logic_vector(3 downto 0);
signal S_0_c5 :  std_logic_vector(3 downto 0);
signal R_0_c5, R_0_c6, R_0_c7, R_0_c8, R_0_c9, R_0_c10, R_0_c11, R_0_c12, R_0_c13, R_0_c14, R_0_c15, R_0_c16, R_0_c17, R_0_c18, R_0_c19, R_0_c20, R_0_c21, R_0_c22, R_0_c23, R_0_c24, R_0_c25, R_0_c26, R_0_c27, R_0_c28, R_0_c29, R_0_c30, R_0_c31, R_0_c32, R_0_c33 :  std_logic_vector(2 downto 0);
signal Cin_1_c5, Cin_1_c6 :  std_logic;
signal X_1_c4, X_1_c5, X_1_c6 :  std_logic_vector(3 downto 0);
signal Y_1_c4, Y_1_c5, Y_1_c6 :  std_logic_vector(3 downto 0);
signal S_1_c6 :  std_logic_vector(3 downto 0);
signal R_1_c6, R_1_c7, R_1_c8, R_1_c9, R_1_c10, R_1_c11, R_1_c12, R_1_c13, R_1_c14, R_1_c15, R_1_c16, R_1_c17, R_1_c18, R_1_c19, R_1_c20, R_1_c21, R_1_c22, R_1_c23, R_1_c24, R_1_c25, R_1_c26, R_1_c27, R_1_c28, R_1_c29, R_1_c30, R_1_c31, R_1_c32, R_1_c33 :  std_logic_vector(2 downto 0);
signal Cin_2_c6, Cin_2_c7 :  std_logic;
signal X_2_c4, X_2_c5, X_2_c6, X_2_c7 :  std_logic_vector(3 downto 0);
signal Y_2_c4, Y_2_c5, Y_2_c6, Y_2_c7 :  std_logic_vector(3 downto 0);
signal S_2_c7 :  std_logic_vector(3 downto 0);
signal R_2_c7, R_2_c8, R_2_c9, R_2_c10, R_2_c11, R_2_c12, R_2_c13, R_2_c14, R_2_c15, R_2_c16, R_2_c17, R_2_c18, R_2_c19, R_2_c20, R_2_c21, R_2_c22, R_2_c23, R_2_c24, R_2_c25, R_2_c26, R_2_c27, R_2_c28, R_2_c29, R_2_c30, R_2_c31, R_2_c32, R_2_c33 :  std_logic_vector(2 downto 0);
signal Cin_3_c7, Cin_3_c8 :  std_logic;
signal X_3_c4, X_3_c5, X_3_c6, X_3_c7, X_3_c8 :  std_logic_vector(3 downto 0);
signal Y_3_c4, Y_3_c5, Y_3_c6, Y_3_c7, Y_3_c8 :  std_logic_vector(3 downto 0);
signal S_3_c8 :  std_logic_vector(3 downto 0);
signal R_3_c8, R_3_c9, R_3_c10, R_3_c11, R_3_c12, R_3_c13, R_3_c14, R_3_c15, R_3_c16, R_3_c17, R_3_c18, R_3_c19, R_3_c20, R_3_c21, R_3_c22, R_3_c23, R_3_c24, R_3_c25, R_3_c26, R_3_c27, R_3_c28, R_3_c29, R_3_c30, R_3_c31, R_3_c32, R_3_c33 :  std_logic_vector(2 downto 0);
signal Cin_4_c8, Cin_4_c9 :  std_logic;
signal X_4_c4, X_4_c5, X_4_c6, X_4_c7, X_4_c8, X_4_c9 :  std_logic_vector(3 downto 0);
signal Y_4_c4, Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8, Y_4_c9 :  std_logic_vector(3 downto 0);
signal S_4_c9 :  std_logic_vector(3 downto 0);
signal R_4_c9, R_4_c10, R_4_c11, R_4_c12, R_4_c13, R_4_c14, R_4_c15, R_4_c16, R_4_c17, R_4_c18, R_4_c19, R_4_c20, R_4_c21, R_4_c22, R_4_c23, R_4_c24, R_4_c25, R_4_c26, R_4_c27, R_4_c28, R_4_c29, R_4_c30, R_4_c31, R_4_c32, R_4_c33 :  std_logic_vector(2 downto 0);
signal Cin_5_c9, Cin_5_c10 :  std_logic;
signal X_5_c4, X_5_c5, X_5_c6, X_5_c7, X_5_c8, X_5_c9, X_5_c10 :  std_logic_vector(3 downto 0);
signal Y_5_c4, Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9, Y_5_c10 :  std_logic_vector(3 downto 0);
signal S_5_c10 :  std_logic_vector(3 downto 0);
signal R_5_c10, R_5_c11, R_5_c12, R_5_c13, R_5_c14, R_5_c15, R_5_c16, R_5_c17, R_5_c18, R_5_c19, R_5_c20, R_5_c21, R_5_c22, R_5_c23, R_5_c24, R_5_c25, R_5_c26, R_5_c27, R_5_c28, R_5_c29, R_5_c30, R_5_c31, R_5_c32, R_5_c33 :  std_logic_vector(2 downto 0);
signal Cin_6_c10, Cin_6_c11 :  std_logic;
signal X_6_c4, X_6_c5, X_6_c6, X_6_c7, X_6_c8, X_6_c9, X_6_c10, X_6_c11 :  std_logic_vector(3 downto 0);
signal Y_6_c4, Y_6_c5, Y_6_c6, Y_6_c7, Y_6_c8, Y_6_c9, Y_6_c10, Y_6_c11 :  std_logic_vector(3 downto 0);
signal S_6_c11 :  std_logic_vector(3 downto 0);
signal R_6_c11, R_6_c12, R_6_c13, R_6_c14, R_6_c15, R_6_c16, R_6_c17, R_6_c18, R_6_c19, R_6_c20, R_6_c21, R_6_c22, R_6_c23, R_6_c24, R_6_c25, R_6_c26, R_6_c27, R_6_c28, R_6_c29, R_6_c30, R_6_c31, R_6_c32, R_6_c33 :  std_logic_vector(2 downto 0);
signal Cin_7_c11, Cin_7_c12 :  std_logic;
signal X_7_c4, X_7_c5, X_7_c6, X_7_c7, X_7_c8, X_7_c9, X_7_c10, X_7_c11, X_7_c12 :  std_logic_vector(3 downto 0);
signal Y_7_c4, Y_7_c5, Y_7_c6, Y_7_c7, Y_7_c8, Y_7_c9, Y_7_c10, Y_7_c11, Y_7_c12 :  std_logic_vector(3 downto 0);
signal S_7_c12 :  std_logic_vector(3 downto 0);
signal R_7_c12, R_7_c13, R_7_c14, R_7_c15, R_7_c16, R_7_c17, R_7_c18, R_7_c19, R_7_c20, R_7_c21, R_7_c22, R_7_c23, R_7_c24, R_7_c25, R_7_c26, R_7_c27, R_7_c28, R_7_c29, R_7_c30, R_7_c31, R_7_c32, R_7_c33 :  std_logic_vector(2 downto 0);
signal Cin_8_c12, Cin_8_c13 :  std_logic;
signal X_8_c4, X_8_c5, X_8_c6, X_8_c7, X_8_c8, X_8_c9, X_8_c10, X_8_c11, X_8_c12, X_8_c13 :  std_logic_vector(3 downto 0);
signal Y_8_c4, Y_8_c5, Y_8_c6, Y_8_c7, Y_8_c8, Y_8_c9, Y_8_c10, Y_8_c11, Y_8_c12, Y_8_c13 :  std_logic_vector(3 downto 0);
signal S_8_c13 :  std_logic_vector(3 downto 0);
signal R_8_c13, R_8_c14, R_8_c15, R_8_c16, R_8_c17, R_8_c18, R_8_c19, R_8_c20, R_8_c21, R_8_c22, R_8_c23, R_8_c24, R_8_c25, R_8_c26, R_8_c27, R_8_c28, R_8_c29, R_8_c30, R_8_c31, R_8_c32, R_8_c33 :  std_logic_vector(2 downto 0);
signal Cin_9_c13, Cin_9_c14 :  std_logic;
signal X_9_c4, X_9_c5, X_9_c6, X_9_c7, X_9_c8, X_9_c9, X_9_c10, X_9_c11, X_9_c12, X_9_c13, X_9_c14 :  std_logic_vector(3 downto 0);
signal Y_9_c4, Y_9_c5, Y_9_c6, Y_9_c7, Y_9_c8, Y_9_c9, Y_9_c10, Y_9_c11, Y_9_c12, Y_9_c13, Y_9_c14 :  std_logic_vector(3 downto 0);
signal S_9_c14 :  std_logic_vector(3 downto 0);
signal R_9_c14, R_9_c15, R_9_c16, R_9_c17, R_9_c18, R_9_c19, R_9_c20, R_9_c21, R_9_c22, R_9_c23, R_9_c24, R_9_c25, R_9_c26, R_9_c27, R_9_c28, R_9_c29, R_9_c30, R_9_c31, R_9_c32, R_9_c33 :  std_logic_vector(2 downto 0);
signal Cin_10_c14, Cin_10_c15 :  std_logic;
signal X_10_c4, X_10_c5, X_10_c6, X_10_c7, X_10_c8, X_10_c9, X_10_c10, X_10_c11, X_10_c12, X_10_c13, X_10_c14, X_10_c15 :  std_logic_vector(3 downto 0);
signal Y_10_c4, Y_10_c5, Y_10_c6, Y_10_c7, Y_10_c8, Y_10_c9, Y_10_c10, Y_10_c11, Y_10_c12, Y_10_c13, Y_10_c14, Y_10_c15 :  std_logic_vector(3 downto 0);
signal S_10_c15 :  std_logic_vector(3 downto 0);
signal R_10_c15, R_10_c16, R_10_c17, R_10_c18, R_10_c19, R_10_c20, R_10_c21, R_10_c22, R_10_c23, R_10_c24, R_10_c25, R_10_c26, R_10_c27, R_10_c28, R_10_c29, R_10_c30, R_10_c31, R_10_c32, R_10_c33 :  std_logic_vector(2 downto 0);
signal Cin_11_c15, Cin_11_c16 :  std_logic;
signal X_11_c4, X_11_c5, X_11_c6, X_11_c7, X_11_c8, X_11_c9, X_11_c10, X_11_c11, X_11_c12, X_11_c13, X_11_c14, X_11_c15, X_11_c16 :  std_logic_vector(3 downto 0);
signal Y_11_c4, Y_11_c5, Y_11_c6, Y_11_c7, Y_11_c8, Y_11_c9, Y_11_c10, Y_11_c11, Y_11_c12, Y_11_c13, Y_11_c14, Y_11_c15, Y_11_c16 :  std_logic_vector(3 downto 0);
signal S_11_c16 :  std_logic_vector(3 downto 0);
signal R_11_c16, R_11_c17, R_11_c18, R_11_c19, R_11_c20, R_11_c21, R_11_c22, R_11_c23, R_11_c24, R_11_c25, R_11_c26, R_11_c27, R_11_c28, R_11_c29, R_11_c30, R_11_c31, R_11_c32, R_11_c33 :  std_logic_vector(2 downto 0);
signal Cin_12_c16, Cin_12_c17 :  std_logic;
signal X_12_c4, X_12_c5, X_12_c6, X_12_c7, X_12_c8, X_12_c9, X_12_c10, X_12_c11, X_12_c12, X_12_c13, X_12_c14, X_12_c15, X_12_c16, X_12_c17 :  std_logic_vector(3 downto 0);
signal Y_12_c4, Y_12_c5, Y_12_c6, Y_12_c7, Y_12_c8, Y_12_c9, Y_12_c10, Y_12_c11, Y_12_c12, Y_12_c13, Y_12_c14, Y_12_c15, Y_12_c16, Y_12_c17 :  std_logic_vector(3 downto 0);
signal S_12_c17 :  std_logic_vector(3 downto 0);
signal R_12_c17, R_12_c18, R_12_c19, R_12_c20, R_12_c21, R_12_c22, R_12_c23, R_12_c24, R_12_c25, R_12_c26, R_12_c27, R_12_c28, R_12_c29, R_12_c30, R_12_c31, R_12_c32, R_12_c33 :  std_logic_vector(2 downto 0);
signal Cin_13_c17, Cin_13_c18 :  std_logic;
signal X_13_c4, X_13_c5, X_13_c6, X_13_c7, X_13_c8, X_13_c9, X_13_c10, X_13_c11, X_13_c12, X_13_c13, X_13_c14, X_13_c15, X_13_c16, X_13_c17, X_13_c18 :  std_logic_vector(3 downto 0);
signal Y_13_c4, Y_13_c5, Y_13_c6, Y_13_c7, Y_13_c8, Y_13_c9, Y_13_c10, Y_13_c11, Y_13_c12, Y_13_c13, Y_13_c14, Y_13_c15, Y_13_c16, Y_13_c17, Y_13_c18 :  std_logic_vector(3 downto 0);
signal S_13_c18 :  std_logic_vector(3 downto 0);
signal R_13_c18, R_13_c19, R_13_c20, R_13_c21, R_13_c22, R_13_c23, R_13_c24, R_13_c25, R_13_c26, R_13_c27, R_13_c28, R_13_c29, R_13_c30, R_13_c31, R_13_c32, R_13_c33 :  std_logic_vector(2 downto 0);
signal Cin_14_c18, Cin_14_c19, Cin_14_c20 :  std_logic;
signal X_14_c4, X_14_c5, X_14_c6, X_14_c7, X_14_c8, X_14_c9, X_14_c10, X_14_c11, X_14_c12, X_14_c13, X_14_c14, X_14_c15, X_14_c16, X_14_c17, X_14_c18, X_14_c19, X_14_c20 :  std_logic_vector(3 downto 0);
signal Y_14_c4, Y_14_c5, Y_14_c6, Y_14_c7, Y_14_c8, Y_14_c9, Y_14_c10, Y_14_c11, Y_14_c12, Y_14_c13, Y_14_c14, Y_14_c15, Y_14_c16, Y_14_c17, Y_14_c18, Y_14_c19, Y_14_c20 :  std_logic_vector(3 downto 0);
signal S_14_c20 :  std_logic_vector(3 downto 0);
signal R_14_c20, R_14_c21, R_14_c22, R_14_c23, R_14_c24, R_14_c25, R_14_c26, R_14_c27, R_14_c28, R_14_c29, R_14_c30, R_14_c31, R_14_c32, R_14_c33 :  std_logic_vector(2 downto 0);
signal Cin_15_c20, Cin_15_c21 :  std_logic;
signal X_15_c4, X_15_c5, X_15_c6, X_15_c7, X_15_c8, X_15_c9, X_15_c10, X_15_c11, X_15_c12, X_15_c13, X_15_c14, X_15_c15, X_15_c16, X_15_c17, X_15_c18, X_15_c19, X_15_c20, X_15_c21 :  std_logic_vector(3 downto 0);
signal Y_15_c4, Y_15_c5, Y_15_c6, Y_15_c7, Y_15_c8, Y_15_c9, Y_15_c10, Y_15_c11, Y_15_c12, Y_15_c13, Y_15_c14, Y_15_c15, Y_15_c16, Y_15_c17, Y_15_c18, Y_15_c19, Y_15_c20, Y_15_c21 :  std_logic_vector(3 downto 0);
signal S_15_c21 :  std_logic_vector(3 downto 0);
signal R_15_c21, R_15_c22, R_15_c23, R_15_c24, R_15_c25, R_15_c26, R_15_c27, R_15_c28, R_15_c29, R_15_c30, R_15_c31, R_15_c32, R_15_c33 :  std_logic_vector(2 downto 0);
signal Cin_16_c21, Cin_16_c22 :  std_logic;
signal X_16_c4, X_16_c5, X_16_c6, X_16_c7, X_16_c8, X_16_c9, X_16_c10, X_16_c11, X_16_c12, X_16_c13, X_16_c14, X_16_c15, X_16_c16, X_16_c17, X_16_c18, X_16_c19, X_16_c20, X_16_c21, X_16_c22 :  std_logic_vector(3 downto 0);
signal Y_16_c4, Y_16_c5, Y_16_c6, Y_16_c7, Y_16_c8, Y_16_c9, Y_16_c10, Y_16_c11, Y_16_c12, Y_16_c13, Y_16_c14, Y_16_c15, Y_16_c16, Y_16_c17, Y_16_c18, Y_16_c19, Y_16_c20, Y_16_c21, Y_16_c22 :  std_logic_vector(3 downto 0);
signal S_16_c22 :  std_logic_vector(3 downto 0);
signal R_16_c22, R_16_c23, R_16_c24, R_16_c25, R_16_c26, R_16_c27, R_16_c28, R_16_c29, R_16_c30, R_16_c31, R_16_c32, R_16_c33 :  std_logic_vector(2 downto 0);
signal Cin_17_c22, Cin_17_c23 :  std_logic;
signal X_17_c4, X_17_c5, X_17_c6, X_17_c7, X_17_c8, X_17_c9, X_17_c10, X_17_c11, X_17_c12, X_17_c13, X_17_c14, X_17_c15, X_17_c16, X_17_c17, X_17_c18, X_17_c19, X_17_c20, X_17_c21, X_17_c22, X_17_c23 :  std_logic_vector(3 downto 0);
signal Y_17_c4, Y_17_c5, Y_17_c6, Y_17_c7, Y_17_c8, Y_17_c9, Y_17_c10, Y_17_c11, Y_17_c12, Y_17_c13, Y_17_c14, Y_17_c15, Y_17_c16, Y_17_c17, Y_17_c18, Y_17_c19, Y_17_c20, Y_17_c21, Y_17_c22, Y_17_c23 :  std_logic_vector(3 downto 0);
signal S_17_c23 :  std_logic_vector(3 downto 0);
signal R_17_c23, R_17_c24, R_17_c25, R_17_c26, R_17_c27, R_17_c28, R_17_c29, R_17_c30, R_17_c31, R_17_c32, R_17_c33 :  std_logic_vector(2 downto 0);
signal Cin_18_c23, Cin_18_c24 :  std_logic;
signal X_18_c4, X_18_c5, X_18_c6, X_18_c7, X_18_c8, X_18_c9, X_18_c10, X_18_c11, X_18_c12, X_18_c13, X_18_c14, X_18_c15, X_18_c16, X_18_c17, X_18_c18, X_18_c19, X_18_c20, X_18_c21, X_18_c22, X_18_c23, X_18_c24 :  std_logic_vector(3 downto 0);
signal Y_18_c4, Y_18_c5, Y_18_c6, Y_18_c7, Y_18_c8, Y_18_c9, Y_18_c10, Y_18_c11, Y_18_c12, Y_18_c13, Y_18_c14, Y_18_c15, Y_18_c16, Y_18_c17, Y_18_c18, Y_18_c19, Y_18_c20, Y_18_c21, Y_18_c22, Y_18_c23, Y_18_c24 :  std_logic_vector(3 downto 0);
signal S_18_c24 :  std_logic_vector(3 downto 0);
signal R_18_c24, R_18_c25, R_18_c26, R_18_c27, R_18_c28, R_18_c29, R_18_c30, R_18_c31, R_18_c32, R_18_c33 :  std_logic_vector(2 downto 0);
signal Cin_19_c24, Cin_19_c25 :  std_logic;
signal X_19_c4, X_19_c5, X_19_c6, X_19_c7, X_19_c8, X_19_c9, X_19_c10, X_19_c11, X_19_c12, X_19_c13, X_19_c14, X_19_c15, X_19_c16, X_19_c17, X_19_c18, X_19_c19, X_19_c20, X_19_c21, X_19_c22, X_19_c23, X_19_c24, X_19_c25 :  std_logic_vector(3 downto 0);
signal Y_19_c4, Y_19_c5, Y_19_c6, Y_19_c7, Y_19_c8, Y_19_c9, Y_19_c10, Y_19_c11, Y_19_c12, Y_19_c13, Y_19_c14, Y_19_c15, Y_19_c16, Y_19_c17, Y_19_c18, Y_19_c19, Y_19_c20, Y_19_c21, Y_19_c22, Y_19_c23, Y_19_c24, Y_19_c25 :  std_logic_vector(3 downto 0);
signal S_19_c25 :  std_logic_vector(3 downto 0);
signal R_19_c25, R_19_c26, R_19_c27, R_19_c28, R_19_c29, R_19_c30, R_19_c31, R_19_c32, R_19_c33 :  std_logic_vector(2 downto 0);
signal Cin_20_c25, Cin_20_c26 :  std_logic;
signal X_20_c4, X_20_c5, X_20_c6, X_20_c7, X_20_c8, X_20_c9, X_20_c10, X_20_c11, X_20_c12, X_20_c13, X_20_c14, X_20_c15, X_20_c16, X_20_c17, X_20_c18, X_20_c19, X_20_c20, X_20_c21, X_20_c22, X_20_c23, X_20_c24, X_20_c25, X_20_c26 :  std_logic_vector(3 downto 0);
signal Y_20_c4, Y_20_c5, Y_20_c6, Y_20_c7, Y_20_c8, Y_20_c9, Y_20_c10, Y_20_c11, Y_20_c12, Y_20_c13, Y_20_c14, Y_20_c15, Y_20_c16, Y_20_c17, Y_20_c18, Y_20_c19, Y_20_c20, Y_20_c21, Y_20_c22, Y_20_c23, Y_20_c24, Y_20_c25, Y_20_c26 :  std_logic_vector(3 downto 0);
signal S_20_c26 :  std_logic_vector(3 downto 0);
signal R_20_c26, R_20_c27, R_20_c28, R_20_c29, R_20_c30, R_20_c31, R_20_c32, R_20_c33 :  std_logic_vector(2 downto 0);
signal Cin_21_c26, Cin_21_c27 :  std_logic;
signal X_21_c4, X_21_c5, X_21_c6, X_21_c7, X_21_c8, X_21_c9, X_21_c10, X_21_c11, X_21_c12, X_21_c13, X_21_c14, X_21_c15, X_21_c16, X_21_c17, X_21_c18, X_21_c19, X_21_c20, X_21_c21, X_21_c22, X_21_c23, X_21_c24, X_21_c25, X_21_c26, X_21_c27 :  std_logic_vector(3 downto 0);
signal Y_21_c4, Y_21_c5, Y_21_c6, Y_21_c7, Y_21_c8, Y_21_c9, Y_21_c10, Y_21_c11, Y_21_c12, Y_21_c13, Y_21_c14, Y_21_c15, Y_21_c16, Y_21_c17, Y_21_c18, Y_21_c19, Y_21_c20, Y_21_c21, Y_21_c22, Y_21_c23, Y_21_c24, Y_21_c25, Y_21_c26, Y_21_c27 :  std_logic_vector(3 downto 0);
signal S_21_c27 :  std_logic_vector(3 downto 0);
signal R_21_c27, R_21_c28, R_21_c29, R_21_c30, R_21_c31, R_21_c32, R_21_c33 :  std_logic_vector(2 downto 0);
signal Cin_22_c27, Cin_22_c28 :  std_logic;
signal X_22_c4, X_22_c5, X_22_c6, X_22_c7, X_22_c8, X_22_c9, X_22_c10, X_22_c11, X_22_c12, X_22_c13, X_22_c14, X_22_c15, X_22_c16, X_22_c17, X_22_c18, X_22_c19, X_22_c20, X_22_c21, X_22_c22, X_22_c23, X_22_c24, X_22_c25, X_22_c26, X_22_c27, X_22_c28 :  std_logic_vector(3 downto 0);
signal Y_22_c4, Y_22_c5, Y_22_c6, Y_22_c7, Y_22_c8, Y_22_c9, Y_22_c10, Y_22_c11, Y_22_c12, Y_22_c13, Y_22_c14, Y_22_c15, Y_22_c16, Y_22_c17, Y_22_c18, Y_22_c19, Y_22_c20, Y_22_c21, Y_22_c22, Y_22_c23, Y_22_c24, Y_22_c25, Y_22_c26, Y_22_c27, Y_22_c28 :  std_logic_vector(3 downto 0);
signal S_22_c28 :  std_logic_vector(3 downto 0);
signal R_22_c28, R_22_c29, R_22_c30, R_22_c31, R_22_c32, R_22_c33 :  std_logic_vector(2 downto 0);
signal Cin_23_c28, Cin_23_c29 :  std_logic;
signal X_23_c4, X_23_c5, X_23_c6, X_23_c7, X_23_c8, X_23_c9, X_23_c10, X_23_c11, X_23_c12, X_23_c13, X_23_c14, X_23_c15, X_23_c16, X_23_c17, X_23_c18, X_23_c19, X_23_c20, X_23_c21, X_23_c22, X_23_c23, X_23_c24, X_23_c25, X_23_c26, X_23_c27, X_23_c28, X_23_c29 :  std_logic_vector(3 downto 0);
signal Y_23_c4, Y_23_c5, Y_23_c6, Y_23_c7, Y_23_c8, Y_23_c9, Y_23_c10, Y_23_c11, Y_23_c12, Y_23_c13, Y_23_c14, Y_23_c15, Y_23_c16, Y_23_c17, Y_23_c18, Y_23_c19, Y_23_c20, Y_23_c21, Y_23_c22, Y_23_c23, Y_23_c24, Y_23_c25, Y_23_c26, Y_23_c27, Y_23_c28, Y_23_c29 :  std_logic_vector(3 downto 0);
signal S_23_c29 :  std_logic_vector(3 downto 0);
signal R_23_c29, R_23_c30, R_23_c31, R_23_c32, R_23_c33 :  std_logic_vector(2 downto 0);
signal Cin_24_c29, Cin_24_c30 :  std_logic;
signal X_24_c4, X_24_c5, X_24_c6, X_24_c7, X_24_c8, X_24_c9, X_24_c10, X_24_c11, X_24_c12, X_24_c13, X_24_c14, X_24_c15, X_24_c16, X_24_c17, X_24_c18, X_24_c19, X_24_c20, X_24_c21, X_24_c22, X_24_c23, X_24_c24, X_24_c25, X_24_c26, X_24_c27, X_24_c28, X_24_c29, X_24_c30 :  std_logic_vector(3 downto 0);
signal Y_24_c4, Y_24_c5, Y_24_c6, Y_24_c7, Y_24_c8, Y_24_c9, Y_24_c10, Y_24_c11, Y_24_c12, Y_24_c13, Y_24_c14, Y_24_c15, Y_24_c16, Y_24_c17, Y_24_c18, Y_24_c19, Y_24_c20, Y_24_c21, Y_24_c22, Y_24_c23, Y_24_c24, Y_24_c25, Y_24_c26, Y_24_c27, Y_24_c28, Y_24_c29, Y_24_c30 :  std_logic_vector(3 downto 0);
signal S_24_c30 :  std_logic_vector(3 downto 0);
signal R_24_c30, R_24_c31, R_24_c32, R_24_c33 :  std_logic_vector(2 downto 0);
signal Cin_25_c30, Cin_25_c31 :  std_logic;
signal X_25_c4, X_25_c5, X_25_c6, X_25_c7, X_25_c8, X_25_c9, X_25_c10, X_25_c11, X_25_c12, X_25_c13, X_25_c14, X_25_c15, X_25_c16, X_25_c17, X_25_c18, X_25_c19, X_25_c20, X_25_c21, X_25_c22, X_25_c23, X_25_c24, X_25_c25, X_25_c26, X_25_c27, X_25_c28, X_25_c29, X_25_c30, X_25_c31 :  std_logic_vector(3 downto 0);
signal Y_25_c4, Y_25_c5, Y_25_c6, Y_25_c7, Y_25_c8, Y_25_c9, Y_25_c10, Y_25_c11, Y_25_c12, Y_25_c13, Y_25_c14, Y_25_c15, Y_25_c16, Y_25_c17, Y_25_c18, Y_25_c19, Y_25_c20, Y_25_c21, Y_25_c22, Y_25_c23, Y_25_c24, Y_25_c25, Y_25_c26, Y_25_c27, Y_25_c28, Y_25_c29, Y_25_c30, Y_25_c31 :  std_logic_vector(3 downto 0);
signal S_25_c31 :  std_logic_vector(3 downto 0);
signal R_25_c31, R_25_c32, R_25_c33 :  std_logic_vector(2 downto 0);
signal Cin_26_c31, Cin_26_c32 :  std_logic;
signal X_26_c4, X_26_c5, X_26_c6, X_26_c7, X_26_c8, X_26_c9, X_26_c10, X_26_c11, X_26_c12, X_26_c13, X_26_c14, X_26_c15, X_26_c16, X_26_c17, X_26_c18, X_26_c19, X_26_c20, X_26_c21, X_26_c22, X_26_c23, X_26_c24, X_26_c25, X_26_c26, X_26_c27, X_26_c28, X_26_c29, X_26_c30, X_26_c31, X_26_c32 :  std_logic_vector(3 downto 0);
signal Y_26_c4, Y_26_c5, Y_26_c6, Y_26_c7, Y_26_c8, Y_26_c9, Y_26_c10, Y_26_c11, Y_26_c12, Y_26_c13, Y_26_c14, Y_26_c15, Y_26_c16, Y_26_c17, Y_26_c18, Y_26_c19, Y_26_c20, Y_26_c21, Y_26_c22, Y_26_c23, Y_26_c24, Y_26_c25, Y_26_c26, Y_26_c27, Y_26_c28, Y_26_c29, Y_26_c30, Y_26_c31, Y_26_c32 :  std_logic_vector(3 downto 0);
signal S_26_c32 :  std_logic_vector(3 downto 0);
signal R_26_c32, R_26_c33 :  std_logic_vector(2 downto 0);
signal Cin_27_c32, Cin_27_c33 :  std_logic;
signal X_27_c4, X_27_c5, X_27_c6, X_27_c7, X_27_c8, X_27_c9, X_27_c10, X_27_c11, X_27_c12, X_27_c13, X_27_c14, X_27_c15, X_27_c16, X_27_c17, X_27_c18, X_27_c19, X_27_c20, X_27_c21, X_27_c22, X_27_c23, X_27_c24, X_27_c25, X_27_c26, X_27_c27, X_27_c28, X_27_c29, X_27_c30, X_27_c31, X_27_c32, X_27_c33 :  std_logic_vector(3 downto 0);
signal Y_27_c4, Y_27_c5, Y_27_c6, Y_27_c7, Y_27_c8, Y_27_c9, Y_27_c10, Y_27_c11, Y_27_c12, Y_27_c13, Y_27_c14, Y_27_c15, Y_27_c16, Y_27_c17, Y_27_c18, Y_27_c19, Y_27_c20, Y_27_c21, Y_27_c22, Y_27_c23, Y_27_c24, Y_27_c25, Y_27_c26, Y_27_c27, Y_27_c28, Y_27_c29, Y_27_c30, Y_27_c31, Y_27_c32, Y_27_c33 :  std_logic_vector(3 downto 0);
signal S_27_c33 :  std_logic_vector(3 downto 0);
signal R_27_c33 :  std_logic_vector(2 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
            end if;
            if ce_4 = '1' then
               Cin_0_c4 <= Cin_0_c3;
            end if;
            if ce_5 = '1' then
               Cin_0_c5 <= Cin_0_c4;
               X_0_c5 <= X_0_c4;
               Y_0_c5 <= Y_0_c4;
               X_1_c5 <= X_1_c4;
               Y_1_c5 <= Y_1_c4;
               X_2_c5 <= X_2_c4;
               Y_2_c5 <= Y_2_c4;
               X_3_c5 <= X_3_c4;
               Y_3_c5 <= Y_3_c4;
               X_4_c5 <= X_4_c4;
               Y_4_c5 <= Y_4_c4;
               X_5_c5 <= X_5_c4;
               Y_5_c5 <= Y_5_c4;
               X_6_c5 <= X_6_c4;
               Y_6_c5 <= Y_6_c4;
               X_7_c5 <= X_7_c4;
               Y_7_c5 <= Y_7_c4;
               X_8_c5 <= X_8_c4;
               Y_8_c5 <= Y_8_c4;
               X_9_c5 <= X_9_c4;
               Y_9_c5 <= Y_9_c4;
               X_10_c5 <= X_10_c4;
               Y_10_c5 <= Y_10_c4;
               X_11_c5 <= X_11_c4;
               Y_11_c5 <= Y_11_c4;
               X_12_c5 <= X_12_c4;
               Y_12_c5 <= Y_12_c4;
               X_13_c5 <= X_13_c4;
               Y_13_c5 <= Y_13_c4;
               X_14_c5 <= X_14_c4;
               Y_14_c5 <= Y_14_c4;
               X_15_c5 <= X_15_c4;
               Y_15_c5 <= Y_15_c4;
               X_16_c5 <= X_16_c4;
               Y_16_c5 <= Y_16_c4;
               X_17_c5 <= X_17_c4;
               Y_17_c5 <= Y_17_c4;
               X_18_c5 <= X_18_c4;
               Y_18_c5 <= Y_18_c4;
               X_19_c5 <= X_19_c4;
               Y_19_c5 <= Y_19_c4;
               X_20_c5 <= X_20_c4;
               Y_20_c5 <= Y_20_c4;
               X_21_c5 <= X_21_c4;
               Y_21_c5 <= Y_21_c4;
               X_22_c5 <= X_22_c4;
               Y_22_c5 <= Y_22_c4;
               X_23_c5 <= X_23_c4;
               Y_23_c5 <= Y_23_c4;
               X_24_c5 <= X_24_c4;
               Y_24_c5 <= Y_24_c4;
               X_25_c5 <= X_25_c4;
               Y_25_c5 <= Y_25_c4;
               X_26_c5 <= X_26_c4;
               Y_26_c5 <= Y_26_c4;
               X_27_c5 <= X_27_c4;
               Y_27_c5 <= Y_27_c4;
            end if;
            if ce_6 = '1' then
               R_0_c6 <= R_0_c5;
               Cin_1_c6 <= Cin_1_c5;
               X_1_c6 <= X_1_c5;
               Y_1_c6 <= Y_1_c5;
               X_2_c6 <= X_2_c5;
               Y_2_c6 <= Y_2_c5;
               X_3_c6 <= X_3_c5;
               Y_3_c6 <= Y_3_c5;
               X_4_c6 <= X_4_c5;
               Y_4_c6 <= Y_4_c5;
               X_5_c6 <= X_5_c5;
               Y_5_c6 <= Y_5_c5;
               X_6_c6 <= X_6_c5;
               Y_6_c6 <= Y_6_c5;
               X_7_c6 <= X_7_c5;
               Y_7_c6 <= Y_7_c5;
               X_8_c6 <= X_8_c5;
               Y_8_c6 <= Y_8_c5;
               X_9_c6 <= X_9_c5;
               Y_9_c6 <= Y_9_c5;
               X_10_c6 <= X_10_c5;
               Y_10_c6 <= Y_10_c5;
               X_11_c6 <= X_11_c5;
               Y_11_c6 <= Y_11_c5;
               X_12_c6 <= X_12_c5;
               Y_12_c6 <= Y_12_c5;
               X_13_c6 <= X_13_c5;
               Y_13_c6 <= Y_13_c5;
               X_14_c6 <= X_14_c5;
               Y_14_c6 <= Y_14_c5;
               X_15_c6 <= X_15_c5;
               Y_15_c6 <= Y_15_c5;
               X_16_c6 <= X_16_c5;
               Y_16_c6 <= Y_16_c5;
               X_17_c6 <= X_17_c5;
               Y_17_c6 <= Y_17_c5;
               X_18_c6 <= X_18_c5;
               Y_18_c6 <= Y_18_c5;
               X_19_c6 <= X_19_c5;
               Y_19_c6 <= Y_19_c5;
               X_20_c6 <= X_20_c5;
               Y_20_c6 <= Y_20_c5;
               X_21_c6 <= X_21_c5;
               Y_21_c6 <= Y_21_c5;
               X_22_c6 <= X_22_c5;
               Y_22_c6 <= Y_22_c5;
               X_23_c6 <= X_23_c5;
               Y_23_c6 <= Y_23_c5;
               X_24_c6 <= X_24_c5;
               Y_24_c6 <= Y_24_c5;
               X_25_c6 <= X_25_c5;
               Y_25_c6 <= Y_25_c5;
               X_26_c6 <= X_26_c5;
               Y_26_c6 <= Y_26_c5;
               X_27_c6 <= X_27_c5;
               Y_27_c6 <= Y_27_c5;
            end if;
            if ce_7 = '1' then
               R_0_c7 <= R_0_c6;
               R_1_c7 <= R_1_c6;
               Cin_2_c7 <= Cin_2_c6;
               X_2_c7 <= X_2_c6;
               Y_2_c7 <= Y_2_c6;
               X_3_c7 <= X_3_c6;
               Y_3_c7 <= Y_3_c6;
               X_4_c7 <= X_4_c6;
               Y_4_c7 <= Y_4_c6;
               X_5_c7 <= X_5_c6;
               Y_5_c7 <= Y_5_c6;
               X_6_c7 <= X_6_c6;
               Y_6_c7 <= Y_6_c6;
               X_7_c7 <= X_7_c6;
               Y_7_c7 <= Y_7_c6;
               X_8_c7 <= X_8_c6;
               Y_8_c7 <= Y_8_c6;
               X_9_c7 <= X_9_c6;
               Y_9_c7 <= Y_9_c6;
               X_10_c7 <= X_10_c6;
               Y_10_c7 <= Y_10_c6;
               X_11_c7 <= X_11_c6;
               Y_11_c7 <= Y_11_c6;
               X_12_c7 <= X_12_c6;
               Y_12_c7 <= Y_12_c6;
               X_13_c7 <= X_13_c6;
               Y_13_c7 <= Y_13_c6;
               X_14_c7 <= X_14_c6;
               Y_14_c7 <= Y_14_c6;
               X_15_c7 <= X_15_c6;
               Y_15_c7 <= Y_15_c6;
               X_16_c7 <= X_16_c6;
               Y_16_c7 <= Y_16_c6;
               X_17_c7 <= X_17_c6;
               Y_17_c7 <= Y_17_c6;
               X_18_c7 <= X_18_c6;
               Y_18_c7 <= Y_18_c6;
               X_19_c7 <= X_19_c6;
               Y_19_c7 <= Y_19_c6;
               X_20_c7 <= X_20_c6;
               Y_20_c7 <= Y_20_c6;
               X_21_c7 <= X_21_c6;
               Y_21_c7 <= Y_21_c6;
               X_22_c7 <= X_22_c6;
               Y_22_c7 <= Y_22_c6;
               X_23_c7 <= X_23_c6;
               Y_23_c7 <= Y_23_c6;
               X_24_c7 <= X_24_c6;
               Y_24_c7 <= Y_24_c6;
               X_25_c7 <= X_25_c6;
               Y_25_c7 <= Y_25_c6;
               X_26_c7 <= X_26_c6;
               Y_26_c7 <= Y_26_c6;
               X_27_c7 <= X_27_c6;
               Y_27_c7 <= Y_27_c6;
            end if;
            if ce_8 = '1' then
               R_0_c8 <= R_0_c7;
               R_1_c8 <= R_1_c7;
               R_2_c8 <= R_2_c7;
               Cin_3_c8 <= Cin_3_c7;
               X_3_c8 <= X_3_c7;
               Y_3_c8 <= Y_3_c7;
               X_4_c8 <= X_4_c7;
               Y_4_c8 <= Y_4_c7;
               X_5_c8 <= X_5_c7;
               Y_5_c8 <= Y_5_c7;
               X_6_c8 <= X_6_c7;
               Y_6_c8 <= Y_6_c7;
               X_7_c8 <= X_7_c7;
               Y_7_c8 <= Y_7_c7;
               X_8_c8 <= X_8_c7;
               Y_8_c8 <= Y_8_c7;
               X_9_c8 <= X_9_c7;
               Y_9_c8 <= Y_9_c7;
               X_10_c8 <= X_10_c7;
               Y_10_c8 <= Y_10_c7;
               X_11_c8 <= X_11_c7;
               Y_11_c8 <= Y_11_c7;
               X_12_c8 <= X_12_c7;
               Y_12_c8 <= Y_12_c7;
               X_13_c8 <= X_13_c7;
               Y_13_c8 <= Y_13_c7;
               X_14_c8 <= X_14_c7;
               Y_14_c8 <= Y_14_c7;
               X_15_c8 <= X_15_c7;
               Y_15_c8 <= Y_15_c7;
               X_16_c8 <= X_16_c7;
               Y_16_c8 <= Y_16_c7;
               X_17_c8 <= X_17_c7;
               Y_17_c8 <= Y_17_c7;
               X_18_c8 <= X_18_c7;
               Y_18_c8 <= Y_18_c7;
               X_19_c8 <= X_19_c7;
               Y_19_c8 <= Y_19_c7;
               X_20_c8 <= X_20_c7;
               Y_20_c8 <= Y_20_c7;
               X_21_c8 <= X_21_c7;
               Y_21_c8 <= Y_21_c7;
               X_22_c8 <= X_22_c7;
               Y_22_c8 <= Y_22_c7;
               X_23_c8 <= X_23_c7;
               Y_23_c8 <= Y_23_c7;
               X_24_c8 <= X_24_c7;
               Y_24_c8 <= Y_24_c7;
               X_25_c8 <= X_25_c7;
               Y_25_c8 <= Y_25_c7;
               X_26_c8 <= X_26_c7;
               Y_26_c8 <= Y_26_c7;
               X_27_c8 <= X_27_c7;
               Y_27_c8 <= Y_27_c7;
            end if;
            if ce_9 = '1' then
               R_0_c9 <= R_0_c8;
               R_1_c9 <= R_1_c8;
               R_2_c9 <= R_2_c8;
               R_3_c9 <= R_3_c8;
               Cin_4_c9 <= Cin_4_c8;
               X_4_c9 <= X_4_c8;
               Y_4_c9 <= Y_4_c8;
               X_5_c9 <= X_5_c8;
               Y_5_c9 <= Y_5_c8;
               X_6_c9 <= X_6_c8;
               Y_6_c9 <= Y_6_c8;
               X_7_c9 <= X_7_c8;
               Y_7_c9 <= Y_7_c8;
               X_8_c9 <= X_8_c8;
               Y_8_c9 <= Y_8_c8;
               X_9_c9 <= X_9_c8;
               Y_9_c9 <= Y_9_c8;
               X_10_c9 <= X_10_c8;
               Y_10_c9 <= Y_10_c8;
               X_11_c9 <= X_11_c8;
               Y_11_c9 <= Y_11_c8;
               X_12_c9 <= X_12_c8;
               Y_12_c9 <= Y_12_c8;
               X_13_c9 <= X_13_c8;
               Y_13_c9 <= Y_13_c8;
               X_14_c9 <= X_14_c8;
               Y_14_c9 <= Y_14_c8;
               X_15_c9 <= X_15_c8;
               Y_15_c9 <= Y_15_c8;
               X_16_c9 <= X_16_c8;
               Y_16_c9 <= Y_16_c8;
               X_17_c9 <= X_17_c8;
               Y_17_c9 <= Y_17_c8;
               X_18_c9 <= X_18_c8;
               Y_18_c9 <= Y_18_c8;
               X_19_c9 <= X_19_c8;
               Y_19_c9 <= Y_19_c8;
               X_20_c9 <= X_20_c8;
               Y_20_c9 <= Y_20_c8;
               X_21_c9 <= X_21_c8;
               Y_21_c9 <= Y_21_c8;
               X_22_c9 <= X_22_c8;
               Y_22_c9 <= Y_22_c8;
               X_23_c9 <= X_23_c8;
               Y_23_c9 <= Y_23_c8;
               X_24_c9 <= X_24_c8;
               Y_24_c9 <= Y_24_c8;
               X_25_c9 <= X_25_c8;
               Y_25_c9 <= Y_25_c8;
               X_26_c9 <= X_26_c8;
               Y_26_c9 <= Y_26_c8;
               X_27_c9 <= X_27_c8;
               Y_27_c9 <= Y_27_c8;
            end if;
            if ce_10 = '1' then
               R_0_c10 <= R_0_c9;
               R_1_c10 <= R_1_c9;
               R_2_c10 <= R_2_c9;
               R_3_c10 <= R_3_c9;
               R_4_c10 <= R_4_c9;
               Cin_5_c10 <= Cin_5_c9;
               X_5_c10 <= X_5_c9;
               Y_5_c10 <= Y_5_c9;
               X_6_c10 <= X_6_c9;
               Y_6_c10 <= Y_6_c9;
               X_7_c10 <= X_7_c9;
               Y_7_c10 <= Y_7_c9;
               X_8_c10 <= X_8_c9;
               Y_8_c10 <= Y_8_c9;
               X_9_c10 <= X_9_c9;
               Y_9_c10 <= Y_9_c9;
               X_10_c10 <= X_10_c9;
               Y_10_c10 <= Y_10_c9;
               X_11_c10 <= X_11_c9;
               Y_11_c10 <= Y_11_c9;
               X_12_c10 <= X_12_c9;
               Y_12_c10 <= Y_12_c9;
               X_13_c10 <= X_13_c9;
               Y_13_c10 <= Y_13_c9;
               X_14_c10 <= X_14_c9;
               Y_14_c10 <= Y_14_c9;
               X_15_c10 <= X_15_c9;
               Y_15_c10 <= Y_15_c9;
               X_16_c10 <= X_16_c9;
               Y_16_c10 <= Y_16_c9;
               X_17_c10 <= X_17_c9;
               Y_17_c10 <= Y_17_c9;
               X_18_c10 <= X_18_c9;
               Y_18_c10 <= Y_18_c9;
               X_19_c10 <= X_19_c9;
               Y_19_c10 <= Y_19_c9;
               X_20_c10 <= X_20_c9;
               Y_20_c10 <= Y_20_c9;
               X_21_c10 <= X_21_c9;
               Y_21_c10 <= Y_21_c9;
               X_22_c10 <= X_22_c9;
               Y_22_c10 <= Y_22_c9;
               X_23_c10 <= X_23_c9;
               Y_23_c10 <= Y_23_c9;
               X_24_c10 <= X_24_c9;
               Y_24_c10 <= Y_24_c9;
               X_25_c10 <= X_25_c9;
               Y_25_c10 <= Y_25_c9;
               X_26_c10 <= X_26_c9;
               Y_26_c10 <= Y_26_c9;
               X_27_c10 <= X_27_c9;
               Y_27_c10 <= Y_27_c9;
            end if;
            if ce_11 = '1' then
               R_0_c11 <= R_0_c10;
               R_1_c11 <= R_1_c10;
               R_2_c11 <= R_2_c10;
               R_3_c11 <= R_3_c10;
               R_4_c11 <= R_4_c10;
               R_5_c11 <= R_5_c10;
               Cin_6_c11 <= Cin_6_c10;
               X_6_c11 <= X_6_c10;
               Y_6_c11 <= Y_6_c10;
               X_7_c11 <= X_7_c10;
               Y_7_c11 <= Y_7_c10;
               X_8_c11 <= X_8_c10;
               Y_8_c11 <= Y_8_c10;
               X_9_c11 <= X_9_c10;
               Y_9_c11 <= Y_9_c10;
               X_10_c11 <= X_10_c10;
               Y_10_c11 <= Y_10_c10;
               X_11_c11 <= X_11_c10;
               Y_11_c11 <= Y_11_c10;
               X_12_c11 <= X_12_c10;
               Y_12_c11 <= Y_12_c10;
               X_13_c11 <= X_13_c10;
               Y_13_c11 <= Y_13_c10;
               X_14_c11 <= X_14_c10;
               Y_14_c11 <= Y_14_c10;
               X_15_c11 <= X_15_c10;
               Y_15_c11 <= Y_15_c10;
               X_16_c11 <= X_16_c10;
               Y_16_c11 <= Y_16_c10;
               X_17_c11 <= X_17_c10;
               Y_17_c11 <= Y_17_c10;
               X_18_c11 <= X_18_c10;
               Y_18_c11 <= Y_18_c10;
               X_19_c11 <= X_19_c10;
               Y_19_c11 <= Y_19_c10;
               X_20_c11 <= X_20_c10;
               Y_20_c11 <= Y_20_c10;
               X_21_c11 <= X_21_c10;
               Y_21_c11 <= Y_21_c10;
               X_22_c11 <= X_22_c10;
               Y_22_c11 <= Y_22_c10;
               X_23_c11 <= X_23_c10;
               Y_23_c11 <= Y_23_c10;
               X_24_c11 <= X_24_c10;
               Y_24_c11 <= Y_24_c10;
               X_25_c11 <= X_25_c10;
               Y_25_c11 <= Y_25_c10;
               X_26_c11 <= X_26_c10;
               Y_26_c11 <= Y_26_c10;
               X_27_c11 <= X_27_c10;
               Y_27_c11 <= Y_27_c10;
            end if;
            if ce_12 = '1' then
               R_0_c12 <= R_0_c11;
               R_1_c12 <= R_1_c11;
               R_2_c12 <= R_2_c11;
               R_3_c12 <= R_3_c11;
               R_4_c12 <= R_4_c11;
               R_5_c12 <= R_5_c11;
               R_6_c12 <= R_6_c11;
               Cin_7_c12 <= Cin_7_c11;
               X_7_c12 <= X_7_c11;
               Y_7_c12 <= Y_7_c11;
               X_8_c12 <= X_8_c11;
               Y_8_c12 <= Y_8_c11;
               X_9_c12 <= X_9_c11;
               Y_9_c12 <= Y_9_c11;
               X_10_c12 <= X_10_c11;
               Y_10_c12 <= Y_10_c11;
               X_11_c12 <= X_11_c11;
               Y_11_c12 <= Y_11_c11;
               X_12_c12 <= X_12_c11;
               Y_12_c12 <= Y_12_c11;
               X_13_c12 <= X_13_c11;
               Y_13_c12 <= Y_13_c11;
               X_14_c12 <= X_14_c11;
               Y_14_c12 <= Y_14_c11;
               X_15_c12 <= X_15_c11;
               Y_15_c12 <= Y_15_c11;
               X_16_c12 <= X_16_c11;
               Y_16_c12 <= Y_16_c11;
               X_17_c12 <= X_17_c11;
               Y_17_c12 <= Y_17_c11;
               X_18_c12 <= X_18_c11;
               Y_18_c12 <= Y_18_c11;
               X_19_c12 <= X_19_c11;
               Y_19_c12 <= Y_19_c11;
               X_20_c12 <= X_20_c11;
               Y_20_c12 <= Y_20_c11;
               X_21_c12 <= X_21_c11;
               Y_21_c12 <= Y_21_c11;
               X_22_c12 <= X_22_c11;
               Y_22_c12 <= Y_22_c11;
               X_23_c12 <= X_23_c11;
               Y_23_c12 <= Y_23_c11;
               X_24_c12 <= X_24_c11;
               Y_24_c12 <= Y_24_c11;
               X_25_c12 <= X_25_c11;
               Y_25_c12 <= Y_25_c11;
               X_26_c12 <= X_26_c11;
               Y_26_c12 <= Y_26_c11;
               X_27_c12 <= X_27_c11;
               Y_27_c12 <= Y_27_c11;
            end if;
            if ce_13 = '1' then
               R_0_c13 <= R_0_c12;
               R_1_c13 <= R_1_c12;
               R_2_c13 <= R_2_c12;
               R_3_c13 <= R_3_c12;
               R_4_c13 <= R_4_c12;
               R_5_c13 <= R_5_c12;
               R_6_c13 <= R_6_c12;
               R_7_c13 <= R_7_c12;
               Cin_8_c13 <= Cin_8_c12;
               X_8_c13 <= X_8_c12;
               Y_8_c13 <= Y_8_c12;
               X_9_c13 <= X_9_c12;
               Y_9_c13 <= Y_9_c12;
               X_10_c13 <= X_10_c12;
               Y_10_c13 <= Y_10_c12;
               X_11_c13 <= X_11_c12;
               Y_11_c13 <= Y_11_c12;
               X_12_c13 <= X_12_c12;
               Y_12_c13 <= Y_12_c12;
               X_13_c13 <= X_13_c12;
               Y_13_c13 <= Y_13_c12;
               X_14_c13 <= X_14_c12;
               Y_14_c13 <= Y_14_c12;
               X_15_c13 <= X_15_c12;
               Y_15_c13 <= Y_15_c12;
               X_16_c13 <= X_16_c12;
               Y_16_c13 <= Y_16_c12;
               X_17_c13 <= X_17_c12;
               Y_17_c13 <= Y_17_c12;
               X_18_c13 <= X_18_c12;
               Y_18_c13 <= Y_18_c12;
               X_19_c13 <= X_19_c12;
               Y_19_c13 <= Y_19_c12;
               X_20_c13 <= X_20_c12;
               Y_20_c13 <= Y_20_c12;
               X_21_c13 <= X_21_c12;
               Y_21_c13 <= Y_21_c12;
               X_22_c13 <= X_22_c12;
               Y_22_c13 <= Y_22_c12;
               X_23_c13 <= X_23_c12;
               Y_23_c13 <= Y_23_c12;
               X_24_c13 <= X_24_c12;
               Y_24_c13 <= Y_24_c12;
               X_25_c13 <= X_25_c12;
               Y_25_c13 <= Y_25_c12;
               X_26_c13 <= X_26_c12;
               Y_26_c13 <= Y_26_c12;
               X_27_c13 <= X_27_c12;
               Y_27_c13 <= Y_27_c12;
            end if;
            if ce_14 = '1' then
               R_0_c14 <= R_0_c13;
               R_1_c14 <= R_1_c13;
               R_2_c14 <= R_2_c13;
               R_3_c14 <= R_3_c13;
               R_4_c14 <= R_4_c13;
               R_5_c14 <= R_5_c13;
               R_6_c14 <= R_6_c13;
               R_7_c14 <= R_7_c13;
               R_8_c14 <= R_8_c13;
               Cin_9_c14 <= Cin_9_c13;
               X_9_c14 <= X_9_c13;
               Y_9_c14 <= Y_9_c13;
               X_10_c14 <= X_10_c13;
               Y_10_c14 <= Y_10_c13;
               X_11_c14 <= X_11_c13;
               Y_11_c14 <= Y_11_c13;
               X_12_c14 <= X_12_c13;
               Y_12_c14 <= Y_12_c13;
               X_13_c14 <= X_13_c13;
               Y_13_c14 <= Y_13_c13;
               X_14_c14 <= X_14_c13;
               Y_14_c14 <= Y_14_c13;
               X_15_c14 <= X_15_c13;
               Y_15_c14 <= Y_15_c13;
               X_16_c14 <= X_16_c13;
               Y_16_c14 <= Y_16_c13;
               X_17_c14 <= X_17_c13;
               Y_17_c14 <= Y_17_c13;
               X_18_c14 <= X_18_c13;
               Y_18_c14 <= Y_18_c13;
               X_19_c14 <= X_19_c13;
               Y_19_c14 <= Y_19_c13;
               X_20_c14 <= X_20_c13;
               Y_20_c14 <= Y_20_c13;
               X_21_c14 <= X_21_c13;
               Y_21_c14 <= Y_21_c13;
               X_22_c14 <= X_22_c13;
               Y_22_c14 <= Y_22_c13;
               X_23_c14 <= X_23_c13;
               Y_23_c14 <= Y_23_c13;
               X_24_c14 <= X_24_c13;
               Y_24_c14 <= Y_24_c13;
               X_25_c14 <= X_25_c13;
               Y_25_c14 <= Y_25_c13;
               X_26_c14 <= X_26_c13;
               Y_26_c14 <= Y_26_c13;
               X_27_c14 <= X_27_c13;
               Y_27_c14 <= Y_27_c13;
            end if;
            if ce_15 = '1' then
               R_0_c15 <= R_0_c14;
               R_1_c15 <= R_1_c14;
               R_2_c15 <= R_2_c14;
               R_3_c15 <= R_3_c14;
               R_4_c15 <= R_4_c14;
               R_5_c15 <= R_5_c14;
               R_6_c15 <= R_6_c14;
               R_7_c15 <= R_7_c14;
               R_8_c15 <= R_8_c14;
               R_9_c15 <= R_9_c14;
               Cin_10_c15 <= Cin_10_c14;
               X_10_c15 <= X_10_c14;
               Y_10_c15 <= Y_10_c14;
               X_11_c15 <= X_11_c14;
               Y_11_c15 <= Y_11_c14;
               X_12_c15 <= X_12_c14;
               Y_12_c15 <= Y_12_c14;
               X_13_c15 <= X_13_c14;
               Y_13_c15 <= Y_13_c14;
               X_14_c15 <= X_14_c14;
               Y_14_c15 <= Y_14_c14;
               X_15_c15 <= X_15_c14;
               Y_15_c15 <= Y_15_c14;
               X_16_c15 <= X_16_c14;
               Y_16_c15 <= Y_16_c14;
               X_17_c15 <= X_17_c14;
               Y_17_c15 <= Y_17_c14;
               X_18_c15 <= X_18_c14;
               Y_18_c15 <= Y_18_c14;
               X_19_c15 <= X_19_c14;
               Y_19_c15 <= Y_19_c14;
               X_20_c15 <= X_20_c14;
               Y_20_c15 <= Y_20_c14;
               X_21_c15 <= X_21_c14;
               Y_21_c15 <= Y_21_c14;
               X_22_c15 <= X_22_c14;
               Y_22_c15 <= Y_22_c14;
               X_23_c15 <= X_23_c14;
               Y_23_c15 <= Y_23_c14;
               X_24_c15 <= X_24_c14;
               Y_24_c15 <= Y_24_c14;
               X_25_c15 <= X_25_c14;
               Y_25_c15 <= Y_25_c14;
               X_26_c15 <= X_26_c14;
               Y_26_c15 <= Y_26_c14;
               X_27_c15 <= X_27_c14;
               Y_27_c15 <= Y_27_c14;
            end if;
            if ce_16 = '1' then
               R_0_c16 <= R_0_c15;
               R_1_c16 <= R_1_c15;
               R_2_c16 <= R_2_c15;
               R_3_c16 <= R_3_c15;
               R_4_c16 <= R_4_c15;
               R_5_c16 <= R_5_c15;
               R_6_c16 <= R_6_c15;
               R_7_c16 <= R_7_c15;
               R_8_c16 <= R_8_c15;
               R_9_c16 <= R_9_c15;
               R_10_c16 <= R_10_c15;
               Cin_11_c16 <= Cin_11_c15;
               X_11_c16 <= X_11_c15;
               Y_11_c16 <= Y_11_c15;
               X_12_c16 <= X_12_c15;
               Y_12_c16 <= Y_12_c15;
               X_13_c16 <= X_13_c15;
               Y_13_c16 <= Y_13_c15;
               X_14_c16 <= X_14_c15;
               Y_14_c16 <= Y_14_c15;
               X_15_c16 <= X_15_c15;
               Y_15_c16 <= Y_15_c15;
               X_16_c16 <= X_16_c15;
               Y_16_c16 <= Y_16_c15;
               X_17_c16 <= X_17_c15;
               Y_17_c16 <= Y_17_c15;
               X_18_c16 <= X_18_c15;
               Y_18_c16 <= Y_18_c15;
               X_19_c16 <= X_19_c15;
               Y_19_c16 <= Y_19_c15;
               X_20_c16 <= X_20_c15;
               Y_20_c16 <= Y_20_c15;
               X_21_c16 <= X_21_c15;
               Y_21_c16 <= Y_21_c15;
               X_22_c16 <= X_22_c15;
               Y_22_c16 <= Y_22_c15;
               X_23_c16 <= X_23_c15;
               Y_23_c16 <= Y_23_c15;
               X_24_c16 <= X_24_c15;
               Y_24_c16 <= Y_24_c15;
               X_25_c16 <= X_25_c15;
               Y_25_c16 <= Y_25_c15;
               X_26_c16 <= X_26_c15;
               Y_26_c16 <= Y_26_c15;
               X_27_c16 <= X_27_c15;
               Y_27_c16 <= Y_27_c15;
            end if;
            if ce_17 = '1' then
               R_0_c17 <= R_0_c16;
               R_1_c17 <= R_1_c16;
               R_2_c17 <= R_2_c16;
               R_3_c17 <= R_3_c16;
               R_4_c17 <= R_4_c16;
               R_5_c17 <= R_5_c16;
               R_6_c17 <= R_6_c16;
               R_7_c17 <= R_7_c16;
               R_8_c17 <= R_8_c16;
               R_9_c17 <= R_9_c16;
               R_10_c17 <= R_10_c16;
               R_11_c17 <= R_11_c16;
               Cin_12_c17 <= Cin_12_c16;
               X_12_c17 <= X_12_c16;
               Y_12_c17 <= Y_12_c16;
               X_13_c17 <= X_13_c16;
               Y_13_c17 <= Y_13_c16;
               X_14_c17 <= X_14_c16;
               Y_14_c17 <= Y_14_c16;
               X_15_c17 <= X_15_c16;
               Y_15_c17 <= Y_15_c16;
               X_16_c17 <= X_16_c16;
               Y_16_c17 <= Y_16_c16;
               X_17_c17 <= X_17_c16;
               Y_17_c17 <= Y_17_c16;
               X_18_c17 <= X_18_c16;
               Y_18_c17 <= Y_18_c16;
               X_19_c17 <= X_19_c16;
               Y_19_c17 <= Y_19_c16;
               X_20_c17 <= X_20_c16;
               Y_20_c17 <= Y_20_c16;
               X_21_c17 <= X_21_c16;
               Y_21_c17 <= Y_21_c16;
               X_22_c17 <= X_22_c16;
               Y_22_c17 <= Y_22_c16;
               X_23_c17 <= X_23_c16;
               Y_23_c17 <= Y_23_c16;
               X_24_c17 <= X_24_c16;
               Y_24_c17 <= Y_24_c16;
               X_25_c17 <= X_25_c16;
               Y_25_c17 <= Y_25_c16;
               X_26_c17 <= X_26_c16;
               Y_26_c17 <= Y_26_c16;
               X_27_c17 <= X_27_c16;
               Y_27_c17 <= Y_27_c16;
            end if;
            if ce_18 = '1' then
               R_0_c18 <= R_0_c17;
               R_1_c18 <= R_1_c17;
               R_2_c18 <= R_2_c17;
               R_3_c18 <= R_3_c17;
               R_4_c18 <= R_4_c17;
               R_5_c18 <= R_5_c17;
               R_6_c18 <= R_6_c17;
               R_7_c18 <= R_7_c17;
               R_8_c18 <= R_8_c17;
               R_9_c18 <= R_9_c17;
               R_10_c18 <= R_10_c17;
               R_11_c18 <= R_11_c17;
               R_12_c18 <= R_12_c17;
               Cin_13_c18 <= Cin_13_c17;
               X_13_c18 <= X_13_c17;
               Y_13_c18 <= Y_13_c17;
               X_14_c18 <= X_14_c17;
               Y_14_c18 <= Y_14_c17;
               X_15_c18 <= X_15_c17;
               Y_15_c18 <= Y_15_c17;
               X_16_c18 <= X_16_c17;
               Y_16_c18 <= Y_16_c17;
               X_17_c18 <= X_17_c17;
               Y_17_c18 <= Y_17_c17;
               X_18_c18 <= X_18_c17;
               Y_18_c18 <= Y_18_c17;
               X_19_c18 <= X_19_c17;
               Y_19_c18 <= Y_19_c17;
               X_20_c18 <= X_20_c17;
               Y_20_c18 <= Y_20_c17;
               X_21_c18 <= X_21_c17;
               Y_21_c18 <= Y_21_c17;
               X_22_c18 <= X_22_c17;
               Y_22_c18 <= Y_22_c17;
               X_23_c18 <= X_23_c17;
               Y_23_c18 <= Y_23_c17;
               X_24_c18 <= X_24_c17;
               Y_24_c18 <= Y_24_c17;
               X_25_c18 <= X_25_c17;
               Y_25_c18 <= Y_25_c17;
               X_26_c18 <= X_26_c17;
               Y_26_c18 <= Y_26_c17;
               X_27_c18 <= X_27_c17;
               Y_27_c18 <= Y_27_c17;
            end if;
            if ce_19 = '1' then
               R_0_c19 <= R_0_c18;
               R_1_c19 <= R_1_c18;
               R_2_c19 <= R_2_c18;
               R_3_c19 <= R_3_c18;
               R_4_c19 <= R_4_c18;
               R_5_c19 <= R_5_c18;
               R_6_c19 <= R_6_c18;
               R_7_c19 <= R_7_c18;
               R_8_c19 <= R_8_c18;
               R_9_c19 <= R_9_c18;
               R_10_c19 <= R_10_c18;
               R_11_c19 <= R_11_c18;
               R_12_c19 <= R_12_c18;
               R_13_c19 <= R_13_c18;
               Cin_14_c19 <= Cin_14_c18;
               X_14_c19 <= X_14_c18;
               Y_14_c19 <= Y_14_c18;
               X_15_c19 <= X_15_c18;
               Y_15_c19 <= Y_15_c18;
               X_16_c19 <= X_16_c18;
               Y_16_c19 <= Y_16_c18;
               X_17_c19 <= X_17_c18;
               Y_17_c19 <= Y_17_c18;
               X_18_c19 <= X_18_c18;
               Y_18_c19 <= Y_18_c18;
               X_19_c19 <= X_19_c18;
               Y_19_c19 <= Y_19_c18;
               X_20_c19 <= X_20_c18;
               Y_20_c19 <= Y_20_c18;
               X_21_c19 <= X_21_c18;
               Y_21_c19 <= Y_21_c18;
               X_22_c19 <= X_22_c18;
               Y_22_c19 <= Y_22_c18;
               X_23_c19 <= X_23_c18;
               Y_23_c19 <= Y_23_c18;
               X_24_c19 <= X_24_c18;
               Y_24_c19 <= Y_24_c18;
               X_25_c19 <= X_25_c18;
               Y_25_c19 <= Y_25_c18;
               X_26_c19 <= X_26_c18;
               Y_26_c19 <= Y_26_c18;
               X_27_c19 <= X_27_c18;
               Y_27_c19 <= Y_27_c18;
            end if;
            if ce_20 = '1' then
               R_0_c20 <= R_0_c19;
               R_1_c20 <= R_1_c19;
               R_2_c20 <= R_2_c19;
               R_3_c20 <= R_3_c19;
               R_4_c20 <= R_4_c19;
               R_5_c20 <= R_5_c19;
               R_6_c20 <= R_6_c19;
               R_7_c20 <= R_7_c19;
               R_8_c20 <= R_8_c19;
               R_9_c20 <= R_9_c19;
               R_10_c20 <= R_10_c19;
               R_11_c20 <= R_11_c19;
               R_12_c20 <= R_12_c19;
               R_13_c20 <= R_13_c19;
               Cin_14_c20 <= Cin_14_c19;
               X_14_c20 <= X_14_c19;
               Y_14_c20 <= Y_14_c19;
               X_15_c20 <= X_15_c19;
               Y_15_c20 <= Y_15_c19;
               X_16_c20 <= X_16_c19;
               Y_16_c20 <= Y_16_c19;
               X_17_c20 <= X_17_c19;
               Y_17_c20 <= Y_17_c19;
               X_18_c20 <= X_18_c19;
               Y_18_c20 <= Y_18_c19;
               X_19_c20 <= X_19_c19;
               Y_19_c20 <= Y_19_c19;
               X_20_c20 <= X_20_c19;
               Y_20_c20 <= Y_20_c19;
               X_21_c20 <= X_21_c19;
               Y_21_c20 <= Y_21_c19;
               X_22_c20 <= X_22_c19;
               Y_22_c20 <= Y_22_c19;
               X_23_c20 <= X_23_c19;
               Y_23_c20 <= Y_23_c19;
               X_24_c20 <= X_24_c19;
               Y_24_c20 <= Y_24_c19;
               X_25_c20 <= X_25_c19;
               Y_25_c20 <= Y_25_c19;
               X_26_c20 <= X_26_c19;
               Y_26_c20 <= Y_26_c19;
               X_27_c20 <= X_27_c19;
               Y_27_c20 <= Y_27_c19;
            end if;
            if ce_21 = '1' then
               R_0_c21 <= R_0_c20;
               R_1_c21 <= R_1_c20;
               R_2_c21 <= R_2_c20;
               R_3_c21 <= R_3_c20;
               R_4_c21 <= R_4_c20;
               R_5_c21 <= R_5_c20;
               R_6_c21 <= R_6_c20;
               R_7_c21 <= R_7_c20;
               R_8_c21 <= R_8_c20;
               R_9_c21 <= R_9_c20;
               R_10_c21 <= R_10_c20;
               R_11_c21 <= R_11_c20;
               R_12_c21 <= R_12_c20;
               R_13_c21 <= R_13_c20;
               R_14_c21 <= R_14_c20;
               Cin_15_c21 <= Cin_15_c20;
               X_15_c21 <= X_15_c20;
               Y_15_c21 <= Y_15_c20;
               X_16_c21 <= X_16_c20;
               Y_16_c21 <= Y_16_c20;
               X_17_c21 <= X_17_c20;
               Y_17_c21 <= Y_17_c20;
               X_18_c21 <= X_18_c20;
               Y_18_c21 <= Y_18_c20;
               X_19_c21 <= X_19_c20;
               Y_19_c21 <= Y_19_c20;
               X_20_c21 <= X_20_c20;
               Y_20_c21 <= Y_20_c20;
               X_21_c21 <= X_21_c20;
               Y_21_c21 <= Y_21_c20;
               X_22_c21 <= X_22_c20;
               Y_22_c21 <= Y_22_c20;
               X_23_c21 <= X_23_c20;
               Y_23_c21 <= Y_23_c20;
               X_24_c21 <= X_24_c20;
               Y_24_c21 <= Y_24_c20;
               X_25_c21 <= X_25_c20;
               Y_25_c21 <= Y_25_c20;
               X_26_c21 <= X_26_c20;
               Y_26_c21 <= Y_26_c20;
               X_27_c21 <= X_27_c20;
               Y_27_c21 <= Y_27_c20;
            end if;
            if ce_22 = '1' then
               R_0_c22 <= R_0_c21;
               R_1_c22 <= R_1_c21;
               R_2_c22 <= R_2_c21;
               R_3_c22 <= R_3_c21;
               R_4_c22 <= R_4_c21;
               R_5_c22 <= R_5_c21;
               R_6_c22 <= R_6_c21;
               R_7_c22 <= R_7_c21;
               R_8_c22 <= R_8_c21;
               R_9_c22 <= R_9_c21;
               R_10_c22 <= R_10_c21;
               R_11_c22 <= R_11_c21;
               R_12_c22 <= R_12_c21;
               R_13_c22 <= R_13_c21;
               R_14_c22 <= R_14_c21;
               R_15_c22 <= R_15_c21;
               Cin_16_c22 <= Cin_16_c21;
               X_16_c22 <= X_16_c21;
               Y_16_c22 <= Y_16_c21;
               X_17_c22 <= X_17_c21;
               Y_17_c22 <= Y_17_c21;
               X_18_c22 <= X_18_c21;
               Y_18_c22 <= Y_18_c21;
               X_19_c22 <= X_19_c21;
               Y_19_c22 <= Y_19_c21;
               X_20_c22 <= X_20_c21;
               Y_20_c22 <= Y_20_c21;
               X_21_c22 <= X_21_c21;
               Y_21_c22 <= Y_21_c21;
               X_22_c22 <= X_22_c21;
               Y_22_c22 <= Y_22_c21;
               X_23_c22 <= X_23_c21;
               Y_23_c22 <= Y_23_c21;
               X_24_c22 <= X_24_c21;
               Y_24_c22 <= Y_24_c21;
               X_25_c22 <= X_25_c21;
               Y_25_c22 <= Y_25_c21;
               X_26_c22 <= X_26_c21;
               Y_26_c22 <= Y_26_c21;
               X_27_c22 <= X_27_c21;
               Y_27_c22 <= Y_27_c21;
            end if;
            if ce_23 = '1' then
               R_0_c23 <= R_0_c22;
               R_1_c23 <= R_1_c22;
               R_2_c23 <= R_2_c22;
               R_3_c23 <= R_3_c22;
               R_4_c23 <= R_4_c22;
               R_5_c23 <= R_5_c22;
               R_6_c23 <= R_6_c22;
               R_7_c23 <= R_7_c22;
               R_8_c23 <= R_8_c22;
               R_9_c23 <= R_9_c22;
               R_10_c23 <= R_10_c22;
               R_11_c23 <= R_11_c22;
               R_12_c23 <= R_12_c22;
               R_13_c23 <= R_13_c22;
               R_14_c23 <= R_14_c22;
               R_15_c23 <= R_15_c22;
               R_16_c23 <= R_16_c22;
               Cin_17_c23 <= Cin_17_c22;
               X_17_c23 <= X_17_c22;
               Y_17_c23 <= Y_17_c22;
               X_18_c23 <= X_18_c22;
               Y_18_c23 <= Y_18_c22;
               X_19_c23 <= X_19_c22;
               Y_19_c23 <= Y_19_c22;
               X_20_c23 <= X_20_c22;
               Y_20_c23 <= Y_20_c22;
               X_21_c23 <= X_21_c22;
               Y_21_c23 <= Y_21_c22;
               X_22_c23 <= X_22_c22;
               Y_22_c23 <= Y_22_c22;
               X_23_c23 <= X_23_c22;
               Y_23_c23 <= Y_23_c22;
               X_24_c23 <= X_24_c22;
               Y_24_c23 <= Y_24_c22;
               X_25_c23 <= X_25_c22;
               Y_25_c23 <= Y_25_c22;
               X_26_c23 <= X_26_c22;
               Y_26_c23 <= Y_26_c22;
               X_27_c23 <= X_27_c22;
               Y_27_c23 <= Y_27_c22;
            end if;
            if ce_24 = '1' then
               R_0_c24 <= R_0_c23;
               R_1_c24 <= R_1_c23;
               R_2_c24 <= R_2_c23;
               R_3_c24 <= R_3_c23;
               R_4_c24 <= R_4_c23;
               R_5_c24 <= R_5_c23;
               R_6_c24 <= R_6_c23;
               R_7_c24 <= R_7_c23;
               R_8_c24 <= R_8_c23;
               R_9_c24 <= R_9_c23;
               R_10_c24 <= R_10_c23;
               R_11_c24 <= R_11_c23;
               R_12_c24 <= R_12_c23;
               R_13_c24 <= R_13_c23;
               R_14_c24 <= R_14_c23;
               R_15_c24 <= R_15_c23;
               R_16_c24 <= R_16_c23;
               R_17_c24 <= R_17_c23;
               Cin_18_c24 <= Cin_18_c23;
               X_18_c24 <= X_18_c23;
               Y_18_c24 <= Y_18_c23;
               X_19_c24 <= X_19_c23;
               Y_19_c24 <= Y_19_c23;
               X_20_c24 <= X_20_c23;
               Y_20_c24 <= Y_20_c23;
               X_21_c24 <= X_21_c23;
               Y_21_c24 <= Y_21_c23;
               X_22_c24 <= X_22_c23;
               Y_22_c24 <= Y_22_c23;
               X_23_c24 <= X_23_c23;
               Y_23_c24 <= Y_23_c23;
               X_24_c24 <= X_24_c23;
               Y_24_c24 <= Y_24_c23;
               X_25_c24 <= X_25_c23;
               Y_25_c24 <= Y_25_c23;
               X_26_c24 <= X_26_c23;
               Y_26_c24 <= Y_26_c23;
               X_27_c24 <= X_27_c23;
               Y_27_c24 <= Y_27_c23;
            end if;
            if ce_25 = '1' then
               R_0_c25 <= R_0_c24;
               R_1_c25 <= R_1_c24;
               R_2_c25 <= R_2_c24;
               R_3_c25 <= R_3_c24;
               R_4_c25 <= R_4_c24;
               R_5_c25 <= R_5_c24;
               R_6_c25 <= R_6_c24;
               R_7_c25 <= R_7_c24;
               R_8_c25 <= R_8_c24;
               R_9_c25 <= R_9_c24;
               R_10_c25 <= R_10_c24;
               R_11_c25 <= R_11_c24;
               R_12_c25 <= R_12_c24;
               R_13_c25 <= R_13_c24;
               R_14_c25 <= R_14_c24;
               R_15_c25 <= R_15_c24;
               R_16_c25 <= R_16_c24;
               R_17_c25 <= R_17_c24;
               R_18_c25 <= R_18_c24;
               Cin_19_c25 <= Cin_19_c24;
               X_19_c25 <= X_19_c24;
               Y_19_c25 <= Y_19_c24;
               X_20_c25 <= X_20_c24;
               Y_20_c25 <= Y_20_c24;
               X_21_c25 <= X_21_c24;
               Y_21_c25 <= Y_21_c24;
               X_22_c25 <= X_22_c24;
               Y_22_c25 <= Y_22_c24;
               X_23_c25 <= X_23_c24;
               Y_23_c25 <= Y_23_c24;
               X_24_c25 <= X_24_c24;
               Y_24_c25 <= Y_24_c24;
               X_25_c25 <= X_25_c24;
               Y_25_c25 <= Y_25_c24;
               X_26_c25 <= X_26_c24;
               Y_26_c25 <= Y_26_c24;
               X_27_c25 <= X_27_c24;
               Y_27_c25 <= Y_27_c24;
            end if;
            if ce_26 = '1' then
               R_0_c26 <= R_0_c25;
               R_1_c26 <= R_1_c25;
               R_2_c26 <= R_2_c25;
               R_3_c26 <= R_3_c25;
               R_4_c26 <= R_4_c25;
               R_5_c26 <= R_5_c25;
               R_6_c26 <= R_6_c25;
               R_7_c26 <= R_7_c25;
               R_8_c26 <= R_8_c25;
               R_9_c26 <= R_9_c25;
               R_10_c26 <= R_10_c25;
               R_11_c26 <= R_11_c25;
               R_12_c26 <= R_12_c25;
               R_13_c26 <= R_13_c25;
               R_14_c26 <= R_14_c25;
               R_15_c26 <= R_15_c25;
               R_16_c26 <= R_16_c25;
               R_17_c26 <= R_17_c25;
               R_18_c26 <= R_18_c25;
               R_19_c26 <= R_19_c25;
               Cin_20_c26 <= Cin_20_c25;
               X_20_c26 <= X_20_c25;
               Y_20_c26 <= Y_20_c25;
               X_21_c26 <= X_21_c25;
               Y_21_c26 <= Y_21_c25;
               X_22_c26 <= X_22_c25;
               Y_22_c26 <= Y_22_c25;
               X_23_c26 <= X_23_c25;
               Y_23_c26 <= Y_23_c25;
               X_24_c26 <= X_24_c25;
               Y_24_c26 <= Y_24_c25;
               X_25_c26 <= X_25_c25;
               Y_25_c26 <= Y_25_c25;
               X_26_c26 <= X_26_c25;
               Y_26_c26 <= Y_26_c25;
               X_27_c26 <= X_27_c25;
               Y_27_c26 <= Y_27_c25;
            end if;
            if ce_27 = '1' then
               R_0_c27 <= R_0_c26;
               R_1_c27 <= R_1_c26;
               R_2_c27 <= R_2_c26;
               R_3_c27 <= R_3_c26;
               R_4_c27 <= R_4_c26;
               R_5_c27 <= R_5_c26;
               R_6_c27 <= R_6_c26;
               R_7_c27 <= R_7_c26;
               R_8_c27 <= R_8_c26;
               R_9_c27 <= R_9_c26;
               R_10_c27 <= R_10_c26;
               R_11_c27 <= R_11_c26;
               R_12_c27 <= R_12_c26;
               R_13_c27 <= R_13_c26;
               R_14_c27 <= R_14_c26;
               R_15_c27 <= R_15_c26;
               R_16_c27 <= R_16_c26;
               R_17_c27 <= R_17_c26;
               R_18_c27 <= R_18_c26;
               R_19_c27 <= R_19_c26;
               R_20_c27 <= R_20_c26;
               Cin_21_c27 <= Cin_21_c26;
               X_21_c27 <= X_21_c26;
               Y_21_c27 <= Y_21_c26;
               X_22_c27 <= X_22_c26;
               Y_22_c27 <= Y_22_c26;
               X_23_c27 <= X_23_c26;
               Y_23_c27 <= Y_23_c26;
               X_24_c27 <= X_24_c26;
               Y_24_c27 <= Y_24_c26;
               X_25_c27 <= X_25_c26;
               Y_25_c27 <= Y_25_c26;
               X_26_c27 <= X_26_c26;
               Y_26_c27 <= Y_26_c26;
               X_27_c27 <= X_27_c26;
               Y_27_c27 <= Y_27_c26;
            end if;
            if ce_28 = '1' then
               R_0_c28 <= R_0_c27;
               R_1_c28 <= R_1_c27;
               R_2_c28 <= R_2_c27;
               R_3_c28 <= R_3_c27;
               R_4_c28 <= R_4_c27;
               R_5_c28 <= R_5_c27;
               R_6_c28 <= R_6_c27;
               R_7_c28 <= R_7_c27;
               R_8_c28 <= R_8_c27;
               R_9_c28 <= R_9_c27;
               R_10_c28 <= R_10_c27;
               R_11_c28 <= R_11_c27;
               R_12_c28 <= R_12_c27;
               R_13_c28 <= R_13_c27;
               R_14_c28 <= R_14_c27;
               R_15_c28 <= R_15_c27;
               R_16_c28 <= R_16_c27;
               R_17_c28 <= R_17_c27;
               R_18_c28 <= R_18_c27;
               R_19_c28 <= R_19_c27;
               R_20_c28 <= R_20_c27;
               R_21_c28 <= R_21_c27;
               Cin_22_c28 <= Cin_22_c27;
               X_22_c28 <= X_22_c27;
               Y_22_c28 <= Y_22_c27;
               X_23_c28 <= X_23_c27;
               Y_23_c28 <= Y_23_c27;
               X_24_c28 <= X_24_c27;
               Y_24_c28 <= Y_24_c27;
               X_25_c28 <= X_25_c27;
               Y_25_c28 <= Y_25_c27;
               X_26_c28 <= X_26_c27;
               Y_26_c28 <= Y_26_c27;
               X_27_c28 <= X_27_c27;
               Y_27_c28 <= Y_27_c27;
            end if;
            if ce_29 = '1' then
               R_0_c29 <= R_0_c28;
               R_1_c29 <= R_1_c28;
               R_2_c29 <= R_2_c28;
               R_3_c29 <= R_3_c28;
               R_4_c29 <= R_4_c28;
               R_5_c29 <= R_5_c28;
               R_6_c29 <= R_6_c28;
               R_7_c29 <= R_7_c28;
               R_8_c29 <= R_8_c28;
               R_9_c29 <= R_9_c28;
               R_10_c29 <= R_10_c28;
               R_11_c29 <= R_11_c28;
               R_12_c29 <= R_12_c28;
               R_13_c29 <= R_13_c28;
               R_14_c29 <= R_14_c28;
               R_15_c29 <= R_15_c28;
               R_16_c29 <= R_16_c28;
               R_17_c29 <= R_17_c28;
               R_18_c29 <= R_18_c28;
               R_19_c29 <= R_19_c28;
               R_20_c29 <= R_20_c28;
               R_21_c29 <= R_21_c28;
               R_22_c29 <= R_22_c28;
               Cin_23_c29 <= Cin_23_c28;
               X_23_c29 <= X_23_c28;
               Y_23_c29 <= Y_23_c28;
               X_24_c29 <= X_24_c28;
               Y_24_c29 <= Y_24_c28;
               X_25_c29 <= X_25_c28;
               Y_25_c29 <= Y_25_c28;
               X_26_c29 <= X_26_c28;
               Y_26_c29 <= Y_26_c28;
               X_27_c29 <= X_27_c28;
               Y_27_c29 <= Y_27_c28;
            end if;
            if ce_30 = '1' then
               R_0_c30 <= R_0_c29;
               R_1_c30 <= R_1_c29;
               R_2_c30 <= R_2_c29;
               R_3_c30 <= R_3_c29;
               R_4_c30 <= R_4_c29;
               R_5_c30 <= R_5_c29;
               R_6_c30 <= R_6_c29;
               R_7_c30 <= R_7_c29;
               R_8_c30 <= R_8_c29;
               R_9_c30 <= R_9_c29;
               R_10_c30 <= R_10_c29;
               R_11_c30 <= R_11_c29;
               R_12_c30 <= R_12_c29;
               R_13_c30 <= R_13_c29;
               R_14_c30 <= R_14_c29;
               R_15_c30 <= R_15_c29;
               R_16_c30 <= R_16_c29;
               R_17_c30 <= R_17_c29;
               R_18_c30 <= R_18_c29;
               R_19_c30 <= R_19_c29;
               R_20_c30 <= R_20_c29;
               R_21_c30 <= R_21_c29;
               R_22_c30 <= R_22_c29;
               R_23_c30 <= R_23_c29;
               Cin_24_c30 <= Cin_24_c29;
               X_24_c30 <= X_24_c29;
               Y_24_c30 <= Y_24_c29;
               X_25_c30 <= X_25_c29;
               Y_25_c30 <= Y_25_c29;
               X_26_c30 <= X_26_c29;
               Y_26_c30 <= Y_26_c29;
               X_27_c30 <= X_27_c29;
               Y_27_c30 <= Y_27_c29;
            end if;
            if ce_31 = '1' then
               R_0_c31 <= R_0_c30;
               R_1_c31 <= R_1_c30;
               R_2_c31 <= R_2_c30;
               R_3_c31 <= R_3_c30;
               R_4_c31 <= R_4_c30;
               R_5_c31 <= R_5_c30;
               R_6_c31 <= R_6_c30;
               R_7_c31 <= R_7_c30;
               R_8_c31 <= R_8_c30;
               R_9_c31 <= R_9_c30;
               R_10_c31 <= R_10_c30;
               R_11_c31 <= R_11_c30;
               R_12_c31 <= R_12_c30;
               R_13_c31 <= R_13_c30;
               R_14_c31 <= R_14_c30;
               R_15_c31 <= R_15_c30;
               R_16_c31 <= R_16_c30;
               R_17_c31 <= R_17_c30;
               R_18_c31 <= R_18_c30;
               R_19_c31 <= R_19_c30;
               R_20_c31 <= R_20_c30;
               R_21_c31 <= R_21_c30;
               R_22_c31 <= R_22_c30;
               R_23_c31 <= R_23_c30;
               R_24_c31 <= R_24_c30;
               Cin_25_c31 <= Cin_25_c30;
               X_25_c31 <= X_25_c30;
               Y_25_c31 <= Y_25_c30;
               X_26_c31 <= X_26_c30;
               Y_26_c31 <= Y_26_c30;
               X_27_c31 <= X_27_c30;
               Y_27_c31 <= Y_27_c30;
            end if;
            if ce_32 = '1' then
               R_0_c32 <= R_0_c31;
               R_1_c32 <= R_1_c31;
               R_2_c32 <= R_2_c31;
               R_3_c32 <= R_3_c31;
               R_4_c32 <= R_4_c31;
               R_5_c32 <= R_5_c31;
               R_6_c32 <= R_6_c31;
               R_7_c32 <= R_7_c31;
               R_8_c32 <= R_8_c31;
               R_9_c32 <= R_9_c31;
               R_10_c32 <= R_10_c31;
               R_11_c32 <= R_11_c31;
               R_12_c32 <= R_12_c31;
               R_13_c32 <= R_13_c31;
               R_14_c32 <= R_14_c31;
               R_15_c32 <= R_15_c31;
               R_16_c32 <= R_16_c31;
               R_17_c32 <= R_17_c31;
               R_18_c32 <= R_18_c31;
               R_19_c32 <= R_19_c31;
               R_20_c32 <= R_20_c31;
               R_21_c32 <= R_21_c31;
               R_22_c32 <= R_22_c31;
               R_23_c32 <= R_23_c31;
               R_24_c32 <= R_24_c31;
               R_25_c32 <= R_25_c31;
               Cin_26_c32 <= Cin_26_c31;
               X_26_c32 <= X_26_c31;
               Y_26_c32 <= Y_26_c31;
               X_27_c32 <= X_27_c31;
               Y_27_c32 <= Y_27_c31;
            end if;
            if ce_33 = '1' then
               R_0_c33 <= R_0_c32;
               R_1_c33 <= R_1_c32;
               R_2_c33 <= R_2_c32;
               R_3_c33 <= R_3_c32;
               R_4_c33 <= R_4_c32;
               R_5_c33 <= R_5_c32;
               R_6_c33 <= R_6_c32;
               R_7_c33 <= R_7_c32;
               R_8_c33 <= R_8_c32;
               R_9_c33 <= R_9_c32;
               R_10_c33 <= R_10_c32;
               R_11_c33 <= R_11_c32;
               R_12_c33 <= R_12_c32;
               R_13_c33 <= R_13_c32;
               R_14_c33 <= R_14_c32;
               R_15_c33 <= R_15_c32;
               R_16_c33 <= R_16_c32;
               R_17_c33 <= R_17_c32;
               R_18_c33 <= R_18_c32;
               R_19_c33 <= R_19_c32;
               R_20_c33 <= R_20_c32;
               R_21_c33 <= R_21_c32;
               R_22_c33 <= R_22_c32;
               R_23_c33 <= R_23_c32;
               R_24_c33 <= R_24_c32;
               R_25_c33 <= R_25_c32;
               R_26_c33 <= R_26_c32;
               Cin_27_c33 <= Cin_27_c32;
               X_27_c33 <= X_27_c32;
               Y_27_c33 <= Y_27_c32;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c4 <= '0' & X(2 downto 0);
   Y_0_c4 <= '0' & Y(2 downto 0);
   S_0_c5 <= X_0_c5 + Y_0_c5 + Cin_0_c5;
   R_0_c5 <= S_0_c5(2 downto 0);
   Cin_1_c5 <= S_0_c5(3);
   X_1_c4 <= '0' & X(5 downto 3);
   Y_1_c4 <= '0' & Y(5 downto 3);
   S_1_c6 <= X_1_c6 + Y_1_c6 + Cin_1_c6;
   R_1_c6 <= S_1_c6(2 downto 0);
   Cin_2_c6 <= S_1_c6(3);
   X_2_c4 <= '0' & X(8 downto 6);
   Y_2_c4 <= '0' & Y(8 downto 6);
   S_2_c7 <= X_2_c7 + Y_2_c7 + Cin_2_c7;
   R_2_c7 <= S_2_c7(2 downto 0);
   Cin_3_c7 <= S_2_c7(3);
   X_3_c4 <= '0' & X(11 downto 9);
   Y_3_c4 <= '0' & Y(11 downto 9);
   S_3_c8 <= X_3_c8 + Y_3_c8 + Cin_3_c8;
   R_3_c8 <= S_3_c8(2 downto 0);
   Cin_4_c8 <= S_3_c8(3);
   X_4_c4 <= '0' & X(14 downto 12);
   Y_4_c4 <= '0' & Y(14 downto 12);
   S_4_c9 <= X_4_c9 + Y_4_c9 + Cin_4_c9;
   R_4_c9 <= S_4_c9(2 downto 0);
   Cin_5_c9 <= S_4_c9(3);
   X_5_c4 <= '0' & X(17 downto 15);
   Y_5_c4 <= '0' & Y(17 downto 15);
   S_5_c10 <= X_5_c10 + Y_5_c10 + Cin_5_c10;
   R_5_c10 <= S_5_c10(2 downto 0);
   Cin_6_c10 <= S_5_c10(3);
   X_6_c4 <= '0' & X(20 downto 18);
   Y_6_c4 <= '0' & Y(20 downto 18);
   S_6_c11 <= X_6_c11 + Y_6_c11 + Cin_6_c11;
   R_6_c11 <= S_6_c11(2 downto 0);
   Cin_7_c11 <= S_6_c11(3);
   X_7_c4 <= '0' & X(23 downto 21);
   Y_7_c4 <= '0' & Y(23 downto 21);
   S_7_c12 <= X_7_c12 + Y_7_c12 + Cin_7_c12;
   R_7_c12 <= S_7_c12(2 downto 0);
   Cin_8_c12 <= S_7_c12(3);
   X_8_c4 <= '0' & X(26 downto 24);
   Y_8_c4 <= '0' & Y(26 downto 24);
   S_8_c13 <= X_8_c13 + Y_8_c13 + Cin_8_c13;
   R_8_c13 <= S_8_c13(2 downto 0);
   Cin_9_c13 <= S_8_c13(3);
   X_9_c4 <= '0' & X(29 downto 27);
   Y_9_c4 <= '0' & Y(29 downto 27);
   S_9_c14 <= X_9_c14 + Y_9_c14 + Cin_9_c14;
   R_9_c14 <= S_9_c14(2 downto 0);
   Cin_10_c14 <= S_9_c14(3);
   X_10_c4 <= '0' & X(32 downto 30);
   Y_10_c4 <= '0' & Y(32 downto 30);
   S_10_c15 <= X_10_c15 + Y_10_c15 + Cin_10_c15;
   R_10_c15 <= S_10_c15(2 downto 0);
   Cin_11_c15 <= S_10_c15(3);
   X_11_c4 <= '0' & X(35 downto 33);
   Y_11_c4 <= '0' & Y(35 downto 33);
   S_11_c16 <= X_11_c16 + Y_11_c16 + Cin_11_c16;
   R_11_c16 <= S_11_c16(2 downto 0);
   Cin_12_c16 <= S_11_c16(3);
   X_12_c4 <= '0' & X(38 downto 36);
   Y_12_c4 <= '0' & Y(38 downto 36);
   S_12_c17 <= X_12_c17 + Y_12_c17 + Cin_12_c17;
   R_12_c17 <= S_12_c17(2 downto 0);
   Cin_13_c17 <= S_12_c17(3);
   X_13_c4 <= '0' & X(41 downto 39);
   Y_13_c4 <= '0' & Y(41 downto 39);
   S_13_c18 <= X_13_c18 + Y_13_c18 + Cin_13_c18;
   R_13_c18 <= S_13_c18(2 downto 0);
   Cin_14_c18 <= S_13_c18(3);
   X_14_c4 <= '0' & X(44 downto 42);
   Y_14_c4 <= '0' & Y(44 downto 42);
   S_14_c20 <= X_14_c20 + Y_14_c20 + Cin_14_c20;
   R_14_c20 <= S_14_c20(2 downto 0);
   Cin_15_c20 <= S_14_c20(3);
   X_15_c4 <= '0' & X(47 downto 45);
   Y_15_c4 <= '0' & Y(47 downto 45);
   S_15_c21 <= X_15_c21 + Y_15_c21 + Cin_15_c21;
   R_15_c21 <= S_15_c21(2 downto 0);
   Cin_16_c21 <= S_15_c21(3);
   X_16_c4 <= '0' & X(50 downto 48);
   Y_16_c4 <= '0' & Y(50 downto 48);
   S_16_c22 <= X_16_c22 + Y_16_c22 + Cin_16_c22;
   R_16_c22 <= S_16_c22(2 downto 0);
   Cin_17_c22 <= S_16_c22(3);
   X_17_c4 <= '0' & X(53 downto 51);
   Y_17_c4 <= '0' & Y(53 downto 51);
   S_17_c23 <= X_17_c23 + Y_17_c23 + Cin_17_c23;
   R_17_c23 <= S_17_c23(2 downto 0);
   Cin_18_c23 <= S_17_c23(3);
   X_18_c4 <= '0' & X(56 downto 54);
   Y_18_c4 <= '0' & Y(56 downto 54);
   S_18_c24 <= X_18_c24 + Y_18_c24 + Cin_18_c24;
   R_18_c24 <= S_18_c24(2 downto 0);
   Cin_19_c24 <= S_18_c24(3);
   X_19_c4 <= '0' & X(59 downto 57);
   Y_19_c4 <= '0' & Y(59 downto 57);
   S_19_c25 <= X_19_c25 + Y_19_c25 + Cin_19_c25;
   R_19_c25 <= S_19_c25(2 downto 0);
   Cin_20_c25 <= S_19_c25(3);
   X_20_c4 <= '0' & X(62 downto 60);
   Y_20_c4 <= '0' & Y(62 downto 60);
   S_20_c26 <= X_20_c26 + Y_20_c26 + Cin_20_c26;
   R_20_c26 <= S_20_c26(2 downto 0);
   Cin_21_c26 <= S_20_c26(3);
   X_21_c4 <= '0' & X(65 downto 63);
   Y_21_c4 <= '0' & Y(65 downto 63);
   S_21_c27 <= X_21_c27 + Y_21_c27 + Cin_21_c27;
   R_21_c27 <= S_21_c27(2 downto 0);
   Cin_22_c27 <= S_21_c27(3);
   X_22_c4 <= '0' & X(68 downto 66);
   Y_22_c4 <= '0' & Y(68 downto 66);
   S_22_c28 <= X_22_c28 + Y_22_c28 + Cin_22_c28;
   R_22_c28 <= S_22_c28(2 downto 0);
   Cin_23_c28 <= S_22_c28(3);
   X_23_c4 <= '0' & X(71 downto 69);
   Y_23_c4 <= '0' & Y(71 downto 69);
   S_23_c29 <= X_23_c29 + Y_23_c29 + Cin_23_c29;
   R_23_c29 <= S_23_c29(2 downto 0);
   Cin_24_c29 <= S_23_c29(3);
   X_24_c4 <= '0' & X(74 downto 72);
   Y_24_c4 <= '0' & Y(74 downto 72);
   S_24_c30 <= X_24_c30 + Y_24_c30 + Cin_24_c30;
   R_24_c30 <= S_24_c30(2 downto 0);
   Cin_25_c30 <= S_24_c30(3);
   X_25_c4 <= '0' & X(77 downto 75);
   Y_25_c4 <= '0' & Y(77 downto 75);
   S_25_c31 <= X_25_c31 + Y_25_c31 + Cin_25_c31;
   R_25_c31 <= S_25_c31(2 downto 0);
   Cin_26_c31 <= S_25_c31(3);
   X_26_c4 <= '0' & X(80 downto 78);
   Y_26_c4 <= '0' & Y(80 downto 78);
   S_26_c32 <= X_26_c32 + Y_26_c32 + Cin_26_c32;
   R_26_c32 <= S_26_c32(2 downto 0);
   Cin_27_c32 <= S_26_c32(3);
   X_27_c4 <= '0' & X(83 downto 81);
   Y_27_c4 <= '0' & Y(83 downto 81);
   S_27_c33 <= X_27_c33 + Y_27_c33 + Cin_27_c33;
   R_27_c33 <= S_27_c33(2 downto 0);
   R <= R_27_c33 & R_26_c33 & R_25_c33 & R_24_c33 & R_23_c33 & R_22_c33 & R_21_c33 & R_20_c33 & R_19_c33 & R_18_c33 & R_17_c33 & R_16_c33 & R_15_c33 & R_14_c33 & R_13_c33 & R_12_c33 & R_11_c33 & R_10_c33 & R_9_c33 & R_8_c33 & R_7_c33 & R_6_c33 & R_5_c33 & R_4_c33 & R_3_c33 & R_2_c33 & R_1_c33 & R_0_c33 ;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_53x53_106_Freq800_uid5
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 33 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_53x53_106_Freq800_uid5 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33 : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          Y : in  std_logic_vector(52 downto 0);
          R : out  std_logic_vector(105 downto 0)   );
end entity;

architecture arch of IntMultiplier_53x53_106_Freq800_uid5 is
   component DSPBlock_17x24_Freq800_uid9 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid11 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid13 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid15 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid20 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid35 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid40 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid45 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid50 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid55 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid57 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq800_uid59 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid61 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid66 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid76 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid81 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid86 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid91 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid96 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid101 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid103 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid105 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid107 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid109 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid111 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid116 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid126 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid131 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid136 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid141 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid146 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid151 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid156 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid161 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid166 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid171 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid173 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid175 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid177 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid179 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid181 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid186 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid191 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid196 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid201 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid206 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid211 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid216 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid221 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid226 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid231 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid236 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq800_uid241 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid243 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid245 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid247 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq800_uid249 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid251 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid256 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid261 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid266 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid271 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid276 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid281 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid286 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid291 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid296 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid301 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq800_uid306 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq800_uid311 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq800_uid316 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq800_uid322 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq800_uid326 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq800_uid334 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq800_uid400 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq800_uid432 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntAdder_84_Freq800_uid972 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33 : in std_logic;
             X : in  std_logic_vector(83 downto 0);
             Y : in  std_logic_vector(83 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(83 downto 0)   );
   end component;

signal XX_m6_c0 :  std_logic_vector(52 downto 0);
signal YY_m6_c0 :  std_logic_vector(52 downto 0);
signal tile_0_X_c0 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_0_output_c2 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w0_0_c2, bh7_w0_0_c3, bh7_w0_0_c4 :  std_logic;
signal bh7_w1_0_c2, bh7_w1_0_c3, bh7_w1_0_c4 :  std_logic;
signal bh7_w2_0_c2, bh7_w2_0_c3, bh7_w2_0_c4 :  std_logic;
signal bh7_w3_0_c2, bh7_w3_0_c3, bh7_w3_0_c4 :  std_logic;
signal bh7_w4_0_c2, bh7_w4_0_c3, bh7_w4_0_c4 :  std_logic;
signal bh7_w5_0_c2, bh7_w5_0_c3, bh7_w5_0_c4 :  std_logic;
signal bh7_w6_0_c2, bh7_w6_0_c3, bh7_w6_0_c4 :  std_logic;
signal bh7_w7_0_c2, bh7_w7_0_c3, bh7_w7_0_c4 :  std_logic;
signal bh7_w8_0_c2, bh7_w8_0_c3, bh7_w8_0_c4 :  std_logic;
signal bh7_w9_0_c2, bh7_w9_0_c3, bh7_w9_0_c4 :  std_logic;
signal bh7_w10_0_c2, bh7_w10_0_c3, bh7_w10_0_c4 :  std_logic;
signal bh7_w11_0_c2, bh7_w11_0_c3, bh7_w11_0_c4 :  std_logic;
signal bh7_w12_0_c2, bh7_w12_0_c3, bh7_w12_0_c4 :  std_logic;
signal bh7_w13_0_c2, bh7_w13_0_c3, bh7_w13_0_c4 :  std_logic;
signal bh7_w14_0_c2, bh7_w14_0_c3, bh7_w14_0_c4 :  std_logic;
signal bh7_w15_0_c2, bh7_w15_0_c3, bh7_w15_0_c4 :  std_logic;
signal bh7_w16_0_c2, bh7_w16_0_c3, bh7_w16_0_c4 :  std_logic;
signal bh7_w17_0_c2 :  std_logic;
signal bh7_w18_0_c2 :  std_logic;
signal bh7_w19_0_c2 :  std_logic;
signal bh7_w20_0_c2 :  std_logic;
signal bh7_w21_0_c2 :  std_logic;
signal bh7_w22_0_c2 :  std_logic;
signal bh7_w23_0_c2 :  std_logic;
signal bh7_w24_0_c2 :  std_logic;
signal bh7_w25_0_c2 :  std_logic;
signal bh7_w26_0_c2 :  std_logic;
signal bh7_w27_0_c2 :  std_logic;
signal bh7_w28_0_c2 :  std_logic;
signal bh7_w29_0_c2 :  std_logic;
signal bh7_w30_0_c2 :  std_logic;
signal bh7_w31_0_c2 :  std_logic;
signal bh7_w32_0_c2 :  std_logic;
signal bh7_w33_0_c2 :  std_logic;
signal bh7_w34_0_c2 :  std_logic;
signal bh7_w35_0_c2 :  std_logic;
signal bh7_w36_0_c2 :  std_logic;
signal bh7_w37_0_c2 :  std_logic;
signal bh7_w38_0_c2 :  std_logic;
signal bh7_w39_0_c2 :  std_logic;
signal bh7_w40_0_c2 :  std_logic;
signal tile_1_X_c0 :  std_logic_vector(16 downto 0);
signal tile_1_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_1_output_c2 :  std_logic_vector(40 downto 0);
signal tile_1_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w17_1_c2 :  std_logic;
signal bh7_w18_1_c2 :  std_logic;
signal bh7_w19_1_c2 :  std_logic;
signal bh7_w20_1_c2 :  std_logic;
signal bh7_w21_1_c2 :  std_logic;
signal bh7_w22_1_c2 :  std_logic;
signal bh7_w23_1_c2 :  std_logic;
signal bh7_w24_1_c2 :  std_logic;
signal bh7_w25_1_c2 :  std_logic;
signal bh7_w26_1_c2 :  std_logic;
signal bh7_w27_1_c2 :  std_logic;
signal bh7_w28_1_c2 :  std_logic;
signal bh7_w29_1_c2 :  std_logic;
signal bh7_w30_1_c2 :  std_logic;
signal bh7_w31_1_c2 :  std_logic;
signal bh7_w32_1_c2 :  std_logic;
signal bh7_w33_1_c2 :  std_logic;
signal bh7_w34_1_c2 :  std_logic;
signal bh7_w35_1_c2 :  std_logic;
signal bh7_w36_1_c2 :  std_logic;
signal bh7_w37_1_c2 :  std_logic;
signal bh7_w38_1_c2 :  std_logic;
signal bh7_w39_1_c2 :  std_logic;
signal bh7_w40_1_c2 :  std_logic;
signal bh7_w41_0_c2 :  std_logic;
signal bh7_w42_0_c2 :  std_logic;
signal bh7_w43_0_c2 :  std_logic;
signal bh7_w44_0_c2 :  std_logic;
signal bh7_w45_0_c2 :  std_logic;
signal bh7_w46_0_c2 :  std_logic;
signal bh7_w47_0_c2 :  std_logic;
signal bh7_w48_0_c2 :  std_logic;
signal bh7_w49_0_c2 :  std_logic;
signal bh7_w50_0_c2 :  std_logic;
signal bh7_w51_0_c2 :  std_logic;
signal bh7_w52_0_c2 :  std_logic;
signal bh7_w53_0_c2 :  std_logic;
signal bh7_w54_0_c2 :  std_logic;
signal bh7_w55_0_c2 :  std_logic;
signal bh7_w56_0_c2 :  std_logic;
signal bh7_w57_0_c2 :  std_logic;
signal tile_2_X_c0 :  std_logic_vector(16 downto 0);
signal tile_2_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_2_output_c2 :  std_logic_vector(40 downto 0);
signal tile_2_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w34_2_c2 :  std_logic;
signal bh7_w35_2_c2 :  std_logic;
signal bh7_w36_2_c2 :  std_logic;
signal bh7_w37_2_c2 :  std_logic;
signal bh7_w38_2_c2 :  std_logic;
signal bh7_w39_2_c2 :  std_logic;
signal bh7_w40_2_c2 :  std_logic;
signal bh7_w41_1_c2 :  std_logic;
signal bh7_w42_1_c2 :  std_logic;
signal bh7_w43_1_c2 :  std_logic;
signal bh7_w44_1_c2 :  std_logic;
signal bh7_w45_1_c2 :  std_logic;
signal bh7_w46_1_c2 :  std_logic;
signal bh7_w47_1_c2 :  std_logic;
signal bh7_w48_1_c2 :  std_logic;
signal bh7_w49_1_c2 :  std_logic;
signal bh7_w50_1_c2 :  std_logic;
signal bh7_w51_1_c2 :  std_logic;
signal bh7_w52_1_c2 :  std_logic;
signal bh7_w53_1_c2 :  std_logic;
signal bh7_w54_1_c2 :  std_logic;
signal bh7_w55_1_c2 :  std_logic;
signal bh7_w56_1_c2 :  std_logic;
signal bh7_w57_1_c2 :  std_logic;
signal bh7_w58_0_c2 :  std_logic;
signal bh7_w59_0_c2, bh7_w59_0_c3 :  std_logic;
signal bh7_w60_0_c2, bh7_w60_0_c3 :  std_logic;
signal bh7_w61_0_c2, bh7_w61_0_c3 :  std_logic;
signal bh7_w62_0_c2, bh7_w62_0_c3 :  std_logic;
signal bh7_w63_0_c2 :  std_logic;
signal bh7_w64_0_c2, bh7_w64_0_c3 :  std_logic;
signal bh7_w65_0_c2, bh7_w65_0_c3 :  std_logic;
signal bh7_w66_0_c2 :  std_logic;
signal bh7_w67_0_c2, bh7_w67_0_c3 :  std_logic;
signal bh7_w68_0_c2 :  std_logic;
signal bh7_w69_0_c2, bh7_w69_0_c3 :  std_logic;
signal bh7_w70_0_c2, bh7_w70_0_c3 :  std_logic;
signal bh7_w71_0_c2 :  std_logic;
signal bh7_w72_0_c2, bh7_w72_0_c3 :  std_logic;
signal bh7_w73_0_c2 :  std_logic;
signal bh7_w74_0_c2, bh7_w74_0_c3 :  std_logic;
signal tile_3_X_c0 :  std_logic_vector(1 downto 0);
signal tile_3_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_3_output_c0 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w72_1_c0 :  std_logic;
signal bh7_w73_1_c0 :  std_logic;
signal bh7_w74_1_c0 :  std_logic;
signal bh7_w75_0_c0 :  std_logic;
signal bh7_w76_0_c0 :  std_logic;
signal tile_4_X_c0 :  std_logic_vector(1 downto 0);
signal tile_4_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_4_output_c0 :  std_logic_vector(4 downto 0);
signal tile_4_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w69_1_c0 :  std_logic;
signal bh7_w70_1_c0 :  std_logic;
signal bh7_w71_1_c0 :  std_logic;
signal bh7_w72_2_c0 :  std_logic;
signal bh7_w73_2_c0 :  std_logic;
signal tile_5_X_c0 :  std_logic_vector(1 downto 0);
signal tile_5_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_5_output_c0 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w66_1_c0 :  std_logic;
signal bh7_w67_1_c0 :  std_logic;
signal bh7_w68_1_c0 :  std_logic;
signal bh7_w69_2_c0 :  std_logic;
signal bh7_w70_2_c0 :  std_logic;
signal tile_6_X_c0 :  std_logic_vector(1 downto 0);
signal tile_6_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_6_output_c0 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w63_1_c0 :  std_logic;
signal bh7_w64_1_c0 :  std_logic;
signal bh7_w65_1_c0 :  std_logic;
signal bh7_w66_2_c0 :  std_logic;
signal bh7_w67_2_c0 :  std_logic;
signal tile_7_X_c0 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_7_output_c0 :  std_logic_vector(4 downto 0);
signal tile_7_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_1_c0 :  std_logic;
signal bh7_w61_1_c0 :  std_logic;
signal bh7_w62_1_c0 :  std_logic;
signal bh7_w63_2_c0 :  std_logic;
signal bh7_w64_2_c0 :  std_logic;
signal tile_8_X_c0 :  std_logic_vector(1 downto 0);
signal tile_8_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_8_output_c0 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_2_c0 :  std_logic;
signal bh7_w58_1_c0 :  std_logic;
signal bh7_w59_1_c0 :  std_logic;
signal bh7_w60_2_c0 :  std_logic;
signal bh7_w61_2_c0 :  std_logic;
signal tile_9_X_c0 :  std_logic_vector(1 downto 0);
signal tile_9_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_9_output_c0 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_2_c0 :  std_logic;
signal bh7_w55_2_c0 :  std_logic;
signal bh7_w56_2_c0 :  std_logic;
signal bh7_w57_3_c0 :  std_logic;
signal bh7_w58_2_c0 :  std_logic;
signal tile_10_X_c0 :  std_logic_vector(1 downto 0);
signal tile_10_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_10_output_c0 :  std_logic_vector(4 downto 0);
signal tile_10_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_2_c0 :  std_logic;
signal bh7_w52_2_c0 :  std_logic;
signal bh7_w53_2_c0 :  std_logic;
signal bh7_w54_3_c0 :  std_logic;
signal bh7_w55_3_c0 :  std_logic;
signal tile_11_X_c0 :  std_logic_vector(16 downto 0);
signal tile_11_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_11_output_c2 :  std_logic_vector(40 downto 0);
signal tile_11_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w24_2_c2 :  std_logic;
signal bh7_w25_2_c2, bh7_w25_2_c3 :  std_logic;
signal bh7_w26_2_c2 :  std_logic;
signal bh7_w27_2_c2, bh7_w27_2_c3 :  std_logic;
signal bh7_w28_2_c2 :  std_logic;
signal bh7_w29_2_c2, bh7_w29_2_c3 :  std_logic;
signal bh7_w30_2_c2 :  std_logic;
signal bh7_w31_2_c2, bh7_w31_2_c3 :  std_logic;
signal bh7_w32_2_c2 :  std_logic;
signal bh7_w33_2_c2, bh7_w33_2_c3 :  std_logic;
signal bh7_w34_3_c2 :  std_logic;
signal bh7_w35_3_c2 :  std_logic;
signal bh7_w36_3_c2 :  std_logic;
signal bh7_w37_3_c2 :  std_logic;
signal bh7_w38_3_c2 :  std_logic;
signal bh7_w39_3_c2 :  std_logic;
signal bh7_w40_3_c2 :  std_logic;
signal bh7_w41_2_c2 :  std_logic;
signal bh7_w42_2_c2 :  std_logic;
signal bh7_w43_2_c2 :  std_logic;
signal bh7_w44_2_c2 :  std_logic;
signal bh7_w45_2_c2 :  std_logic;
signal bh7_w46_2_c2 :  std_logic;
signal bh7_w47_2_c2 :  std_logic;
signal bh7_w48_2_c2 :  std_logic;
signal bh7_w49_2_c2 :  std_logic;
signal bh7_w50_2_c2 :  std_logic;
signal bh7_w51_3_c2 :  std_logic;
signal bh7_w52_3_c2 :  std_logic;
signal bh7_w53_3_c2 :  std_logic;
signal bh7_w54_4_c2 :  std_logic;
signal bh7_w55_4_c2 :  std_logic;
signal bh7_w56_3_c2 :  std_logic;
signal bh7_w57_4_c2 :  std_logic;
signal bh7_w58_3_c2 :  std_logic;
signal bh7_w59_2_c2, bh7_w59_2_c3 :  std_logic;
signal bh7_w60_3_c2, bh7_w60_3_c3 :  std_logic;
signal bh7_w61_3_c2, bh7_w61_3_c3 :  std_logic;
signal bh7_w62_2_c2, bh7_w62_2_c3 :  std_logic;
signal bh7_w63_3_c2 :  std_logic;
signal bh7_w64_3_c2, bh7_w64_3_c3 :  std_logic;
signal tile_12_X_c0 :  std_logic_vector(16 downto 0);
signal tile_12_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_12_output_c2 :  std_logic_vector(40 downto 0);
signal tile_12_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w41_3_c2 :  std_logic;
signal bh7_w42_3_c2 :  std_logic;
signal bh7_w43_3_c2 :  std_logic;
signal bh7_w44_3_c2 :  std_logic;
signal bh7_w45_3_c2 :  std_logic;
signal bh7_w46_3_c2 :  std_logic;
signal bh7_w47_3_c2 :  std_logic;
signal bh7_w48_3_c2, bh7_w48_3_c3 :  std_logic;
signal bh7_w49_3_c2 :  std_logic;
signal bh7_w50_3_c2 :  std_logic;
signal bh7_w51_4_c2 :  std_logic;
signal bh7_w52_4_c2 :  std_logic;
signal bh7_w53_4_c2 :  std_logic;
signal bh7_w54_5_c2 :  std_logic;
signal bh7_w55_5_c2 :  std_logic;
signal bh7_w56_4_c2 :  std_logic;
signal bh7_w57_5_c2 :  std_logic;
signal bh7_w58_4_c2 :  std_logic;
signal bh7_w59_3_c2, bh7_w59_3_c3 :  std_logic;
signal bh7_w60_4_c2, bh7_w60_4_c3 :  std_logic;
signal bh7_w61_4_c2, bh7_w61_4_c3 :  std_logic;
signal bh7_w62_3_c2, bh7_w62_3_c3 :  std_logic;
signal bh7_w63_4_c2 :  std_logic;
signal bh7_w64_4_c2, bh7_w64_4_c3 :  std_logic;
signal bh7_w65_2_c2, bh7_w65_2_c3 :  std_logic;
signal bh7_w66_3_c2 :  std_logic;
signal bh7_w67_3_c2, bh7_w67_3_c3 :  std_logic;
signal bh7_w68_2_c2 :  std_logic;
signal bh7_w69_3_c2, bh7_w69_3_c3 :  std_logic;
signal bh7_w70_3_c2, bh7_w70_3_c3 :  std_logic;
signal bh7_w71_2_c2 :  std_logic;
signal bh7_w72_3_c2, bh7_w72_3_c3 :  std_logic;
signal bh7_w73_3_c2 :  std_logic;
signal bh7_w74_2_c2, bh7_w74_2_c3 :  std_logic;
signal bh7_w75_1_c2 :  std_logic;
signal bh7_w76_1_c2, bh7_w76_1_c3 :  std_logic;
signal bh7_w77_0_c2, bh7_w77_0_c3 :  std_logic;
signal bh7_w78_0_c2, bh7_w78_0_c3 :  std_logic;
signal bh7_w79_0_c2, bh7_w79_0_c3 :  std_logic;
signal bh7_w80_0_c2, bh7_w80_0_c3 :  std_logic;
signal bh7_w81_0_c2, bh7_w81_0_c3 :  std_logic;
signal tile_13_X_c0 :  std_logic_vector(16 downto 0);
signal tile_13_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_13_output_c2 :  std_logic_vector(40 downto 0);
signal tile_13_filtered_output_c2 :  unsigned(40-0 downto 0);
signal bh7_w58_5_c2, bh7_w58_5_c3 :  std_logic;
signal bh7_w59_4_c2, bh7_w59_4_c3 :  std_logic;
signal bh7_w60_5_c2, bh7_w60_5_c3 :  std_logic;
signal bh7_w61_5_c2, bh7_w61_5_c3 :  std_logic;
signal bh7_w62_4_c2, bh7_w62_4_c3 :  std_logic;
signal bh7_w63_5_c2, bh7_w63_5_c3 :  std_logic;
signal bh7_w64_5_c2, bh7_w64_5_c3 :  std_logic;
signal bh7_w65_3_c2, bh7_w65_3_c3 :  std_logic;
signal bh7_w66_4_c2 :  std_logic;
signal bh7_w67_4_c2, bh7_w67_4_c3 :  std_logic;
signal bh7_w68_3_c2 :  std_logic;
signal bh7_w69_4_c2, bh7_w69_4_c3 :  std_logic;
signal bh7_w70_4_c2, bh7_w70_4_c3 :  std_logic;
signal bh7_w71_3_c2 :  std_logic;
signal bh7_w72_4_c2, bh7_w72_4_c3 :  std_logic;
signal bh7_w73_4_c2 :  std_logic;
signal bh7_w74_3_c2, bh7_w74_3_c3 :  std_logic;
signal bh7_w75_2_c2, bh7_w75_2_c3 :  std_logic;
signal bh7_w76_2_c2, bh7_w76_2_c3 :  std_logic;
signal bh7_w77_1_c2, bh7_w77_1_c3 :  std_logic;
signal bh7_w78_1_c2, bh7_w78_1_c3 :  std_logic;
signal bh7_w79_1_c2, bh7_w79_1_c3 :  std_logic;
signal bh7_w80_1_c2, bh7_w80_1_c3 :  std_logic;
signal bh7_w81_1_c2, bh7_w81_1_c3 :  std_logic;
signal bh7_w82_0_c2, bh7_w82_0_c3 :  std_logic;
signal bh7_w83_0_c2, bh7_w83_0_c3 :  std_logic;
signal bh7_w84_0_c2, bh7_w84_0_c3 :  std_logic;
signal bh7_w85_0_c2, bh7_w85_0_c3 :  std_logic;
signal bh7_w86_0_c2, bh7_w86_0_c3 :  std_logic;
signal bh7_w87_0_c2, bh7_w87_0_c3 :  std_logic;
signal bh7_w88_0_c2, bh7_w88_0_c3 :  std_logic;
signal bh7_w89_0_c2, bh7_w89_0_c3 :  std_logic;
signal bh7_w90_0_c2, bh7_w90_0_c3 :  std_logic;
signal bh7_w91_0_c2, bh7_w91_0_c3 :  std_logic;
signal bh7_w92_0_c2, bh7_w92_0_c3 :  std_logic;
signal bh7_w93_0_c2, bh7_w93_0_c3 :  std_logic;
signal bh7_w94_0_c2, bh7_w94_0_c3 :  std_logic;
signal bh7_w95_0_c2, bh7_w95_0_c3 :  std_logic;
signal bh7_w96_0_c2, bh7_w96_0_c3 :  std_logic;
signal bh7_w97_0_c2, bh7_w97_0_c3 :  std_logic;
signal bh7_w98_0_c2, bh7_w98_0_c3 :  std_logic;
signal tile_14_X_c0 :  std_logic_vector(1 downto 0);
signal tile_14_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_14_output_c0 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_1_c0 :  std_logic;
signal bh7_w97_1_c0 :  std_logic;
signal bh7_w98_1_c0 :  std_logic;
signal bh7_w99_0_c0 :  std_logic;
signal bh7_w100_0_c0 :  std_logic;
signal tile_15_X_c0 :  std_logic_vector(1 downto 0);
signal tile_15_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_15_output_c0 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_1_c0 :  std_logic;
signal bh7_w94_1_c0 :  std_logic;
signal bh7_w95_1_c0 :  std_logic;
signal bh7_w96_2_c0 :  std_logic;
signal bh7_w97_2_c0 :  std_logic;
signal tile_16_X_c0 :  std_logic_vector(1 downto 0);
signal tile_16_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_16_output_c0 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_1_c0 :  std_logic;
signal bh7_w91_1_c0 :  std_logic;
signal bh7_w92_1_c0 :  std_logic;
signal bh7_w93_2_c0 :  std_logic;
signal bh7_w94_2_c0 :  std_logic;
signal tile_17_X_c0 :  std_logic_vector(1 downto 0);
signal tile_17_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_17_output_c0 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_1_c0 :  std_logic;
signal bh7_w88_1_c0 :  std_logic;
signal bh7_w89_1_c0 :  std_logic;
signal bh7_w90_2_c0 :  std_logic;
signal bh7_w91_2_c0 :  std_logic;
signal tile_18_X_c0 :  std_logic_vector(1 downto 0);
signal tile_18_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_18_output_c0 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_1_c0 :  std_logic;
signal bh7_w85_1_c0 :  std_logic;
signal bh7_w86_1_c0 :  std_logic;
signal bh7_w87_2_c0 :  std_logic;
signal bh7_w88_2_c0 :  std_logic;
signal tile_19_X_c0 :  std_logic_vector(1 downto 0);
signal tile_19_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_19_output_c0 :  std_logic_vector(4 downto 0);
signal tile_19_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w81_2_c0 :  std_logic;
signal bh7_w82_1_c0 :  std_logic;
signal bh7_w83_1_c0 :  std_logic;
signal bh7_w84_2_c0 :  std_logic;
signal bh7_w85_2_c0 :  std_logic;
signal tile_20_X_c0 :  std_logic_vector(1 downto 0);
signal tile_20_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_20_output_c0 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w78_2_c0 :  std_logic;
signal bh7_w79_2_c0 :  std_logic;
signal bh7_w80_2_c0 :  std_logic;
signal bh7_w81_3_c0 :  std_logic;
signal bh7_w82_2_c0 :  std_logic;
signal tile_21_X_c0 :  std_logic_vector(1 downto 0);
signal tile_21_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_21_output_c0 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w75_3_c0 :  std_logic;
signal bh7_w76_3_c0 :  std_logic;
signal bh7_w77_2_c0 :  std_logic;
signal bh7_w78_3_c0 :  std_logic;
signal bh7_w79_3_c0 :  std_logic;
signal tile_22_X_c0 :  std_logic_vector(0 downto 0);
signal tile_22_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_22_output_c0 :  std_logic_vector(0 downto 0);
signal tile_22_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w68_4_c0 :  std_logic;
signal tile_23_X_c0 :  std_logic_vector(3 downto 0);
signal tile_23_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_23_output_c0 :  std_logic_vector(3 downto 0);
signal tile_23_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w64_6_c0 :  std_logic;
signal bh7_w65_4_c0 :  std_logic;
signal bh7_w66_5_c0 :  std_logic;
signal bh7_w67_5_c0 :  std_logic;
signal tile_24_X_c0 :  std_logic_vector(3 downto 0);
signal tile_24_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_24_output_c0 :  std_logic_vector(3 downto 0);
signal tile_24_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w60_6_c0 :  std_logic;
signal bh7_w61_6_c0 :  std_logic;
signal bh7_w62_5_c0 :  std_logic;
signal bh7_w63_6_c0 :  std_logic;
signal tile_25_X_c0 :  std_logic_vector(3 downto 0);
signal tile_25_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_25_output_c0 :  std_logic_vector(3 downto 0);
signal tile_25_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w56_5_c0 :  std_logic;
signal bh7_w57_6_c0 :  std_logic;
signal bh7_w58_6_c0 :  std_logic;
signal bh7_w59_5_c0 :  std_logic;
signal tile_26_X_c0 :  std_logic_vector(3 downto 0);
signal tile_26_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_26_output_c0 :  std_logic_vector(3 downto 0);
signal tile_26_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w52_5_c0 :  std_logic;
signal bh7_w53_5_c0 :  std_logic;
signal bh7_w54_6_c0 :  std_logic;
signal bh7_w55_6_c0 :  std_logic;
signal tile_27_X_c0 :  std_logic_vector(1 downto 0);
signal tile_27_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_27_output_c0 :  std_logic_vector(3 downto 0);
signal tile_27_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w65_5_c0 :  std_logic;
signal bh7_w66_6_c0 :  std_logic;
signal bh7_w67_6_c0 :  std_logic;
signal bh7_w68_5_c0 :  std_logic;
signal tile_28_X_c0 :  std_logic_vector(2 downto 0);
signal tile_28_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_28_output_c0 :  std_logic_vector(4 downto 0);
signal tile_28_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w62_6_c0 :  std_logic;
signal bh7_w63_7_c0 :  std_logic;
signal bh7_w64_7_c0 :  std_logic;
signal bh7_w65_6_c0 :  std_logic;
signal bh7_w66_7_c0 :  std_logic;
signal tile_29_X_c0 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_29_output_c0 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w59_6_c0 :  std_logic;
signal bh7_w60_7_c0 :  std_logic;
signal bh7_w61_7_c0 :  std_logic;
signal bh7_w62_7_c0 :  std_logic;
signal bh7_w63_8_c0 :  std_logic;
signal tile_30_X_c0 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_30_output_c0 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w56_6_c0 :  std_logic;
signal bh7_w57_7_c0 :  std_logic;
signal bh7_w58_7_c0 :  std_logic;
signal bh7_w59_7_c0 :  std_logic;
signal bh7_w60_8_c0 :  std_logic;
signal tile_31_X_c0 :  std_logic_vector(2 downto 0);
signal tile_31_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_31_output_c0 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w53_6_c0 :  std_logic;
signal bh7_w54_7_c0 :  std_logic;
signal bh7_w55_7_c0 :  std_logic;
signal bh7_w56_7_c0 :  std_logic;
signal bh7_w57_8_c0 :  std_logic;
signal tile_32_X_c0 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_32_output_c0 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w50_4_c0 :  std_logic;
signal bh7_w51_5_c0 :  std_logic;
signal bh7_w52_6_c0 :  std_logic;
signal bh7_w53_7_c0 :  std_logic;
signal bh7_w54_8_c0 :  std_logic;
signal tile_33_X_c0 :  std_logic_vector(1 downto 0);
signal tile_33_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_33_output_c0 :  std_logic_vector(3 downto 0);
signal tile_33_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w63_9_c0 :  std_logic;
signal bh7_w64_8_c0 :  std_logic;
signal bh7_w65_7_c0 :  std_logic;
signal bh7_w66_8_c0 :  std_logic;
signal tile_34_X_c0 :  std_logic_vector(2 downto 0);
signal tile_34_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_34_output_c0 :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_9_c0 :  std_logic;
signal bh7_w61_8_c0 :  std_logic;
signal bh7_w62_8_c0, bh7_w62_8_c1 :  std_logic;
signal bh7_w63_10_c0 :  std_logic;
signal bh7_w64_9_c0 :  std_logic;
signal tile_35_X_c0 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_35_output_c0 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_9_c0 :  std_logic;
signal bh7_w58_8_c0 :  std_logic;
signal bh7_w59_8_c0, bh7_w59_8_c1 :  std_logic;
signal bh7_w60_10_c0 :  std_logic;
signal bh7_w61_9_c0 :  std_logic;
signal tile_36_X_c0 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_36_output_c0 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_9_c0 :  std_logic;
signal bh7_w55_8_c0 :  std_logic;
signal bh7_w56_8_c0, bh7_w56_8_c1 :  std_logic;
signal bh7_w57_10_c0 :  std_logic;
signal bh7_w58_9_c0 :  std_logic;
signal tile_37_X_c0 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_37_output_c0 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_6_c0 :  std_logic;
signal bh7_w52_7_c0 :  std_logic;
signal bh7_w53_8_c0 :  std_logic;
signal bh7_w54_10_c0 :  std_logic;
signal bh7_w55_9_c0 :  std_logic;
signal tile_38_X_c0 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_38_output_c0 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w48_4_c0, bh7_w48_4_c1, bh7_w48_4_c2 :  std_logic;
signal bh7_w49_4_c0 :  std_logic;
signal bh7_w50_5_c0 :  std_logic;
signal bh7_w51_7_c0 :  std_logic;
signal bh7_w52_8_c0 :  std_logic;
signal tile_39_X_c0 :  std_logic_vector(0 downto 0);
signal tile_39_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_39_output_c0 :  std_logic_vector(0 downto 0);
signal tile_39_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w85_3_c0 :  std_logic;
signal tile_40_X_c0 :  std_logic_vector(3 downto 0);
signal tile_40_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_40_output_c0 :  std_logic_vector(3 downto 0);
signal tile_40_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w81_4_c0 :  std_logic;
signal bh7_w82_3_c0 :  std_logic;
signal bh7_w83_2_c0 :  std_logic;
signal bh7_w84_3_c0 :  std_logic;
signal tile_41_X_c0 :  std_logic_vector(3 downto 0);
signal tile_41_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_41_output_c0 :  std_logic_vector(3 downto 0);
signal tile_41_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w77_3_c0 :  std_logic;
signal bh7_w78_4_c0 :  std_logic;
signal bh7_w79_4_c0 :  std_logic;
signal bh7_w80_3_c0 :  std_logic;
signal tile_42_X_c0 :  std_logic_vector(3 downto 0);
signal tile_42_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_42_output_c0 :  std_logic_vector(3 downto 0);
signal tile_42_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w73_5_c0 :  std_logic;
signal bh7_w74_4_c0 :  std_logic;
signal bh7_w75_4_c0 :  std_logic;
signal bh7_w76_4_c0 :  std_logic;
signal tile_43_X_c0 :  std_logic_vector(3 downto 0);
signal tile_43_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_43_output_c0 :  std_logic_vector(3 downto 0);
signal tile_43_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w69_5_c0 :  std_logic;
signal bh7_w70_5_c0 :  std_logic;
signal bh7_w71_4_c0 :  std_logic;
signal bh7_w72_5_c0 :  std_logic;
signal tile_44_X_c0 :  std_logic_vector(1 downto 0);
signal tile_44_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_44_output_c0 :  std_logic_vector(3 downto 0);
signal tile_44_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w82_4_c0 :  std_logic;
signal bh7_w83_3_c0 :  std_logic;
signal bh7_w84_4_c0 :  std_logic;
signal bh7_w85_4_c0 :  std_logic;
signal tile_45_X_c0 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_45_output_c0 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w79_5_c0 :  std_logic;
signal bh7_w80_4_c0 :  std_logic;
signal bh7_w81_5_c0 :  std_logic;
signal bh7_w82_5_c0 :  std_logic;
signal bh7_w83_4_c0 :  std_logic;
signal tile_46_X_c0 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_46_output_c0 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w76_5_c0 :  std_logic;
signal bh7_w77_4_c0 :  std_logic;
signal bh7_w78_5_c0 :  std_logic;
signal bh7_w79_6_c0 :  std_logic;
signal bh7_w80_5_c0 :  std_logic;
signal tile_47_X_c0 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_47_output_c0 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w73_6_c0 :  std_logic;
signal bh7_w74_5_c0 :  std_logic;
signal bh7_w75_5_c0 :  std_logic;
signal bh7_w76_6_c0 :  std_logic;
signal bh7_w77_5_c0 :  std_logic;
signal tile_48_X_c0 :  std_logic_vector(2 downto 0);
signal tile_48_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_48_output_c0 :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w70_6_c0 :  std_logic;
signal bh7_w71_5_c0 :  std_logic;
signal bh7_w72_6_c0 :  std_logic;
signal bh7_w73_7_c0 :  std_logic;
signal bh7_w74_6_c0 :  std_logic;
signal tile_49_X_c0 :  std_logic_vector(2 downto 0);
signal tile_49_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_49_output_c0 :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w67_7_c0 :  std_logic;
signal bh7_w68_6_c0 :  std_logic;
signal bh7_w69_6_c0 :  std_logic;
signal bh7_w70_7_c0 :  std_logic;
signal bh7_w71_6_c0 :  std_logic;
signal tile_50_X_c0 :  std_logic_vector(1 downto 0);
signal tile_50_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_50_output_c0 :  std_logic_vector(3 downto 0);
signal tile_50_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w80_6_c0 :  std_logic;
signal bh7_w81_6_c0 :  std_logic;
signal bh7_w82_6_c0 :  std_logic;
signal bh7_w83_5_c0 :  std_logic;
signal tile_51_X_c0 :  std_logic_vector(2 downto 0);
signal tile_51_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_51_output_c0 :  std_logic_vector(4 downto 0);
signal tile_51_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w77_6_c0 :  std_logic;
signal bh7_w78_6_c0 :  std_logic;
signal bh7_w79_7_c0 :  std_logic;
signal bh7_w80_7_c0 :  std_logic;
signal bh7_w81_7_c0 :  std_logic;
signal tile_52_X_c0 :  std_logic_vector(2 downto 0);
signal tile_52_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_52_output_c0 :  std_logic_vector(4 downto 0);
signal tile_52_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w74_7_c0 :  std_logic;
signal bh7_w75_6_c0 :  std_logic;
signal bh7_w76_7_c0 :  std_logic;
signal bh7_w77_7_c0 :  std_logic;
signal bh7_w78_7_c0 :  std_logic;
signal tile_53_X_c0 :  std_logic_vector(2 downto 0);
signal tile_53_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_53_output_c0 :  std_logic_vector(4 downto 0);
signal tile_53_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w71_7_c0 :  std_logic;
signal bh7_w72_7_c0 :  std_logic;
signal bh7_w73_8_c0 :  std_logic;
signal bh7_w74_8_c0 :  std_logic;
signal bh7_w75_7_c0 :  std_logic;
signal tile_54_X_c0 :  std_logic_vector(2 downto 0);
signal tile_54_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_54_output_c0 :  std_logic_vector(4 downto 0);
signal tile_54_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w68_7_c0 :  std_logic;
signal bh7_w69_7_c0 :  std_logic;
signal bh7_w70_8_c0 :  std_logic;
signal bh7_w71_8_c0 :  std_logic;
signal bh7_w72_8_c0 :  std_logic;
signal tile_55_X_c0 :  std_logic_vector(2 downto 0);
signal tile_55_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_55_output_c0 :  std_logic_vector(4 downto 0);
signal tile_55_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w65_8_c0 :  std_logic;
signal bh7_w66_9_c0, bh7_w66_9_c1 :  std_logic;
signal bh7_w67_8_c0 :  std_logic;
signal bh7_w68_8_c0 :  std_logic;
signal bh7_w69_8_c0 :  std_logic;
signal tile_56_X_c0 :  std_logic_vector(0 downto 0);
signal tile_56_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_56_output_c0 :  std_logic_vector(0 downto 0);
signal tile_56_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w102_0_c0 :  std_logic;
signal tile_57_X_c0 :  std_logic_vector(3 downto 0);
signal tile_57_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_57_output_c0 :  std_logic_vector(3 downto 0);
signal tile_57_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w98_2_c0 :  std_logic;
signal bh7_w99_1_c0 :  std_logic;
signal bh7_w100_1_c0 :  std_logic;
signal bh7_w101_0_c0 :  std_logic;
signal tile_58_X_c0 :  std_logic_vector(3 downto 0);
signal tile_58_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_58_output_c0 :  std_logic_vector(3 downto 0);
signal tile_58_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w94_3_c0 :  std_logic;
signal bh7_w95_2_c0 :  std_logic;
signal bh7_w96_3_c0 :  std_logic;
signal bh7_w97_3_c0 :  std_logic;
signal tile_59_X_c0 :  std_logic_vector(3 downto 0);
signal tile_59_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_59_output_c0 :  std_logic_vector(3 downto 0);
signal tile_59_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w90_3_c0 :  std_logic;
signal bh7_w91_3_c0 :  std_logic;
signal bh7_w92_2_c0 :  std_logic;
signal bh7_w93_3_c0 :  std_logic;
signal tile_60_X_c0 :  std_logic_vector(3 downto 0);
signal tile_60_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_60_output_c0 :  std_logic_vector(3 downto 0);
signal tile_60_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w86_2_c0 :  std_logic;
signal bh7_w87_3_c0 :  std_logic;
signal bh7_w88_3_c0 :  std_logic;
signal bh7_w89_2_c0 :  std_logic;
signal tile_61_X_c0 :  std_logic_vector(1 downto 0);
signal tile_61_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_61_output_c0 :  std_logic_vector(3 downto 0);
signal tile_61_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w99_2_c0 :  std_logic;
signal bh7_w100_2_c0 :  std_logic;
signal bh7_w101_1_c0 :  std_logic;
signal bh7_w102_1_c0 :  std_logic;
signal tile_62_X_c0 :  std_logic_vector(2 downto 0);
signal tile_62_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_62_output_c0 :  std_logic_vector(4 downto 0);
signal tile_62_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_4_c0 :  std_logic;
signal bh7_w97_4_c0 :  std_logic;
signal bh7_w98_3_c0 :  std_logic;
signal bh7_w99_3_c0 :  std_logic;
signal bh7_w100_3_c0 :  std_logic;
signal tile_63_X_c0 :  std_logic_vector(2 downto 0);
signal tile_63_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_63_output_c0 :  std_logic_vector(4 downto 0);
signal tile_63_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_4_c0 :  std_logic;
signal bh7_w94_4_c0 :  std_logic;
signal bh7_w95_3_c0 :  std_logic;
signal bh7_w96_5_c0 :  std_logic;
signal bh7_w97_5_c0 :  std_logic;
signal tile_64_X_c0 :  std_logic_vector(2 downto 0);
signal tile_64_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_64_output_c0 :  std_logic_vector(4 downto 0);
signal tile_64_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_4_c0 :  std_logic;
signal bh7_w91_4_c0 :  std_logic;
signal bh7_w92_3_c0 :  std_logic;
signal bh7_w93_5_c0 :  std_logic;
signal bh7_w94_5_c0 :  std_logic;
signal tile_65_X_c0 :  std_logic_vector(2 downto 0);
signal tile_65_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_65_output_c0 :  std_logic_vector(4 downto 0);
signal tile_65_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_4_c0 :  std_logic;
signal bh7_w88_4_c0 :  std_logic;
signal bh7_w89_3_c0 :  std_logic;
signal bh7_w90_5_c0 :  std_logic;
signal bh7_w91_5_c0 :  std_logic;
signal tile_66_X_c0 :  std_logic_vector(2 downto 0);
signal tile_66_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_66_output_c0 :  std_logic_vector(4 downto 0);
signal tile_66_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_5_c0 :  std_logic;
signal bh7_w85_5_c0 :  std_logic;
signal bh7_w86_3_c0 :  std_logic;
signal bh7_w87_5_c0 :  std_logic;
signal bh7_w88_5_c0 :  std_logic;
signal tile_67_X_c0 :  std_logic_vector(1 downto 0);
signal tile_67_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_67_output_c0 :  std_logic_vector(3 downto 0);
signal tile_67_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w97_6_c0 :  std_logic;
signal bh7_w98_4_c0 :  std_logic;
signal bh7_w99_4_c0 :  std_logic;
signal bh7_w100_4_c0 :  std_logic;
signal tile_68_X_c0 :  std_logic_vector(2 downto 0);
signal tile_68_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_68_output_c0 :  std_logic_vector(4 downto 0);
signal tile_68_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w94_6_c0 :  std_logic;
signal bh7_w95_4_c0 :  std_logic;
signal bh7_w96_6_c0 :  std_logic;
signal bh7_w97_7_c0, bh7_w97_7_c1 :  std_logic;
signal bh7_w98_5_c0 :  std_logic;
signal tile_69_X_c0 :  std_logic_vector(2 downto 0);
signal tile_69_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_69_output_c0 :  std_logic_vector(4 downto 0);
signal tile_69_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w91_6_c0 :  std_logic;
signal bh7_w92_4_c0 :  std_logic;
signal bh7_w93_6_c0 :  std_logic;
signal bh7_w94_7_c0, bh7_w94_7_c1 :  std_logic;
signal bh7_w95_5_c0 :  std_logic;
signal tile_70_X_c0 :  std_logic_vector(2 downto 0);
signal tile_70_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_70_output_c0 :  std_logic_vector(4 downto 0);
signal tile_70_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w88_6_c0 :  std_logic;
signal bh7_w89_4_c0 :  std_logic;
signal bh7_w90_6_c0 :  std_logic;
signal bh7_w91_7_c0, bh7_w91_7_c1 :  std_logic;
signal bh7_w92_5_c0 :  std_logic;
signal tile_71_X_c0 :  std_logic_vector(2 downto 0);
signal tile_71_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_71_output_c0 :  std_logic_vector(4 downto 0);
signal tile_71_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w85_6_c0 :  std_logic;
signal bh7_w86_4_c0 :  std_logic;
signal bh7_w87_6_c0 :  std_logic;
signal bh7_w88_7_c0, bh7_w88_7_c1 :  std_logic;
signal bh7_w89_5_c0 :  std_logic;
signal tile_72_X_c0 :  std_logic_vector(2 downto 0);
signal tile_72_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_72_output_c0 :  std_logic_vector(4 downto 0);
signal tile_72_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w82_7_c0, bh7_w82_7_c1 :  std_logic;
signal bh7_w83_6_c0 :  std_logic;
signal bh7_w84_6_c0 :  std_logic;
signal bh7_w85_7_c0, bh7_w85_7_c1 :  std_logic;
signal bh7_w86_5_c0 :  std_logic;
signal tile_73_X_c0 :  std_logic_vector(1 downto 0);
signal tile_73_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_73_output_c0 :  std_logic_vector(3 downto 0);
signal tile_73_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w102_2_c0 :  std_logic;
signal bh7_w103_0_c0 :  std_logic;
signal bh7_w104_0_c0, bh7_w104_0_c1 :  std_logic;
signal bh7_w105_0_c0, bh7_w105_0_c1 :  std_logic;
signal tile_74_X_c0 :  std_logic_vector(1 downto 0);
signal tile_74_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_74_output_c0 :  std_logic_vector(4 downto 0);
signal tile_74_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w99_5_c0 :  std_logic;
signal bh7_w100_5_c0 :  std_logic;
signal bh7_w101_2_c0 :  std_logic;
signal bh7_w102_3_c0 :  std_logic;
signal bh7_w103_1_c0, bh7_w103_1_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid323_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid323_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w49_5_c1 :  std_logic;
signal bh7_w50_6_c1 :  std_logic;
signal bh7_w51_8_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c0, Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid327_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid327_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w51_9_c1 :  std_logic;
signal bh7_w52_9_c1 :  std_logic;
signal bh7_w53_9_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c0, Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid329_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid329_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w52_10_c1 :  std_logic;
signal bh7_w53_10_c1 :  std_logic;
signal bh7_w54_11_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c0, Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid331_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid331_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w53_11_c1 :  std_logic;
signal bh7_w54_12_c1 :  std_logic;
signal bh7_w55_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c0, Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid335_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w54_13_c1 :  std_logic;
signal bh7_w55_11_c1 :  std_logic;
signal bh7_w56_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c0, Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid337_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w55_12_c1 :  std_logic;
signal bh7_w56_10_c1 :  std_logic;
signal bh7_w57_11_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c0, Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid339_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid339_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_11_c1 :  std_logic;
signal bh7_w57_12_c1 :  std_logic;
signal bh7_w58_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c0, Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid341_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w57_13_c1 :  std_logic;
signal bh7_w58_11_c1 :  std_logic;
signal bh7_w59_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c0, Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid343_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w58_12_c1 :  std_logic;
signal bh7_w59_10_c1 :  std_logic;
signal bh7_w60_11_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c0, Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid345_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid345_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_11_c1 :  std_logic;
signal bh7_w60_12_c1 :  std_logic;
signal bh7_w61_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c0, Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid347_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w60_13_c1 :  std_logic;
signal bh7_w61_11_c1 :  std_logic;
signal bh7_w62_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c0, Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid349_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w61_12_c1 :  std_logic;
signal bh7_w62_10_c1 :  std_logic;
signal bh7_w63_11_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c0, Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid351_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid351_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_11_c1 :  std_logic;
signal bh7_w63_12_c1 :  std_logic;
signal bh7_w64_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c0, Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid353_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w63_13_c1 :  std_logic;
signal bh7_w64_11_c1 :  std_logic;
signal bh7_w65_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c0, Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid355_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_12_c1 :  std_logic;
signal bh7_w65_10_c1 :  std_logic;
signal bh7_w66_10_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c0, Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid357_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w65_11_c1 :  std_logic;
signal bh7_w66_11_c1 :  std_logic;
signal bh7_w67_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c0, Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid359_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w66_12_c1 :  std_logic;
signal bh7_w67_10_c1 :  std_logic;
signal bh7_w68_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c0, Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid361_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w67_11_c1 :  std_logic;
signal bh7_w68_10_c1 :  std_logic;
signal bh7_w69_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c0, Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid363_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_11_c1 :  std_logic;
signal bh7_w69_10_c1 :  std_logic;
signal bh7_w70_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c0, Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid365_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w69_11_c1 :  std_logic;
signal bh7_w70_10_c1 :  std_logic;
signal bh7_w71_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c0, Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid367_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_11_c1 :  std_logic;
signal bh7_w71_10_c1 :  std_logic;
signal bh7_w72_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c0, Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid369_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w71_11_c1 :  std_logic;
signal bh7_w72_10_c1 :  std_logic;
signal bh7_w73_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c0, Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid371_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_11_c1 :  std_logic;
signal bh7_w73_10_c1 :  std_logic;
signal bh7_w74_9_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c0, Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid373_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w73_11_c1 :  std_logic;
signal bh7_w74_10_c1 :  std_logic;
signal bh7_w75_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c0, Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid375_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_11_c1 :  std_logic;
signal bh7_w75_9_c1 :  std_logic;
signal bh7_w76_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c0, Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid377_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w75_10_c1 :  std_logic;
signal bh7_w76_9_c1 :  std_logic;
signal bh7_w77_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c0, Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid379_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_10_c1 :  std_logic;
signal bh7_w77_9_c1 :  std_logic;
signal bh7_w78_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c0, Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid381_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w77_10_c1 :  std_logic;
signal bh7_w78_9_c1 :  std_logic;
signal bh7_w79_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c0, Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid383_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_10_c1 :  std_logic;
signal bh7_w79_9_c1 :  std_logic;
signal bh7_w80_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c0, Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid385_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w79_10_c1 :  std_logic;
signal bh7_w80_9_c1 :  std_logic;
signal bh7_w81_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c0, Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid387_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_10_c1 :  std_logic;
signal bh7_w81_9_c1 :  std_logic;
signal bh7_w82_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c0, Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid389_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w81_10_c1 :  std_logic;
signal bh7_w82_9_c1 :  std_logic;
signal bh7_w83_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c0, Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid391_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_10_c1 :  std_logic;
signal bh7_w83_8_c1 :  std_logic;
signal bh7_w84_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c0, Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid393_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w83_9_c1 :  std_logic;
signal bh7_w84_8_c1 :  std_logic;
signal bh7_w85_8_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c0, Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid395_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_9_c1 :  std_logic;
signal bh7_w85_9_c1 :  std_logic;
signal bh7_w86_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c0, Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid397_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w85_10_c1 :  std_logic;
signal bh7_w86_7_c1 :  std_logic;
signal bh7_w87_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c0, Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid401_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_8_c1 :  std_logic;
signal bh7_w87_8_c1 :  std_logic;
signal bh7_w88_8_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c0, Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid403_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w87_9_c1 :  std_logic;
signal bh7_w88_9_c1 :  std_logic;
signal bh7_w89_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c0, Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid405_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_10_c1 :  std_logic;
signal bh7_w89_7_c1 :  std_logic;
signal bh7_w90_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c0, Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid407_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w89_8_c1 :  std_logic;
signal bh7_w90_8_c1 :  std_logic;
signal bh7_w91_8_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c0, Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid409_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w90_9_c1 :  std_logic;
signal bh7_w91_9_c1 :  std_logic;
signal bh7_w92_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c0, Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid411_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w91_10_c1 :  std_logic;
signal bh7_w92_7_c1 :  std_logic;
signal bh7_w93_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c0, Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid413_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w92_8_c1 :  std_logic;
signal bh7_w93_8_c1 :  std_logic;
signal bh7_w94_8_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c0, Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid415_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w93_9_c1 :  std_logic;
signal bh7_w94_9_c1 :  std_logic;
signal bh7_w95_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c0, Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid417_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w94_10_c1 :  std_logic;
signal bh7_w95_7_c1 :  std_logic;
signal bh7_w96_7_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c0, Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid419_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w95_8_c1 :  std_logic;
signal bh7_w96_8_c1 :  std_logic;
signal bh7_w97_8_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c0, Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid421_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w96_9_c1 :  std_logic;
signal bh7_w97_9_c1 :  std_logic;
signal bh7_w98_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c0, Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid423_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w97_10_c1 :  std_logic;
signal bh7_w98_7_c1 :  std_logic;
signal bh7_w99_6_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c0, Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid425_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w98_8_c1 :  std_logic;
signal bh7_w99_7_c1 :  std_logic;
signal bh7_w100_6_c1 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c0, Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid427_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w99_8_c1 :  std_logic;
signal bh7_w100_7_c1 :  std_logic;
signal bh7_w101_3_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c0, Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid429_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w100_8_c1 :  std_logic;
signal bh7_w101_4_c1 :  std_logic;
signal bh7_w102_4_c1 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c0, Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid433_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w101_5_c1 :  std_logic;
signal bh7_w102_5_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c0, Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid435_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid435_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w102_6_c1 :  std_logic;
signal bh7_w103_2_c1 :  std_logic;
signal bh7_w104_1_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c0, Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid437_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid437_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w51_10_c1 :  std_logic;
signal bh7_w52_11_c1 :  std_logic;
signal bh7_w53_12_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_copy438_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid439_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid439_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w53_13_c1 :  std_logic;
signal bh7_w54_14_c1 :  std_logic;
signal bh7_w55_13_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_copy440_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid441_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w55_14_c1 :  std_logic;
signal bh7_w56_12_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_copy442_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid443_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_13_c1 :  std_logic;
signal bh7_w57_14_c1 :  std_logic;
signal bh7_w58_13_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_copy444_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid445_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w57_15_c1 :  std_logic;
signal bh7_w58_14_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_copy446_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid447_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w58_15_c1 :  std_logic;
signal bh7_w59_12_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_copy448_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid449_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_13_c1 :  std_logic;
signal bh7_w60_14_c1 :  std_logic;
signal bh7_w61_13_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_copy450_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid451_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w60_15_c1 :  std_logic;
signal bh7_w61_14_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_copy452_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid453_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w61_15_c1 :  std_logic;
signal bh7_w62_12_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_copy454_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid455_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_13_c1 :  std_logic;
signal bh7_w63_14_c1 :  std_logic;
signal bh7_w64_13_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_copy456_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid457_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w63_15_c1 :  std_logic;
signal bh7_w64_14_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_copy458_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid459_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid459_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_15_c1 :  std_logic;
signal bh7_w65_12_c1 :  std_logic;
signal bh7_w66_13_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_copy460_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid461_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w66_14_c1 :  std_logic;
signal bh7_w67_12_c1 :  std_logic;
signal bh7_w68_12_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_copy462_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid463_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w67_13_c1 :  std_logic;
signal bh7_w68_13_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_copy464_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid465_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid465_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_14_c1 :  std_logic;
signal bh7_w69_12_c1 :  std_logic;
signal bh7_w70_12_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_copy466_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid467_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid467_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_13_c1 :  std_logic;
signal bh7_w71_12_c1 :  std_logic;
signal bh7_w72_12_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_copy468_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid469_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid469_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_13_c1 :  std_logic;
signal bh7_w73_12_c1 :  std_logic;
signal bh7_w74_12_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_copy470_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid471_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid471_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_13_c1 :  std_logic;
signal bh7_w75_11_c1 :  std_logic;
signal bh7_w76_11_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_copy472_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid473_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid473_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_12_c1 :  std_logic;
signal bh7_w77_11_c1 :  std_logic;
signal bh7_w78_11_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_copy474_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid475_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid475_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_12_c1 :  std_logic;
signal bh7_w79_11_c1 :  std_logic;
signal bh7_w80_11_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_copy476_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid477_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid477_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_12_c1 :  std_logic;
signal bh7_w81_11_c1 :  std_logic;
signal bh7_w82_11_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_copy478_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid479_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_12_c1 :  std_logic;
signal bh7_w83_10_c1 :  std_logic;
signal bh7_w84_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_copy480_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid481_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w83_11_c1 :  std_logic;
signal bh7_w84_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_copy482_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid483_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w84_12_c1 :  std_logic;
signal bh7_w85_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_copy484_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid485_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w85_12_c1 :  std_logic;
signal bh7_w86_9_c1 :  std_logic;
signal bh7_w87_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_copy486_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid487_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w86_10_c1 :  std_logic;
signal bh7_w87_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_copy488_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid489_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w87_12_c1 :  std_logic;
signal bh7_w88_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_copy490_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid491_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_12_c1 :  std_logic;
signal bh7_w89_9_c1 :  std_logic;
signal bh7_w90_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_copy492_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid493_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w89_10_c1 :  std_logic;
signal bh7_w90_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_copy494_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid495_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w90_12_c1 :  std_logic;
signal bh7_w91_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_copy496_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid497_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w91_12_c1 :  std_logic;
signal bh7_w92_9_c1 :  std_logic;
signal bh7_w93_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_copy498_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid499_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w92_10_c1 :  std_logic;
signal bh7_w93_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_copy500_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid501_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w93_12_c1 :  std_logic;
signal bh7_w94_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_copy502_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid503_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w94_12_c1 :  std_logic;
signal bh7_w95_9_c1 :  std_logic;
signal bh7_w96_10_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_copy504_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid505_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w95_10_c1 :  std_logic;
signal bh7_w96_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_copy506_c1 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid507_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w96_12_c1 :  std_logic;
signal bh7_w97_11_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_copy508_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid509_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w97_12_c1 :  std_logic;
signal bh7_w98_9_c1 :  std_logic;
signal bh7_w99_9_c1 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_copy510_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid511_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w98_10_c1 :  std_logic;
signal bh7_w99_10_c1 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_copy512_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid513_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid513_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w99_11_c1 :  std_logic;
signal bh7_w100_9_c1 :  std_logic;
signal bh7_w101_6_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_copy514_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid515_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid515_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w101_7_c1 :  std_logic;
signal bh7_w102_7_c1 :  std_logic;
signal bh7_w103_3_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_copy516_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid517_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid517_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w103_4_c1 :  std_logic;
signal bh7_w104_2_c1 :  std_logic;
signal bh7_w105_1_c1 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_copy518_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid519_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid519_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w53_14_c2 :  std_logic;
signal bh7_w54_15_c2 :  std_logic;
signal bh7_w55_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c1, Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid521_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid521_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w55_16_c2 :  std_logic;
signal bh7_w56_14_c2 :  std_logic;
signal bh7_w57_16_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c1, Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid523_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w57_17_c2 :  std_logic;
signal bh7_w58_16_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c1, Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid525_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid525_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w58_17_c2 :  std_logic;
signal bh7_w59_14_c2 :  std_logic;
signal bh7_w60_16_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c1, Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid527_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w60_17_c2 :  std_logic;
signal bh7_w61_16_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c1, Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid529_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid529_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w61_17_c2 :  std_logic;
signal bh7_w62_14_c2 :  std_logic;
signal bh7_w63_16_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c1, Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid531_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w63_17_c2 :  std_logic;
signal bh7_w64_16_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c1, Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid533_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid533_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w64_17_c2 :  std_logic;
signal bh7_w65_13_c2 :  std_logic;
signal bh7_w66_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c1, Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid535_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid535_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w66_16_c2 :  std_logic;
signal bh7_w67_14_c2 :  std_logic;
signal bh7_w68_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c1, Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid537_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid537_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w68_16_c2 :  std_logic;
signal bh7_w69_13_c2 :  std_logic;
signal bh7_w70_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c1, Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid539_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid539_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w70_15_c2 :  std_logic;
signal bh7_w71_13_c2 :  std_logic;
signal bh7_w72_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c1, Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid541_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid541_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w72_15_c2 :  std_logic;
signal bh7_w73_13_c2 :  std_logic;
signal bh7_w74_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c1, Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid543_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid543_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w74_15_c2 :  std_logic;
signal bh7_w75_12_c2 :  std_logic;
signal bh7_w76_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c1, Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid545_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid545_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w76_14_c2 :  std_logic;
signal bh7_w77_12_c2 :  std_logic;
signal bh7_w78_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c1, Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid547_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid547_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w78_14_c2 :  std_logic;
signal bh7_w79_12_c2 :  std_logic;
signal bh7_w80_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c1, Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid549_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid549_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w80_14_c2 :  std_logic;
signal bh7_w81_12_c2 :  std_logic;
signal bh7_w82_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c1, Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid551_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid551_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w82_14_c2 :  std_logic;
signal bh7_w83_12_c2 :  std_logic;
signal bh7_w84_13_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c1, Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid553_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid553_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w84_14_c2 :  std_logic;
signal bh7_w85_13_c2 :  std_logic;
signal bh7_w86_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c1, Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid555_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w86_12_c2 :  std_logic;
signal bh7_w87_13_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c1, Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid557_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid557_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w87_14_c2 :  std_logic;
signal bh7_w88_13_c2 :  std_logic;
signal bh7_w89_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c1, Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid559_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w89_12_c2 :  std_logic;
signal bh7_w90_13_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c1, Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid561_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid561_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w90_14_c2 :  std_logic;
signal bh7_w91_13_c2 :  std_logic;
signal bh7_w92_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c1, Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid563_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w92_12_c2 :  std_logic;
signal bh7_w93_13_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c1, Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid565_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid565_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w93_14_c2 :  std_logic;
signal bh7_w94_13_c2 :  std_logic;
signal bh7_w95_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c1, Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid567_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w95_12_c2 :  std_logic;
signal bh7_w96_13_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c1, Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid569_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid569_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w96_14_c2 :  std_logic;
signal bh7_w97_13_c2 :  std_logic;
signal bh7_w98_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c1, Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid571_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w98_12_c2 :  std_logic;
signal bh7_w99_12_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c1, Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid573_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid573_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w99_13_c2 :  std_logic;
signal bh7_w100_10_c2 :  std_logic;
signal bh7_w101_8_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c1, Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid575_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid575_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w101_9_c2 :  std_logic;
signal bh7_w102_8_c2 :  std_logic;
signal bh7_w103_5_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c1, Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid577_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid577_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w103_6_c2 :  std_logic;
signal bh7_w104_3_c2 :  std_logic;
signal bh7_w105_2_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c1, Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid579_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w105_3_c2 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c1, Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c2 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid581_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid581_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w55_17_c2 :  std_logic;
signal bh7_w56_15_c2 :  std_logic;
signal bh7_w57_18_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_copy582_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid583_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid583_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w57_19_c2 :  std_logic;
signal bh7_w58_18_c2 :  std_logic;
signal bh7_w59_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_copy584_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid585_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid585_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w60_18_c2 :  std_logic;
signal bh7_w61_18_c2, bh7_w61_18_c3 :  std_logic;
signal bh7_w62_15_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_copy586_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid587_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid587_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w63_18_c2 :  std_logic;
signal bh7_w64_18_c2, bh7_w64_18_c3 :  std_logic;
signal bh7_w65_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_copy588_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid589_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid589_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w66_17_c2 :  std_logic;
signal bh7_w67_15_c2, bh7_w67_15_c3 :  std_logic;
signal bh7_w68_17_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_copy590_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid591_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid591_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w68_18_c2 :  std_logic;
signal bh7_w69_14_c2 :  std_logic;
signal bh7_w70_16_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_copy592_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid593_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid593_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w70_17_c2 :  std_logic;
signal bh7_w71_14_c2 :  std_logic;
signal bh7_w72_16_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_copy594_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid595_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid595_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w72_17_c2 :  std_logic;
signal bh7_w73_14_c2 :  std_logic;
signal bh7_w74_16_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_copy596_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid597_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid597_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w74_17_c2 :  std_logic;
signal bh7_w75_13_c2 :  std_logic;
signal bh7_w76_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_copy598_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid599_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid599_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w76_16_c2 :  std_logic;
signal bh7_w77_13_c2 :  std_logic;
signal bh7_w78_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_copy600_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid601_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid601_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w78_16_c2 :  std_logic;
signal bh7_w79_13_c2 :  std_logic;
signal bh7_w80_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_copy602_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid603_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid603_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w80_16_c2 :  std_logic;
signal bh7_w81_13_c2 :  std_logic;
signal bh7_w82_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_copy604_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid605_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid605_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w82_16_c2 :  std_logic;
signal bh7_w83_13_c2 :  std_logic;
signal bh7_w84_15_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_copy606_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid607_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid607_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w84_16_c2 :  std_logic;
signal bh7_w85_14_c2 :  std_logic;
signal bh7_w86_13_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_copy608_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid609_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid609_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w86_14_c2 :  std_logic;
signal bh7_w87_15_c2 :  std_logic;
signal bh7_w88_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_copy610_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid611_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid611_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w89_13_c2 :  std_logic;
signal bh7_w90_15_c2, bh7_w90_15_c3 :  std_logic;
signal bh7_w91_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_copy612_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid613_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid613_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w92_13_c2 :  std_logic;
signal bh7_w93_15_c2, bh7_w93_15_c3 :  std_logic;
signal bh7_w94_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_copy614_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid615_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid615_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w95_13_c2 :  std_logic;
signal bh7_w96_15_c2, bh7_w96_15_c3 :  std_logic;
signal bh7_w97_14_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_copy616_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid617_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid617_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w98_13_c2 :  std_logic;
signal bh7_w99_14_c2, bh7_w99_14_c3 :  std_logic;
signal bh7_w100_11_c2 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_copy618_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid619_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid619_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w101_10_c2 :  std_logic;
signal bh7_w102_9_c2, bh7_w102_9_c3 :  std_logic;
signal bh7_w103_7_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_copy620_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid621_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid621_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w103_8_c2 :  std_logic;
signal bh7_w104_4_c2 :  std_logic;
signal bh7_w105_4_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_copy622_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid623_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w105_5_c2 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_copy624_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid625_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid625_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w57_20_c3 :  std_logic;
signal bh7_w58_19_c3 :  std_logic;
signal bh7_w59_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c2, Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid627_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid627_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w59_17_c3 :  std_logic;
signal bh7_w60_19_c3 :  std_logic;
signal bh7_w61_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c2, Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid629_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid629_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w62_16_c3 :  std_logic;
signal bh7_w63_19_c3 :  std_logic;
signal bh7_w64_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c2, Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid631_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid631_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w65_15_c3 :  std_logic;
signal bh7_w66_18_c3 :  std_logic;
signal bh7_w67_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c2, Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid633_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid633_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w68_19_c3 :  std_logic;
signal bh7_w69_15_c3 :  std_logic;
signal bh7_w70_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c2, Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid635_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid635_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w70_19_c3 :  std_logic;
signal bh7_w71_15_c3 :  std_logic;
signal bh7_w72_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c2, Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid637_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid637_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w72_19_c3 :  std_logic;
signal bh7_w73_15_c3 :  std_logic;
signal bh7_w74_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c2, Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid639_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid639_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w74_19_c3 :  std_logic;
signal bh7_w75_14_c3 :  std_logic;
signal bh7_w76_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c2, Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid641_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid641_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w76_18_c3 :  std_logic;
signal bh7_w77_14_c3 :  std_logic;
signal bh7_w78_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c2, Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid643_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid643_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w78_18_c3 :  std_logic;
signal bh7_w79_14_c3 :  std_logic;
signal bh7_w80_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c2, Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid645_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid645_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w80_18_c3 :  std_logic;
signal bh7_w81_14_c3 :  std_logic;
signal bh7_w82_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c2, Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid647_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid647_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w82_18_c3 :  std_logic;
signal bh7_w83_14_c3 :  std_logic;
signal bh7_w84_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c2, Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid649_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid649_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w84_18_c3 :  std_logic;
signal bh7_w85_15_c3 :  std_logic;
signal bh7_w86_15_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c2, Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid651_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid651_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w86_16_c3 :  std_logic;
signal bh7_w87_16_c3 :  std_logic;
signal bh7_w88_15_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c2, Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid653_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid653_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w88_16_c3 :  std_logic;
signal bh7_w89_14_c3 :  std_logic;
signal bh7_w90_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c2, Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid655_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid655_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w91_15_c3 :  std_logic;
signal bh7_w92_14_c3 :  std_logic;
signal bh7_w93_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c2, Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid657_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid657_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w94_15_c3 :  std_logic;
signal bh7_w95_14_c3 :  std_logic;
signal bh7_w96_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c2, Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid659_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid659_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w97_15_c3 :  std_logic;
signal bh7_w98_14_c3 :  std_logic;
signal bh7_w99_15_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c2, Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid661_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid661_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w100_12_c3 :  std_logic;
signal bh7_w101_11_c3 :  std_logic;
signal bh7_w102_10_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c2, Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid663_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid663_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w103_9_c3 :  std_logic;
signal bh7_w104_5_c3 :  std_logic;
signal bh7_w105_6_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c2, Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid665_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w105_7_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c2, Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid667_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid667_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w17_2_c3, bh7_w17_2_c4 :  std_logic;
signal bh7_w18_2_c3, bh7_w18_2_c4 :  std_logic;
signal bh7_w19_2_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c2, Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid669_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid669_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w19_3_c3 :  std_logic;
signal bh7_w20_2_c3 :  std_logic;
signal bh7_w21_2_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c2, Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid671_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid671_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w21_3_c3 :  std_logic;
signal bh7_w22_2_c3 :  std_logic;
signal bh7_w23_2_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c2, Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid673_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w23_3_c3 :  std_logic;
signal bh7_w24_3_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c2, Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid675_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid675_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w24_4_c3 :  std_logic;
signal bh7_w25_3_c3 :  std_logic;
signal bh7_w26_3_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c2, Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid677_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid677_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w26_4_c3 :  std_logic;
signal bh7_w27_3_c3 :  std_logic;
signal bh7_w28_3_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c2, Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid679_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid679_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w28_4_c3 :  std_logic;
signal bh7_w29_3_c3 :  std_logic;
signal bh7_w30_3_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c2, Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid681_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid681_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w30_4_c3 :  std_logic;
signal bh7_w31_3_c3 :  std_logic;
signal bh7_w32_3_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c2, Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid683_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid683_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w32_4_c3 :  std_logic;
signal bh7_w33_3_c3 :  std_logic;
signal bh7_w34_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c2, Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid685_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid685_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w34_5_c3 :  std_logic;
signal bh7_w35_4_c3 :  std_logic;
signal bh7_w36_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c2, Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid687_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w35_5_c3 :  std_logic;
signal bh7_w36_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c2, Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid689_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid689_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w36_6_c3 :  std_logic;
signal bh7_w37_4_c3 :  std_logic;
signal bh7_w38_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c2, Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid691_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w37_5_c3 :  std_logic;
signal bh7_w38_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c2, Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid693_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid693_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w38_6_c3 :  std_logic;
signal bh7_w39_4_c3 :  std_logic;
signal bh7_w40_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c2, Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid695_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w39_5_c3 :  std_logic;
signal bh7_w40_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c2, Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid697_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid697_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w40_6_c3 :  std_logic;
signal bh7_w41_4_c3 :  std_logic;
signal bh7_w42_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c2, Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid699_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w41_5_c3 :  std_logic;
signal bh7_w42_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c2, Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid701_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid701_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w42_6_c3 :  std_logic;
signal bh7_w43_4_c3 :  std_logic;
signal bh7_w44_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c2, Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid703_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w43_5_c3 :  std_logic;
signal bh7_w44_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c2, Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid705_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid705_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w44_6_c3 :  std_logic;
signal bh7_w45_4_c3 :  std_logic;
signal bh7_w46_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c2, Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid707_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w45_5_c3 :  std_logic;
signal bh7_w46_5_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c2, Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid709_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid709_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w46_6_c3 :  std_logic;
signal bh7_w47_4_c3 :  std_logic;
signal bh7_w48_5_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c2, Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid711_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w47_5_c3 :  std_logic;
signal bh7_w48_6_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c2, Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid713_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w48_7_c3 :  std_logic;
signal bh7_w49_6_c3 :  std_logic;
signal bh7_w50_7_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c2, Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid715_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w49_7_c3 :  std_logic;
signal bh7_w50_8_c3 :  std_logic;
signal bh7_w51_11_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c2, Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid717_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w50_9_c3 :  std_logic;
signal bh7_w51_12_c3 :  std_logic;
signal bh7_w52_12_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c2, Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid719_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w51_13_c3 :  std_logic;
signal bh7_w52_13_c3 :  std_logic;
signal bh7_w53_15_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c2, Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid721_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid721_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w52_14_c3 :  std_logic;
signal bh7_w53_16_c3 :  std_logic;
signal bh7_w54_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c2, Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid723_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid723_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w53_17_c3 :  std_logic;
signal bh7_w54_17_c3 :  std_logic;
signal bh7_w55_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c2, Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid725_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid725_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w54_18_c3 :  std_logic;
signal bh7_w55_19_c3 :  std_logic;
signal bh7_w56_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c2, Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid727_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid727_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w55_20_c3 :  std_logic;
signal bh7_w56_17_c3 :  std_logic;
signal bh7_w57_21_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c2, Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c2, Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid729_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w56_18_c3 :  std_logic;
signal bh7_w57_22_c3 :  std_logic;
signal bh7_w58_20_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_copy730_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c2, Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid731_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w57_23_c3, bh7_w57_23_c4 :  std_logic;
signal bh7_w58_21_c3 :  std_logic;
signal bh7_w59_18_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_copy732_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid733_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w58_22_c3 :  std_logic;
signal bh7_w59_19_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c2, Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c3 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid735_In0_c3 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w59_20_c3 :  std_logic;
signal bh7_w60_20_c3 :  std_logic;
signal bh7_w61_20_c3 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_copy736_c3 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid737_In0_c3 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w60_21_c3 :  std_logic;
signal bh7_w61_21_c3 :  std_logic;
signal bh7_w62_17_c3 :  std_logic;
signal Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_copy738_c3 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid739_In0_c3 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w61_22_c3 :  std_logic;
signal bh7_w62_18_c3 :  std_logic;
signal bh7_w63_20_c3 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_copy740_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid741_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid741_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w62_19_c3 :  std_logic;
signal bh7_w63_21_c3 :  std_logic;
signal bh7_w64_20_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_copy742_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid743_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w63_22_c3 :  std_logic;
signal bh7_w64_21_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c2, Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c3 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid745_In0_c3 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w64_22_c3 :  std_logic;
signal bh7_w65_16_c3 :  std_logic;
signal bh7_w66_19_c3 :  std_logic;
signal Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_copy746_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid747_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid747_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w65_17_c3 :  std_logic;
signal bh7_w66_20_c3 :  std_logic;
signal bh7_w67_17_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_copy748_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid749_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w66_21_c3 :  std_logic;
signal bh7_w67_18_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c2, Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid751_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid751_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w67_19_c3 :  std_logic;
signal bh7_w68_20_c3 :  std_logic;
signal bh7_w69_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_copy752_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid753_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w68_21_c3, bh7_w68_21_c4 :  std_logic;
signal bh7_w69_17_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c2, Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid755_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid755_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w69_18_c3 :  std_logic;
signal bh7_w70_20_c3 :  std_logic;
signal bh7_w71_16_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_copy756_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid757_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid757_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w70_21_c3 :  std_logic;
signal bh7_w71_17_c3 :  std_logic;
signal bh7_w72_20_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_copy758_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid759_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w71_18_c3 :  std_logic;
signal bh7_w72_21_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c2, Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid761_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid761_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w72_22_c3 :  std_logic;
signal bh7_w73_16_c3 :  std_logic;
signal bh7_w74_20_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_copy762_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid763_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w73_17_c3, bh7_w73_17_c4 :  std_logic;
signal bh7_w74_21_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c2, Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid765_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w74_22_c3 :  std_logic;
signal bh7_w75_15_c3 :  std_logic;
signal bh7_w76_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_copy766_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid767_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid767_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w74_23_c3 :  std_logic;
signal bh7_w75_16_c3, bh7_w75_16_c4 :  std_logic;
signal bh7_w76_20_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_copy768_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid769_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w76_21_c3 :  std_logic;
signal bh7_w77_15_c3 :  std_logic;
signal bh7_w78_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_copy770_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid771_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w77_16_c3 :  std_logic;
signal bh7_w78_20_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_copy772_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid773_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w78_21_c3 :  std_logic;
signal bh7_w79_15_c3 :  std_logic;
signal bh7_w80_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_copy774_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid775_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w79_16_c3 :  std_logic;
signal bh7_w80_20_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_copy776_c3 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid777_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w80_21_c3 :  std_logic;
signal bh7_w81_15_c3 :  std_logic;
signal bh7_w82_19_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_copy778_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid779_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w81_16_c3 :  std_logic;
signal bh7_w82_20_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_copy780_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid781_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid781_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w82_21_c3 :  std_logic;
signal bh7_w83_15_c3, bh7_w83_15_c4 :  std_logic;
signal bh7_w84_19_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_copy782_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid783_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid783_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w84_20_c3 :  std_logic;
signal bh7_w85_16_c3 :  std_logic;
signal bh7_w86_17_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_copy784_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid785_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid785_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w86_18_c3 :  std_logic;
signal bh7_w87_17_c3 :  std_logic;
signal bh7_w88_17_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_copy786_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid787_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid787_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w88_18_c3 :  std_logic;
signal bh7_w89_15_c3 :  std_logic;
signal bh7_w90_17_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_copy788_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid789_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid789_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w90_18_c3 :  std_logic;
signal bh7_w91_16_c3 :  std_logic;
signal bh7_w92_15_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_copy790_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid791_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w92_16_c3 :  std_logic;
signal bh7_w93_17_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_copy792_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid793_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid793_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w93_18_c3 :  std_logic;
signal bh7_w94_16_c3, bh7_w94_16_c4 :  std_logic;
signal bh7_w95_15_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_copy794_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid795_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w95_16_c3 :  std_logic;
signal bh7_w96_17_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_copy796_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid797_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid797_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w96_18_c3 :  std_logic;
signal bh7_w97_16_c3, bh7_w97_16_c4 :  std_logic;
signal bh7_w98_15_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_copy798_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid799_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid799_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w98_16_c3 :  std_logic;
signal bh7_w99_16_c3 :  std_logic;
signal bh7_w100_13_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_copy800_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid801_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid801_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w102_11_c3, bh7_w102_11_c4 :  std_logic;
signal bh7_w103_10_c3 :  std_logic;
signal bh7_w104_6_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_copy802_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid803_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w105_8_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_copy804_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid805_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid805_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w19_4_c3, bh7_w19_4_c4 :  std_logic;
signal bh7_w20_3_c3, bh7_w20_3_c4 :  std_logic;
signal bh7_w21_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_copy806_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid807_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid807_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w21_5_c3 :  std_logic;
signal bh7_w22_3_c3 :  std_logic;
signal bh7_w23_4_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_copy808_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid809_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid809_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w23_5_c3 :  std_logic;
signal bh7_w24_5_c3 :  std_logic;
signal bh7_w25_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_copy810_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid811_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid811_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w25_5_c3 :  std_logic;
signal bh7_w26_5_c3 :  std_logic;
signal bh7_w27_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_copy812_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid813_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid813_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w27_5_c3 :  std_logic;
signal bh7_w28_5_c3 :  std_logic;
signal bh7_w29_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_copy814_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid815_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid815_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w29_5_c3 :  std_logic;
signal bh7_w30_5_c3 :  std_logic;
signal bh7_w31_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_copy816_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid817_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid817_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w31_5_c3 :  std_logic;
signal bh7_w32_5_c3 :  std_logic;
signal bh7_w33_4_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_copy818_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid819_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid819_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w33_5_c3 :  std_logic;
signal bh7_w34_6_c3 :  std_logic;
signal bh7_w35_6_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_copy820_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid821_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_c3 :  std_logic_vector(1 downto 0);
signal bh7_w35_7_c3 :  std_logic;
signal bh7_w36_7_c3 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_copy822_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid823_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid823_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w36_8_c3 :  std_logic;
signal bh7_w37_6_c3, bh7_w37_6_c4 :  std_logic;
signal bh7_w38_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_copy824_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid825_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid825_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w38_8_c3 :  std_logic;
signal bh7_w39_6_c3 :  std_logic;
signal bh7_w40_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_copy826_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid827_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid827_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w40_8_c3 :  std_logic;
signal bh7_w41_6_c3 :  std_logic;
signal bh7_w42_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_copy828_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid829_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid829_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w42_8_c3 :  std_logic;
signal bh7_w43_6_c3 :  std_logic;
signal bh7_w44_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_copy830_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid831_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid831_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w44_8_c3 :  std_logic;
signal bh7_w45_6_c3 :  std_logic;
signal bh7_w46_7_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_copy832_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid833_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid833_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w46_8_c3 :  std_logic;
signal bh7_w47_6_c3 :  std_logic;
signal bh7_w48_8_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_copy834_c3 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid835_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid835_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w48_9_c3 :  std_logic;
signal bh7_w49_8_c3 :  std_logic;
signal bh7_w50_10_c3 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_copy836_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid837_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid837_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w50_11_c3 :  std_logic;
signal bh7_w51_14_c3 :  std_logic;
signal bh7_w52_15_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_copy838_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid839_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid839_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w52_16_c3 :  std_logic;
signal bh7_w53_18_c3 :  std_logic;
signal bh7_w54_19_c3 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_copy840_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid841_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid841_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3 :  std_logic_vector(2 downto 0);
signal bh7_w54_20_c3 :  std_logic;
signal bh7_w55_21_c3 :  std_logic;
signal bh7_w56_19_c3, bh7_w56_19_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_copy842_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid843_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid843_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w56_20_c4 :  std_logic;
signal bh7_w57_24_c4 :  std_logic;
signal bh7_w58_23_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c3, Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid845_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c0, Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c1, Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c2, Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w58_24_c4 :  std_logic;
signal bh7_w59_21_c4 :  std_logic;
signal bh7_w60_22_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c3, Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid847_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid847_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w59_22_c4 :  std_logic;
signal bh7_w60_23_c4 :  std_logic;
signal bh7_w61_23_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c3, Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid849_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh7_w61_24_c4 :  std_logic;
signal bh7_w62_20_c4 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c3, Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid851_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid851_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w62_21_c4 :  std_logic;
signal bh7_w63_23_c4 :  std_logic;
signal bh7_w64_23_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c3, Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid853_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c0, Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c1, Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c2, Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w63_24_c4 :  std_logic;
signal bh7_w64_24_c4 :  std_logic;
signal bh7_w65_18_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c3, Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid855_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid855_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w64_25_c4 :  std_logic;
signal bh7_w65_19_c4 :  std_logic;
signal bh7_w66_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c3, Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid857_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh7_w66_23_c4 :  std_logic;
signal bh7_w67_20_c4 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c3, Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid859_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid859_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w67_21_c4 :  std_logic;
signal bh7_w68_22_c4 :  std_logic;
signal bh7_w69_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c3, Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid861_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid861_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w69_20_c4 :  std_logic;
signal bh7_w70_22_c4 :  std_logic;
signal bh7_w71_19_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c3, Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid863_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh7_w71_20_c4 :  std_logic;
signal bh7_w72_23_c4 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c3, Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid865_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid865_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w72_24_c4 :  std_logic;
signal bh7_w73_18_c4 :  std_logic;
signal bh7_w74_24_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c3, Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid867_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid867_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w74_25_c4 :  std_logic;
signal bh7_w75_17_c4 :  std_logic;
signal bh7_w76_22_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c3, Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid869_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid869_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w76_23_c4 :  std_logic;
signal bh7_w77_17_c4 :  std_logic;
signal bh7_w78_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c3, Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid871_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid871_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w78_23_c4 :  std_logic;
signal bh7_w79_17_c4 :  std_logic;
signal bh7_w80_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c3, Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid873_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid873_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w80_23_c4 :  std_logic;
signal bh7_w81_17_c4 :  std_logic;
signal bh7_w82_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c3, Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c4 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid875_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_c4 :  std_logic_vector(1 downto 0);
signal bh7_w82_23_c4 :  std_logic;
signal bh7_w83_16_c4 :  std_logic;
signal Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c3, Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c4 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid877_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid877_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w84_21_c4 :  std_logic;
signal bh7_w85_17_c4 :  std_logic;
signal bh7_w86_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c3, Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid879_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid879_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w86_20_c4 :  std_logic;
signal bh7_w87_18_c4 :  std_logic;
signal bh7_w88_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c3, Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid881_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid881_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w88_20_c4 :  std_logic;
signal bh7_w89_16_c4 :  std_logic;
signal bh7_w90_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c3, Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid883_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid883_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w90_20_c4 :  std_logic;
signal bh7_w91_17_c4 :  std_logic;
signal bh7_w92_17_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c3, Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid885_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid885_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w92_18_c4 :  std_logic;
signal bh7_w93_19_c4 :  std_logic;
signal bh7_w94_17_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c3, Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid887_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid887_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w95_17_c4 :  std_logic;
signal bh7_w96_19_c4 :  std_logic;
signal bh7_w97_17_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c3, Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid889_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid889_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w98_17_c4 :  std_logic;
signal bh7_w99_17_c4 :  std_logic;
signal bh7_w100_14_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c3, Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid891_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid891_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w100_15_c4 :  std_logic;
signal bh7_w101_12_c4 :  std_logic;
signal bh7_w102_12_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c3, Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid893_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid893_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w104_7_c4 :  std_logic;
signal bh7_w105_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c3, Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid895_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid895_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w21_6_c4 :  std_logic;
signal bh7_w22_4_c4 :  std_logic;
signal bh7_w23_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c3, Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid897_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid897_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w23_7_c4 :  std_logic;
signal bh7_w24_6_c4 :  std_logic;
signal bh7_w25_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c3, Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid899_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid899_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w25_7_c4 :  std_logic;
signal bh7_w26_6_c4 :  std_logic;
signal bh7_w27_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c3, Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid901_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid901_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w27_7_c4 :  std_logic;
signal bh7_w28_6_c4 :  std_logic;
signal bh7_w29_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c3, Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid903_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid903_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w29_7_c4 :  std_logic;
signal bh7_w30_6_c4 :  std_logic;
signal bh7_w31_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c3, Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid905_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid905_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w31_7_c4 :  std_logic;
signal bh7_w32_6_c4 :  std_logic;
signal bh7_w33_6_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c3, Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid907_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid907_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w33_7_c4 :  std_logic;
signal bh7_w34_7_c4 :  std_logic;
signal bh7_w35_8_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c3, Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid909_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid909_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w35_9_c4 :  std_logic;
signal bh7_w36_9_c4 :  std_logic;
signal bh7_w37_7_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c3, Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid911_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid911_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w38_9_c4 :  std_logic;
signal bh7_w39_7_c4 :  std_logic;
signal bh7_w40_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c3, Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid913_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid913_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w40_10_c4 :  std_logic;
signal bh7_w41_7_c4 :  std_logic;
signal bh7_w42_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c3, Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid915_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid915_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w42_10_c4 :  std_logic;
signal bh7_w43_7_c4 :  std_logic;
signal bh7_w44_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c3, Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid917_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid917_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w44_10_c4 :  std_logic;
signal bh7_w45_7_c4 :  std_logic;
signal bh7_w46_9_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c3, Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid919_In0_c3 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid919_In1_c3 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w46_10_c4 :  std_logic;
signal bh7_w47_7_c4 :  std_logic;
signal bh7_w48_10_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c3, Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid921_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid921_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w48_11_c4 :  std_logic;
signal bh7_w49_9_c4 :  std_logic;
signal bh7_w50_12_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c3, Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid923_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid923_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w50_13_c4 :  std_logic;
signal bh7_w51_15_c4 :  std_logic;
signal bh7_w52_17_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c3, Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid925_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid925_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w52_18_c4 :  std_logic;
signal bh7_w53_19_c4 :  std_logic;
signal bh7_w54_21_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c3, Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid927_In0_c3 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid927_In1_c3 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w54_22_c4 :  std_logic;
signal bh7_w55_22_c4 :  std_logic;
signal bh7_w56_21_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c3, Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid929_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid929_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w56_22_c4 :  std_logic;
signal bh7_w57_25_c4 :  std_logic;
signal bh7_w58_25_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_copy930_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid931_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid931_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w58_26_c4 :  std_logic;
signal bh7_w59_23_c4 :  std_logic;
signal bh7_w60_24_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_copy932_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid933_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid933_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w60_25_c4 :  std_logic;
signal bh7_w61_25_c4 :  std_logic;
signal bh7_w62_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_copy934_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid935_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid935_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w62_23_c4 :  std_logic;
signal bh7_w63_25_c4 :  std_logic;
signal bh7_w64_26_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_copy936_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid937_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid937_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w64_27_c4 :  std_logic;
signal bh7_w65_20_c4 :  std_logic;
signal bh7_w66_24_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_copy938_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid939_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid939_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w66_25_c4 :  std_logic;
signal bh7_w67_22_c4 :  std_logic;
signal bh7_w68_23_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_copy940_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid941_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid941_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w68_24_c4 :  std_logic;
signal bh7_w69_21_c4 :  std_logic;
signal bh7_w70_23_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_copy942_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid943_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid943_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w71_21_c4 :  std_logic;
signal bh7_w72_25_c4 :  std_logic;
signal bh7_w73_19_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_copy944_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid945_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid945_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w73_20_c4 :  std_logic;
signal bh7_w74_26_c4 :  std_logic;
signal bh7_w75_18_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_copy946_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid947_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid947_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w75_19_c4 :  std_logic;
signal bh7_w76_24_c4 :  std_logic;
signal bh7_w77_18_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_copy948_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid949_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid949_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w78_24_c4 :  std_logic;
signal bh7_w79_18_c4 :  std_logic;
signal bh7_w80_24_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_copy950_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid951_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid951_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w80_25_c4 :  std_logic;
signal bh7_w81_18_c4 :  std_logic;
signal bh7_w82_24_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_copy952_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid953_In0_c4 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid953_In1_c4 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w82_25_c4 :  std_logic;
signal bh7_w83_17_c4 :  std_logic;
signal bh7_w84_22_c4 :  std_logic;
signal Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_copy954_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid955_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid955_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w86_21_c4 :  std_logic;
signal bh7_w87_19_c4 :  std_logic;
signal bh7_w88_21_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_copy956_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid957_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid957_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w88_22_c4 :  std_logic;
signal bh7_w89_17_c4 :  std_logic;
signal bh7_w90_21_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_copy958_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid959_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid959_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w90_22_c4 :  std_logic;
signal bh7_w91_18_c4 :  std_logic;
signal bh7_w92_19_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_copy960_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid961_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid961_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w92_20_c4 :  std_logic;
signal bh7_w93_20_c4 :  std_logic;
signal bh7_w94_18_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_copy962_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid963_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid963_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w94_19_c4 :  std_logic;
signal bh7_w95_18_c4 :  std_logic;
signal bh7_w96_20_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_copy964_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid965_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid965_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w97_18_c4 :  std_logic;
signal bh7_w98_18_c4 :  std_logic;
signal bh7_w99_18_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_copy966_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid967_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid967_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w100_16_c4 :  std_logic;
signal bh7_w101_13_c4 :  std_logic;
signal bh7_w102_13_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_copy968_c4 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid969_In0_c4 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c3, Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c4 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4 :  std_logic_vector(2 downto 0);
signal bh7_w102_14_c4 :  std_logic;
signal bh7_w103_11_c4 :  std_logic;
signal bh7_w104_8_c4 :  std_logic;
signal Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_copy970_c4 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh7_22_c4, tmp_bitheapResult_bh7_22_c5, tmp_bitheapResult_bh7_22_c6, tmp_bitheapResult_bh7_22_c7, tmp_bitheapResult_bh7_22_c8, tmp_bitheapResult_bh7_22_c9, tmp_bitheapResult_bh7_22_c10, tmp_bitheapResult_bh7_22_c11, tmp_bitheapResult_bh7_22_c12, tmp_bitheapResult_bh7_22_c13, tmp_bitheapResult_bh7_22_c14, tmp_bitheapResult_bh7_22_c15, tmp_bitheapResult_bh7_22_c16, tmp_bitheapResult_bh7_22_c17, tmp_bitheapResult_bh7_22_c18, tmp_bitheapResult_bh7_22_c19, tmp_bitheapResult_bh7_22_c20, tmp_bitheapResult_bh7_22_c21, tmp_bitheapResult_bh7_22_c22, tmp_bitheapResult_bh7_22_c23, tmp_bitheapResult_bh7_22_c24, tmp_bitheapResult_bh7_22_c25, tmp_bitheapResult_bh7_22_c26, tmp_bitheapResult_bh7_22_c27, tmp_bitheapResult_bh7_22_c28, tmp_bitheapResult_bh7_22_c29, tmp_bitheapResult_bh7_22_c30, tmp_bitheapResult_bh7_22_c31, tmp_bitheapResult_bh7_22_c32, tmp_bitheapResult_bh7_22_c33 :  std_logic_vector(22 downto 0);
signal bitheapFinalAdd_bh7_In0_c4 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_In1_c4 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh7_Out_c33 :  std_logic_vector(83 downto 0);
signal bitheapResult_bh7_c33 :  std_logic_vector(105 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               bh7_w62_8_c1 <= bh7_w62_8_c0;
               bh7_w59_8_c1 <= bh7_w59_8_c0;
               bh7_w56_8_c1 <= bh7_w56_8_c0;
               bh7_w48_4_c1 <= bh7_w48_4_c0;
               bh7_w66_9_c1 <= bh7_w66_9_c0;
               bh7_w97_7_c1 <= bh7_w97_7_c0;
               bh7_w94_7_c1 <= bh7_w94_7_c0;
               bh7_w91_7_c1 <= bh7_w91_7_c0;
               bh7_w88_7_c1 <= bh7_w88_7_c0;
               bh7_w82_7_c1 <= bh7_w82_7_c0;
               bh7_w85_7_c1 <= bh7_w85_7_c0;
               bh7_w104_0_c1 <= bh7_w104_0_c0;
               bh7_w105_0_c1 <= bh7_w105_0_c0;
               bh7_w103_1_c1 <= bh7_w103_1_c0;
               Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c0;
               Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c0;
               Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c0;
               Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c0;
               Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c0;
               Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c0;
            end if;
            if ce_2 = '1' then
               bh7_w48_4_c2 <= bh7_w48_4_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c1;
               Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c1;
               Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c1;
               Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c1;
            end if;
            if ce_3 = '1' then
               bh7_w0_0_c3 <= bh7_w0_0_c2;
               bh7_w1_0_c3 <= bh7_w1_0_c2;
               bh7_w2_0_c3 <= bh7_w2_0_c2;
               bh7_w3_0_c3 <= bh7_w3_0_c2;
               bh7_w4_0_c3 <= bh7_w4_0_c2;
               bh7_w5_0_c3 <= bh7_w5_0_c2;
               bh7_w6_0_c3 <= bh7_w6_0_c2;
               bh7_w7_0_c3 <= bh7_w7_0_c2;
               bh7_w8_0_c3 <= bh7_w8_0_c2;
               bh7_w9_0_c3 <= bh7_w9_0_c2;
               bh7_w10_0_c3 <= bh7_w10_0_c2;
               bh7_w11_0_c3 <= bh7_w11_0_c2;
               bh7_w12_0_c3 <= bh7_w12_0_c2;
               bh7_w13_0_c3 <= bh7_w13_0_c2;
               bh7_w14_0_c3 <= bh7_w14_0_c2;
               bh7_w15_0_c3 <= bh7_w15_0_c2;
               bh7_w16_0_c3 <= bh7_w16_0_c2;
               bh7_w59_0_c3 <= bh7_w59_0_c2;
               bh7_w60_0_c3 <= bh7_w60_0_c2;
               bh7_w61_0_c3 <= bh7_w61_0_c2;
               bh7_w62_0_c3 <= bh7_w62_0_c2;
               bh7_w64_0_c3 <= bh7_w64_0_c2;
               bh7_w65_0_c3 <= bh7_w65_0_c2;
               bh7_w67_0_c3 <= bh7_w67_0_c2;
               bh7_w69_0_c3 <= bh7_w69_0_c2;
               bh7_w70_0_c3 <= bh7_w70_0_c2;
               bh7_w72_0_c3 <= bh7_w72_0_c2;
               bh7_w74_0_c3 <= bh7_w74_0_c2;
               bh7_w25_2_c3 <= bh7_w25_2_c2;
               bh7_w27_2_c3 <= bh7_w27_2_c2;
               bh7_w29_2_c3 <= bh7_w29_2_c2;
               bh7_w31_2_c3 <= bh7_w31_2_c2;
               bh7_w33_2_c3 <= bh7_w33_2_c2;
               bh7_w59_2_c3 <= bh7_w59_2_c2;
               bh7_w60_3_c3 <= bh7_w60_3_c2;
               bh7_w61_3_c3 <= bh7_w61_3_c2;
               bh7_w62_2_c3 <= bh7_w62_2_c2;
               bh7_w64_3_c3 <= bh7_w64_3_c2;
               bh7_w48_3_c3 <= bh7_w48_3_c2;
               bh7_w59_3_c3 <= bh7_w59_3_c2;
               bh7_w60_4_c3 <= bh7_w60_4_c2;
               bh7_w61_4_c3 <= bh7_w61_4_c2;
               bh7_w62_3_c3 <= bh7_w62_3_c2;
               bh7_w64_4_c3 <= bh7_w64_4_c2;
               bh7_w65_2_c3 <= bh7_w65_2_c2;
               bh7_w67_3_c3 <= bh7_w67_3_c2;
               bh7_w69_3_c3 <= bh7_w69_3_c2;
               bh7_w70_3_c3 <= bh7_w70_3_c2;
               bh7_w72_3_c3 <= bh7_w72_3_c2;
               bh7_w74_2_c3 <= bh7_w74_2_c2;
               bh7_w76_1_c3 <= bh7_w76_1_c2;
               bh7_w77_0_c3 <= bh7_w77_0_c2;
               bh7_w78_0_c3 <= bh7_w78_0_c2;
               bh7_w79_0_c3 <= bh7_w79_0_c2;
               bh7_w80_0_c3 <= bh7_w80_0_c2;
               bh7_w81_0_c3 <= bh7_w81_0_c2;
               bh7_w58_5_c3 <= bh7_w58_5_c2;
               bh7_w59_4_c3 <= bh7_w59_4_c2;
               bh7_w60_5_c3 <= bh7_w60_5_c2;
               bh7_w61_5_c3 <= bh7_w61_5_c2;
               bh7_w62_4_c3 <= bh7_w62_4_c2;
               bh7_w63_5_c3 <= bh7_w63_5_c2;
               bh7_w64_5_c3 <= bh7_w64_5_c2;
               bh7_w65_3_c3 <= bh7_w65_3_c2;
               bh7_w67_4_c3 <= bh7_w67_4_c2;
               bh7_w69_4_c3 <= bh7_w69_4_c2;
               bh7_w70_4_c3 <= bh7_w70_4_c2;
               bh7_w72_4_c3 <= bh7_w72_4_c2;
               bh7_w74_3_c3 <= bh7_w74_3_c2;
               bh7_w75_2_c3 <= bh7_w75_2_c2;
               bh7_w76_2_c3 <= bh7_w76_2_c2;
               bh7_w77_1_c3 <= bh7_w77_1_c2;
               bh7_w78_1_c3 <= bh7_w78_1_c2;
               bh7_w79_1_c3 <= bh7_w79_1_c2;
               bh7_w80_1_c3 <= bh7_w80_1_c2;
               bh7_w81_1_c3 <= bh7_w81_1_c2;
               bh7_w82_0_c3 <= bh7_w82_0_c2;
               bh7_w83_0_c3 <= bh7_w83_0_c2;
               bh7_w84_0_c3 <= bh7_w84_0_c2;
               bh7_w85_0_c3 <= bh7_w85_0_c2;
               bh7_w86_0_c3 <= bh7_w86_0_c2;
               bh7_w87_0_c3 <= bh7_w87_0_c2;
               bh7_w88_0_c3 <= bh7_w88_0_c2;
               bh7_w89_0_c3 <= bh7_w89_0_c2;
               bh7_w90_0_c3 <= bh7_w90_0_c2;
               bh7_w91_0_c3 <= bh7_w91_0_c2;
               bh7_w92_0_c3 <= bh7_w92_0_c2;
               bh7_w93_0_c3 <= bh7_w93_0_c2;
               bh7_w94_0_c3 <= bh7_w94_0_c2;
               bh7_w95_0_c3 <= bh7_w95_0_c2;
               bh7_w96_0_c3 <= bh7_w96_0_c2;
               bh7_w97_0_c3 <= bh7_w97_0_c2;
               bh7_w98_0_c3 <= bh7_w98_0_c2;
               bh7_w61_18_c3 <= bh7_w61_18_c2;
               bh7_w64_18_c3 <= bh7_w64_18_c2;
               bh7_w67_15_c3 <= bh7_w67_15_c2;
               bh7_w90_15_c3 <= bh7_w90_15_c2;
               bh7_w93_15_c3 <= bh7_w93_15_c2;
               bh7_w96_15_c3 <= bh7_w96_15_c2;
               bh7_w99_14_c3 <= bh7_w99_14_c2;
               bh7_w102_9_c3 <= bh7_w102_9_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c2;
               Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c2;
               Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c2;
               Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c2;
            end if;
            if ce_4 = '1' then
               bh7_w0_0_c4 <= bh7_w0_0_c3;
               bh7_w1_0_c4 <= bh7_w1_0_c3;
               bh7_w2_0_c4 <= bh7_w2_0_c3;
               bh7_w3_0_c4 <= bh7_w3_0_c3;
               bh7_w4_0_c4 <= bh7_w4_0_c3;
               bh7_w5_0_c4 <= bh7_w5_0_c3;
               bh7_w6_0_c4 <= bh7_w6_0_c3;
               bh7_w7_0_c4 <= bh7_w7_0_c3;
               bh7_w8_0_c4 <= bh7_w8_0_c3;
               bh7_w9_0_c4 <= bh7_w9_0_c3;
               bh7_w10_0_c4 <= bh7_w10_0_c3;
               bh7_w11_0_c4 <= bh7_w11_0_c3;
               bh7_w12_0_c4 <= bh7_w12_0_c3;
               bh7_w13_0_c4 <= bh7_w13_0_c3;
               bh7_w14_0_c4 <= bh7_w14_0_c3;
               bh7_w15_0_c4 <= bh7_w15_0_c3;
               bh7_w16_0_c4 <= bh7_w16_0_c3;
               bh7_w17_2_c4 <= bh7_w17_2_c3;
               bh7_w18_2_c4 <= bh7_w18_2_c3;
               bh7_w57_23_c4 <= bh7_w57_23_c3;
               bh7_w68_21_c4 <= bh7_w68_21_c3;
               bh7_w73_17_c4 <= bh7_w73_17_c3;
               bh7_w75_16_c4 <= bh7_w75_16_c3;
               bh7_w83_15_c4 <= bh7_w83_15_c3;
               bh7_w94_16_c4 <= bh7_w94_16_c3;
               bh7_w97_16_c4 <= bh7_w97_16_c3;
               bh7_w102_11_c4 <= bh7_w102_11_c3;
               bh7_w19_4_c4 <= bh7_w19_4_c3;
               bh7_w20_3_c4 <= bh7_w20_3_c3;
               bh7_w37_6_c4 <= bh7_w37_6_c3;
               bh7_w56_19_c4 <= bh7_w56_19_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c3;
               Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c3;
               Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c3;
               Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c3;
               Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c3;
               Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c3;
               Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c3;
            end if;
            if ce_5 = '1' then
               tmp_bitheapResult_bh7_22_c5 <= tmp_bitheapResult_bh7_22_c4;
            end if;
            if ce_6 = '1' then
               tmp_bitheapResult_bh7_22_c6 <= tmp_bitheapResult_bh7_22_c5;
            end if;
            if ce_7 = '1' then
               tmp_bitheapResult_bh7_22_c7 <= tmp_bitheapResult_bh7_22_c6;
            end if;
            if ce_8 = '1' then
               tmp_bitheapResult_bh7_22_c8 <= tmp_bitheapResult_bh7_22_c7;
            end if;
            if ce_9 = '1' then
               tmp_bitheapResult_bh7_22_c9 <= tmp_bitheapResult_bh7_22_c8;
            end if;
            if ce_10 = '1' then
               tmp_bitheapResult_bh7_22_c10 <= tmp_bitheapResult_bh7_22_c9;
            end if;
            if ce_11 = '1' then
               tmp_bitheapResult_bh7_22_c11 <= tmp_bitheapResult_bh7_22_c10;
            end if;
            if ce_12 = '1' then
               tmp_bitheapResult_bh7_22_c12 <= tmp_bitheapResult_bh7_22_c11;
            end if;
            if ce_13 = '1' then
               tmp_bitheapResult_bh7_22_c13 <= tmp_bitheapResult_bh7_22_c12;
            end if;
            if ce_14 = '1' then
               tmp_bitheapResult_bh7_22_c14 <= tmp_bitheapResult_bh7_22_c13;
            end if;
            if ce_15 = '1' then
               tmp_bitheapResult_bh7_22_c15 <= tmp_bitheapResult_bh7_22_c14;
            end if;
            if ce_16 = '1' then
               tmp_bitheapResult_bh7_22_c16 <= tmp_bitheapResult_bh7_22_c15;
            end if;
            if ce_17 = '1' then
               tmp_bitheapResult_bh7_22_c17 <= tmp_bitheapResult_bh7_22_c16;
            end if;
            if ce_18 = '1' then
               tmp_bitheapResult_bh7_22_c18 <= tmp_bitheapResult_bh7_22_c17;
            end if;
            if ce_19 = '1' then
               tmp_bitheapResult_bh7_22_c19 <= tmp_bitheapResult_bh7_22_c18;
            end if;
            if ce_20 = '1' then
               tmp_bitheapResult_bh7_22_c20 <= tmp_bitheapResult_bh7_22_c19;
            end if;
            if ce_21 = '1' then
               tmp_bitheapResult_bh7_22_c21 <= tmp_bitheapResult_bh7_22_c20;
            end if;
            if ce_22 = '1' then
               tmp_bitheapResult_bh7_22_c22 <= tmp_bitheapResult_bh7_22_c21;
            end if;
            if ce_23 = '1' then
               tmp_bitheapResult_bh7_22_c23 <= tmp_bitheapResult_bh7_22_c22;
            end if;
            if ce_24 = '1' then
               tmp_bitheapResult_bh7_22_c24 <= tmp_bitheapResult_bh7_22_c23;
            end if;
            if ce_25 = '1' then
               tmp_bitheapResult_bh7_22_c25 <= tmp_bitheapResult_bh7_22_c24;
            end if;
            if ce_26 = '1' then
               tmp_bitheapResult_bh7_22_c26 <= tmp_bitheapResult_bh7_22_c25;
            end if;
            if ce_27 = '1' then
               tmp_bitheapResult_bh7_22_c27 <= tmp_bitheapResult_bh7_22_c26;
            end if;
            if ce_28 = '1' then
               tmp_bitheapResult_bh7_22_c28 <= tmp_bitheapResult_bh7_22_c27;
            end if;
            if ce_29 = '1' then
               tmp_bitheapResult_bh7_22_c29 <= tmp_bitheapResult_bh7_22_c28;
            end if;
            if ce_30 = '1' then
               tmp_bitheapResult_bh7_22_c30 <= tmp_bitheapResult_bh7_22_c29;
            end if;
            if ce_31 = '1' then
               tmp_bitheapResult_bh7_22_c31 <= tmp_bitheapResult_bh7_22_c30;
            end if;
            if ce_32 = '1' then
               tmp_bitheapResult_bh7_22_c32 <= tmp_bitheapResult_bh7_22_c31;
            end if;
            if ce_33 = '1' then
               tmp_bitheapResult_bh7_22_c33 <= tmp_bitheapResult_bh7_22_c32;
            end if;
         end if;
      end process;
   XX_m6_c0 <= X ;
   YY_m6_c0 <= Y ;
   tile_0_X_c0 <= X(16 downto 0);
   tile_0_Y_c0 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq800_uid9
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_0_X_c0,
                 Y => tile_0_Y_c0,
                 R => tile_0_output_c2);

   tile_0_filtered_output_c2 <= unsigned(tile_0_output_c2(40 downto 0));
   bh7_w0_0_c2 <= tile_0_filtered_output_c2(0);
   bh7_w1_0_c2 <= tile_0_filtered_output_c2(1);
   bh7_w2_0_c2 <= tile_0_filtered_output_c2(2);
   bh7_w3_0_c2 <= tile_0_filtered_output_c2(3);
   bh7_w4_0_c2 <= tile_0_filtered_output_c2(4);
   bh7_w5_0_c2 <= tile_0_filtered_output_c2(5);
   bh7_w6_0_c2 <= tile_0_filtered_output_c2(6);
   bh7_w7_0_c2 <= tile_0_filtered_output_c2(7);
   bh7_w8_0_c2 <= tile_0_filtered_output_c2(8);
   bh7_w9_0_c2 <= tile_0_filtered_output_c2(9);
   bh7_w10_0_c2 <= tile_0_filtered_output_c2(10);
   bh7_w11_0_c2 <= tile_0_filtered_output_c2(11);
   bh7_w12_0_c2 <= tile_0_filtered_output_c2(12);
   bh7_w13_0_c2 <= tile_0_filtered_output_c2(13);
   bh7_w14_0_c2 <= tile_0_filtered_output_c2(14);
   bh7_w15_0_c2 <= tile_0_filtered_output_c2(15);
   bh7_w16_0_c2 <= tile_0_filtered_output_c2(16);
   bh7_w17_0_c2 <= tile_0_filtered_output_c2(17);
   bh7_w18_0_c2 <= tile_0_filtered_output_c2(18);
   bh7_w19_0_c2 <= tile_0_filtered_output_c2(19);
   bh7_w20_0_c2 <= tile_0_filtered_output_c2(20);
   bh7_w21_0_c2 <= tile_0_filtered_output_c2(21);
   bh7_w22_0_c2 <= tile_0_filtered_output_c2(22);
   bh7_w23_0_c2 <= tile_0_filtered_output_c2(23);
   bh7_w24_0_c2 <= tile_0_filtered_output_c2(24);
   bh7_w25_0_c2 <= tile_0_filtered_output_c2(25);
   bh7_w26_0_c2 <= tile_0_filtered_output_c2(26);
   bh7_w27_0_c2 <= tile_0_filtered_output_c2(27);
   bh7_w28_0_c2 <= tile_0_filtered_output_c2(28);
   bh7_w29_0_c2 <= tile_0_filtered_output_c2(29);
   bh7_w30_0_c2 <= tile_0_filtered_output_c2(30);
   bh7_w31_0_c2 <= tile_0_filtered_output_c2(31);
   bh7_w32_0_c2 <= tile_0_filtered_output_c2(32);
   bh7_w33_0_c2 <= tile_0_filtered_output_c2(33);
   bh7_w34_0_c2 <= tile_0_filtered_output_c2(34);
   bh7_w35_0_c2 <= tile_0_filtered_output_c2(35);
   bh7_w36_0_c2 <= tile_0_filtered_output_c2(36);
   bh7_w37_0_c2 <= tile_0_filtered_output_c2(37);
   bh7_w38_0_c2 <= tile_0_filtered_output_c2(38);
   bh7_w39_0_c2 <= tile_0_filtered_output_c2(39);
   bh7_w40_0_c2 <= tile_0_filtered_output_c2(40);
   tile_1_X_c0 <= X(33 downto 17);
   tile_1_Y_c0 <= Y(23 downto 0);
   tile_1_mult: DSPBlock_17x24_Freq800_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_1_X_c0,
                 Y => tile_1_Y_c0,
                 R => tile_1_output_c2);

   tile_1_filtered_output_c2 <= unsigned(tile_1_output_c2(40 downto 0));
   bh7_w17_1_c2 <= tile_1_filtered_output_c2(0);
   bh7_w18_1_c2 <= tile_1_filtered_output_c2(1);
   bh7_w19_1_c2 <= tile_1_filtered_output_c2(2);
   bh7_w20_1_c2 <= tile_1_filtered_output_c2(3);
   bh7_w21_1_c2 <= tile_1_filtered_output_c2(4);
   bh7_w22_1_c2 <= tile_1_filtered_output_c2(5);
   bh7_w23_1_c2 <= tile_1_filtered_output_c2(6);
   bh7_w24_1_c2 <= tile_1_filtered_output_c2(7);
   bh7_w25_1_c2 <= tile_1_filtered_output_c2(8);
   bh7_w26_1_c2 <= tile_1_filtered_output_c2(9);
   bh7_w27_1_c2 <= tile_1_filtered_output_c2(10);
   bh7_w28_1_c2 <= tile_1_filtered_output_c2(11);
   bh7_w29_1_c2 <= tile_1_filtered_output_c2(12);
   bh7_w30_1_c2 <= tile_1_filtered_output_c2(13);
   bh7_w31_1_c2 <= tile_1_filtered_output_c2(14);
   bh7_w32_1_c2 <= tile_1_filtered_output_c2(15);
   bh7_w33_1_c2 <= tile_1_filtered_output_c2(16);
   bh7_w34_1_c2 <= tile_1_filtered_output_c2(17);
   bh7_w35_1_c2 <= tile_1_filtered_output_c2(18);
   bh7_w36_1_c2 <= tile_1_filtered_output_c2(19);
   bh7_w37_1_c2 <= tile_1_filtered_output_c2(20);
   bh7_w38_1_c2 <= tile_1_filtered_output_c2(21);
   bh7_w39_1_c2 <= tile_1_filtered_output_c2(22);
   bh7_w40_1_c2 <= tile_1_filtered_output_c2(23);
   bh7_w41_0_c2 <= tile_1_filtered_output_c2(24);
   bh7_w42_0_c2 <= tile_1_filtered_output_c2(25);
   bh7_w43_0_c2 <= tile_1_filtered_output_c2(26);
   bh7_w44_0_c2 <= tile_1_filtered_output_c2(27);
   bh7_w45_0_c2 <= tile_1_filtered_output_c2(28);
   bh7_w46_0_c2 <= tile_1_filtered_output_c2(29);
   bh7_w47_0_c2 <= tile_1_filtered_output_c2(30);
   bh7_w48_0_c2 <= tile_1_filtered_output_c2(31);
   bh7_w49_0_c2 <= tile_1_filtered_output_c2(32);
   bh7_w50_0_c2 <= tile_1_filtered_output_c2(33);
   bh7_w51_0_c2 <= tile_1_filtered_output_c2(34);
   bh7_w52_0_c2 <= tile_1_filtered_output_c2(35);
   bh7_w53_0_c2 <= tile_1_filtered_output_c2(36);
   bh7_w54_0_c2 <= tile_1_filtered_output_c2(37);
   bh7_w55_0_c2 <= tile_1_filtered_output_c2(38);
   bh7_w56_0_c2 <= tile_1_filtered_output_c2(39);
   bh7_w57_0_c2 <= tile_1_filtered_output_c2(40);
   tile_2_X_c0 <= X(50 downto 34);
   tile_2_Y_c0 <= Y(23 downto 0);
   tile_2_mult: DSPBlock_17x24_Freq800_uid13
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_2_X_c0,
                 Y => tile_2_Y_c0,
                 R => tile_2_output_c2);

   tile_2_filtered_output_c2 <= unsigned(tile_2_output_c2(40 downto 0));
   bh7_w34_2_c2 <= tile_2_filtered_output_c2(0);
   bh7_w35_2_c2 <= tile_2_filtered_output_c2(1);
   bh7_w36_2_c2 <= tile_2_filtered_output_c2(2);
   bh7_w37_2_c2 <= tile_2_filtered_output_c2(3);
   bh7_w38_2_c2 <= tile_2_filtered_output_c2(4);
   bh7_w39_2_c2 <= tile_2_filtered_output_c2(5);
   bh7_w40_2_c2 <= tile_2_filtered_output_c2(6);
   bh7_w41_1_c2 <= tile_2_filtered_output_c2(7);
   bh7_w42_1_c2 <= tile_2_filtered_output_c2(8);
   bh7_w43_1_c2 <= tile_2_filtered_output_c2(9);
   bh7_w44_1_c2 <= tile_2_filtered_output_c2(10);
   bh7_w45_1_c2 <= tile_2_filtered_output_c2(11);
   bh7_w46_1_c2 <= tile_2_filtered_output_c2(12);
   bh7_w47_1_c2 <= tile_2_filtered_output_c2(13);
   bh7_w48_1_c2 <= tile_2_filtered_output_c2(14);
   bh7_w49_1_c2 <= tile_2_filtered_output_c2(15);
   bh7_w50_1_c2 <= tile_2_filtered_output_c2(16);
   bh7_w51_1_c2 <= tile_2_filtered_output_c2(17);
   bh7_w52_1_c2 <= tile_2_filtered_output_c2(18);
   bh7_w53_1_c2 <= tile_2_filtered_output_c2(19);
   bh7_w54_1_c2 <= tile_2_filtered_output_c2(20);
   bh7_w55_1_c2 <= tile_2_filtered_output_c2(21);
   bh7_w56_1_c2 <= tile_2_filtered_output_c2(22);
   bh7_w57_1_c2 <= tile_2_filtered_output_c2(23);
   bh7_w58_0_c2 <= tile_2_filtered_output_c2(24);
   bh7_w59_0_c2 <= tile_2_filtered_output_c2(25);
   bh7_w60_0_c2 <= tile_2_filtered_output_c2(26);
   bh7_w61_0_c2 <= tile_2_filtered_output_c2(27);
   bh7_w62_0_c2 <= tile_2_filtered_output_c2(28);
   bh7_w63_0_c2 <= tile_2_filtered_output_c2(29);
   bh7_w64_0_c2 <= tile_2_filtered_output_c2(30);
   bh7_w65_0_c2 <= tile_2_filtered_output_c2(31);
   bh7_w66_0_c2 <= tile_2_filtered_output_c2(32);
   bh7_w67_0_c2 <= tile_2_filtered_output_c2(33);
   bh7_w68_0_c2 <= tile_2_filtered_output_c2(34);
   bh7_w69_0_c2 <= tile_2_filtered_output_c2(35);
   bh7_w70_0_c2 <= tile_2_filtered_output_c2(36);
   bh7_w71_0_c2 <= tile_2_filtered_output_c2(37);
   bh7_w72_0_c2 <= tile_2_filtered_output_c2(38);
   bh7_w73_0_c2 <= tile_2_filtered_output_c2(39);
   bh7_w74_0_c2 <= tile_2_filtered_output_c2(40);
   tile_3_X_c0 <= X(52 downto 51);
   tile_3_Y_c0 <= Y(23 downto 21);
   tile_3_mult: IntMultiplierLUT_2x3_Freq800_uid15
      port map ( clk  => clk,
                 X => tile_3_X_c0,
                 Y => tile_3_Y_c0,
                 R => tile_3_output_c0);

   tile_3_filtered_output_c0 <= unsigned(tile_3_output_c0(4 downto 0));
   bh7_w72_1_c0 <= tile_3_filtered_output_c0(0);
   bh7_w73_1_c0 <= tile_3_filtered_output_c0(1);
   bh7_w74_1_c0 <= tile_3_filtered_output_c0(2);
   bh7_w75_0_c0 <= tile_3_filtered_output_c0(3);
   bh7_w76_0_c0 <= tile_3_filtered_output_c0(4);
   tile_4_X_c0 <= X(52 downto 51);
   tile_4_Y_c0 <= Y(20 downto 18);
   tile_4_mult: IntMultiplierLUT_2x3_Freq800_uid20
      port map ( clk  => clk,
                 X => tile_4_X_c0,
                 Y => tile_4_Y_c0,
                 R => tile_4_output_c0);

   tile_4_filtered_output_c0 <= unsigned(tile_4_output_c0(4 downto 0));
   bh7_w69_1_c0 <= tile_4_filtered_output_c0(0);
   bh7_w70_1_c0 <= tile_4_filtered_output_c0(1);
   bh7_w71_1_c0 <= tile_4_filtered_output_c0(2);
   bh7_w72_2_c0 <= tile_4_filtered_output_c0(3);
   bh7_w73_2_c0 <= tile_4_filtered_output_c0(4);
   tile_5_X_c0 <= X(52 downto 51);
   tile_5_Y_c0 <= Y(17 downto 15);
   tile_5_mult: IntMultiplierLUT_2x3_Freq800_uid25
      port map ( clk  => clk,
                 X => tile_5_X_c0,
                 Y => tile_5_Y_c0,
                 R => tile_5_output_c0);

   tile_5_filtered_output_c0 <= unsigned(tile_5_output_c0(4 downto 0));
   bh7_w66_1_c0 <= tile_5_filtered_output_c0(0);
   bh7_w67_1_c0 <= tile_5_filtered_output_c0(1);
   bh7_w68_1_c0 <= tile_5_filtered_output_c0(2);
   bh7_w69_2_c0 <= tile_5_filtered_output_c0(3);
   bh7_w70_2_c0 <= tile_5_filtered_output_c0(4);
   tile_6_X_c0 <= X(52 downto 51);
   tile_6_Y_c0 <= Y(14 downto 12);
   tile_6_mult: IntMultiplierLUT_2x3_Freq800_uid30
      port map ( clk  => clk,
                 X => tile_6_X_c0,
                 Y => tile_6_Y_c0,
                 R => tile_6_output_c0);

   tile_6_filtered_output_c0 <= unsigned(tile_6_output_c0(4 downto 0));
   bh7_w63_1_c0 <= tile_6_filtered_output_c0(0);
   bh7_w64_1_c0 <= tile_6_filtered_output_c0(1);
   bh7_w65_1_c0 <= tile_6_filtered_output_c0(2);
   bh7_w66_2_c0 <= tile_6_filtered_output_c0(3);
   bh7_w67_2_c0 <= tile_6_filtered_output_c0(4);
   tile_7_X_c0 <= X(52 downto 51);
   tile_7_Y_c0 <= Y(11 downto 9);
   tile_7_mult: IntMultiplierLUT_2x3_Freq800_uid35
      port map ( clk  => clk,
                 X => tile_7_X_c0,
                 Y => tile_7_Y_c0,
                 R => tile_7_output_c0);

   tile_7_filtered_output_c0 <= unsigned(tile_7_output_c0(4 downto 0));
   bh7_w60_1_c0 <= tile_7_filtered_output_c0(0);
   bh7_w61_1_c0 <= tile_7_filtered_output_c0(1);
   bh7_w62_1_c0 <= tile_7_filtered_output_c0(2);
   bh7_w63_2_c0 <= tile_7_filtered_output_c0(3);
   bh7_w64_2_c0 <= tile_7_filtered_output_c0(4);
   tile_8_X_c0 <= X(52 downto 51);
   tile_8_Y_c0 <= Y(8 downto 6);
   tile_8_mult: IntMultiplierLUT_2x3_Freq800_uid40
      port map ( clk  => clk,
                 X => tile_8_X_c0,
                 Y => tile_8_Y_c0,
                 R => tile_8_output_c0);

   tile_8_filtered_output_c0 <= unsigned(tile_8_output_c0(4 downto 0));
   bh7_w57_2_c0 <= tile_8_filtered_output_c0(0);
   bh7_w58_1_c0 <= tile_8_filtered_output_c0(1);
   bh7_w59_1_c0 <= tile_8_filtered_output_c0(2);
   bh7_w60_2_c0 <= tile_8_filtered_output_c0(3);
   bh7_w61_2_c0 <= tile_8_filtered_output_c0(4);
   tile_9_X_c0 <= X(52 downto 51);
   tile_9_Y_c0 <= Y(5 downto 3);
   tile_9_mult: IntMultiplierLUT_2x3_Freq800_uid45
      port map ( clk  => clk,
                 X => tile_9_X_c0,
                 Y => tile_9_Y_c0,
                 R => tile_9_output_c0);

   tile_9_filtered_output_c0 <= unsigned(tile_9_output_c0(4 downto 0));
   bh7_w54_2_c0 <= tile_9_filtered_output_c0(0);
   bh7_w55_2_c0 <= tile_9_filtered_output_c0(1);
   bh7_w56_2_c0 <= tile_9_filtered_output_c0(2);
   bh7_w57_3_c0 <= tile_9_filtered_output_c0(3);
   bh7_w58_2_c0 <= tile_9_filtered_output_c0(4);
   tile_10_X_c0 <= X(52 downto 51);
   tile_10_Y_c0 <= Y(2 downto 0);
   tile_10_mult: IntMultiplierLUT_2x3_Freq800_uid50
      port map ( clk  => clk,
                 X => tile_10_X_c0,
                 Y => tile_10_Y_c0,
                 R => tile_10_output_c0);

   tile_10_filtered_output_c0 <= unsigned(tile_10_output_c0(4 downto 0));
   bh7_w51_2_c0 <= tile_10_filtered_output_c0(0);
   bh7_w52_2_c0 <= tile_10_filtered_output_c0(1);
   bh7_w53_2_c0 <= tile_10_filtered_output_c0(2);
   bh7_w54_3_c0 <= tile_10_filtered_output_c0(3);
   bh7_w55_3_c0 <= tile_10_filtered_output_c0(4);
   tile_11_X_c0 <= X(16 downto 0);
   tile_11_Y_c0 <= Y(47 downto 24);
   tile_11_mult: DSPBlock_17x24_Freq800_uid55
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_11_X_c0,
                 Y => tile_11_Y_c0,
                 R => tile_11_output_c2);

   tile_11_filtered_output_c2 <= unsigned(tile_11_output_c2(40 downto 0));
   bh7_w24_2_c2 <= tile_11_filtered_output_c2(0);
   bh7_w25_2_c2 <= tile_11_filtered_output_c2(1);
   bh7_w26_2_c2 <= tile_11_filtered_output_c2(2);
   bh7_w27_2_c2 <= tile_11_filtered_output_c2(3);
   bh7_w28_2_c2 <= tile_11_filtered_output_c2(4);
   bh7_w29_2_c2 <= tile_11_filtered_output_c2(5);
   bh7_w30_2_c2 <= tile_11_filtered_output_c2(6);
   bh7_w31_2_c2 <= tile_11_filtered_output_c2(7);
   bh7_w32_2_c2 <= tile_11_filtered_output_c2(8);
   bh7_w33_2_c2 <= tile_11_filtered_output_c2(9);
   bh7_w34_3_c2 <= tile_11_filtered_output_c2(10);
   bh7_w35_3_c2 <= tile_11_filtered_output_c2(11);
   bh7_w36_3_c2 <= tile_11_filtered_output_c2(12);
   bh7_w37_3_c2 <= tile_11_filtered_output_c2(13);
   bh7_w38_3_c2 <= tile_11_filtered_output_c2(14);
   bh7_w39_3_c2 <= tile_11_filtered_output_c2(15);
   bh7_w40_3_c2 <= tile_11_filtered_output_c2(16);
   bh7_w41_2_c2 <= tile_11_filtered_output_c2(17);
   bh7_w42_2_c2 <= tile_11_filtered_output_c2(18);
   bh7_w43_2_c2 <= tile_11_filtered_output_c2(19);
   bh7_w44_2_c2 <= tile_11_filtered_output_c2(20);
   bh7_w45_2_c2 <= tile_11_filtered_output_c2(21);
   bh7_w46_2_c2 <= tile_11_filtered_output_c2(22);
   bh7_w47_2_c2 <= tile_11_filtered_output_c2(23);
   bh7_w48_2_c2 <= tile_11_filtered_output_c2(24);
   bh7_w49_2_c2 <= tile_11_filtered_output_c2(25);
   bh7_w50_2_c2 <= tile_11_filtered_output_c2(26);
   bh7_w51_3_c2 <= tile_11_filtered_output_c2(27);
   bh7_w52_3_c2 <= tile_11_filtered_output_c2(28);
   bh7_w53_3_c2 <= tile_11_filtered_output_c2(29);
   bh7_w54_4_c2 <= tile_11_filtered_output_c2(30);
   bh7_w55_4_c2 <= tile_11_filtered_output_c2(31);
   bh7_w56_3_c2 <= tile_11_filtered_output_c2(32);
   bh7_w57_4_c2 <= tile_11_filtered_output_c2(33);
   bh7_w58_3_c2 <= tile_11_filtered_output_c2(34);
   bh7_w59_2_c2 <= tile_11_filtered_output_c2(35);
   bh7_w60_3_c2 <= tile_11_filtered_output_c2(36);
   bh7_w61_3_c2 <= tile_11_filtered_output_c2(37);
   bh7_w62_2_c2 <= tile_11_filtered_output_c2(38);
   bh7_w63_3_c2 <= tile_11_filtered_output_c2(39);
   bh7_w64_3_c2 <= tile_11_filtered_output_c2(40);
   tile_12_X_c0 <= X(33 downto 17);
   tile_12_Y_c0 <= Y(47 downto 24);
   tile_12_mult: DSPBlock_17x24_Freq800_uid57
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_12_X_c0,
                 Y => tile_12_Y_c0,
                 R => tile_12_output_c2);

   tile_12_filtered_output_c2 <= unsigned(tile_12_output_c2(40 downto 0));
   bh7_w41_3_c2 <= tile_12_filtered_output_c2(0);
   bh7_w42_3_c2 <= tile_12_filtered_output_c2(1);
   bh7_w43_3_c2 <= tile_12_filtered_output_c2(2);
   bh7_w44_3_c2 <= tile_12_filtered_output_c2(3);
   bh7_w45_3_c2 <= tile_12_filtered_output_c2(4);
   bh7_w46_3_c2 <= tile_12_filtered_output_c2(5);
   bh7_w47_3_c2 <= tile_12_filtered_output_c2(6);
   bh7_w48_3_c2 <= tile_12_filtered_output_c2(7);
   bh7_w49_3_c2 <= tile_12_filtered_output_c2(8);
   bh7_w50_3_c2 <= tile_12_filtered_output_c2(9);
   bh7_w51_4_c2 <= tile_12_filtered_output_c2(10);
   bh7_w52_4_c2 <= tile_12_filtered_output_c2(11);
   bh7_w53_4_c2 <= tile_12_filtered_output_c2(12);
   bh7_w54_5_c2 <= tile_12_filtered_output_c2(13);
   bh7_w55_5_c2 <= tile_12_filtered_output_c2(14);
   bh7_w56_4_c2 <= tile_12_filtered_output_c2(15);
   bh7_w57_5_c2 <= tile_12_filtered_output_c2(16);
   bh7_w58_4_c2 <= tile_12_filtered_output_c2(17);
   bh7_w59_3_c2 <= tile_12_filtered_output_c2(18);
   bh7_w60_4_c2 <= tile_12_filtered_output_c2(19);
   bh7_w61_4_c2 <= tile_12_filtered_output_c2(20);
   bh7_w62_3_c2 <= tile_12_filtered_output_c2(21);
   bh7_w63_4_c2 <= tile_12_filtered_output_c2(22);
   bh7_w64_4_c2 <= tile_12_filtered_output_c2(23);
   bh7_w65_2_c2 <= tile_12_filtered_output_c2(24);
   bh7_w66_3_c2 <= tile_12_filtered_output_c2(25);
   bh7_w67_3_c2 <= tile_12_filtered_output_c2(26);
   bh7_w68_2_c2 <= tile_12_filtered_output_c2(27);
   bh7_w69_3_c2 <= tile_12_filtered_output_c2(28);
   bh7_w70_3_c2 <= tile_12_filtered_output_c2(29);
   bh7_w71_2_c2 <= tile_12_filtered_output_c2(30);
   bh7_w72_3_c2 <= tile_12_filtered_output_c2(31);
   bh7_w73_3_c2 <= tile_12_filtered_output_c2(32);
   bh7_w74_2_c2 <= tile_12_filtered_output_c2(33);
   bh7_w75_1_c2 <= tile_12_filtered_output_c2(34);
   bh7_w76_1_c2 <= tile_12_filtered_output_c2(35);
   bh7_w77_0_c2 <= tile_12_filtered_output_c2(36);
   bh7_w78_0_c2 <= tile_12_filtered_output_c2(37);
   bh7_w79_0_c2 <= tile_12_filtered_output_c2(38);
   bh7_w80_0_c2 <= tile_12_filtered_output_c2(39);
   bh7_w81_0_c2 <= tile_12_filtered_output_c2(40);
   tile_13_X_c0 <= X(50 downto 34);
   tile_13_Y_c0 <= Y(47 downto 24);
   tile_13_mult: DSPBlock_17x24_Freq800_uid59
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => tile_13_X_c0,
                 Y => tile_13_Y_c0,
                 R => tile_13_output_c2);

   tile_13_filtered_output_c2 <= unsigned(tile_13_output_c2(40 downto 0));
   bh7_w58_5_c2 <= tile_13_filtered_output_c2(0);
   bh7_w59_4_c2 <= tile_13_filtered_output_c2(1);
   bh7_w60_5_c2 <= tile_13_filtered_output_c2(2);
   bh7_w61_5_c2 <= tile_13_filtered_output_c2(3);
   bh7_w62_4_c2 <= tile_13_filtered_output_c2(4);
   bh7_w63_5_c2 <= tile_13_filtered_output_c2(5);
   bh7_w64_5_c2 <= tile_13_filtered_output_c2(6);
   bh7_w65_3_c2 <= tile_13_filtered_output_c2(7);
   bh7_w66_4_c2 <= tile_13_filtered_output_c2(8);
   bh7_w67_4_c2 <= tile_13_filtered_output_c2(9);
   bh7_w68_3_c2 <= tile_13_filtered_output_c2(10);
   bh7_w69_4_c2 <= tile_13_filtered_output_c2(11);
   bh7_w70_4_c2 <= tile_13_filtered_output_c2(12);
   bh7_w71_3_c2 <= tile_13_filtered_output_c2(13);
   bh7_w72_4_c2 <= tile_13_filtered_output_c2(14);
   bh7_w73_4_c2 <= tile_13_filtered_output_c2(15);
   bh7_w74_3_c2 <= tile_13_filtered_output_c2(16);
   bh7_w75_2_c2 <= tile_13_filtered_output_c2(17);
   bh7_w76_2_c2 <= tile_13_filtered_output_c2(18);
   bh7_w77_1_c2 <= tile_13_filtered_output_c2(19);
   bh7_w78_1_c2 <= tile_13_filtered_output_c2(20);
   bh7_w79_1_c2 <= tile_13_filtered_output_c2(21);
   bh7_w80_1_c2 <= tile_13_filtered_output_c2(22);
   bh7_w81_1_c2 <= tile_13_filtered_output_c2(23);
   bh7_w82_0_c2 <= tile_13_filtered_output_c2(24);
   bh7_w83_0_c2 <= tile_13_filtered_output_c2(25);
   bh7_w84_0_c2 <= tile_13_filtered_output_c2(26);
   bh7_w85_0_c2 <= tile_13_filtered_output_c2(27);
   bh7_w86_0_c2 <= tile_13_filtered_output_c2(28);
   bh7_w87_0_c2 <= tile_13_filtered_output_c2(29);
   bh7_w88_0_c2 <= tile_13_filtered_output_c2(30);
   bh7_w89_0_c2 <= tile_13_filtered_output_c2(31);
   bh7_w90_0_c2 <= tile_13_filtered_output_c2(32);
   bh7_w91_0_c2 <= tile_13_filtered_output_c2(33);
   bh7_w92_0_c2 <= tile_13_filtered_output_c2(34);
   bh7_w93_0_c2 <= tile_13_filtered_output_c2(35);
   bh7_w94_0_c2 <= tile_13_filtered_output_c2(36);
   bh7_w95_0_c2 <= tile_13_filtered_output_c2(37);
   bh7_w96_0_c2 <= tile_13_filtered_output_c2(38);
   bh7_w97_0_c2 <= tile_13_filtered_output_c2(39);
   bh7_w98_0_c2 <= tile_13_filtered_output_c2(40);
   tile_14_X_c0 <= X(52 downto 51);
   tile_14_Y_c0 <= Y(47 downto 45);
   tile_14_mult: IntMultiplierLUT_2x3_Freq800_uid61
      port map ( clk  => clk,
                 X => tile_14_X_c0,
                 Y => tile_14_Y_c0,
                 R => tile_14_output_c0);

   tile_14_filtered_output_c0 <= unsigned(tile_14_output_c0(4 downto 0));
   bh7_w96_1_c0 <= tile_14_filtered_output_c0(0);
   bh7_w97_1_c0 <= tile_14_filtered_output_c0(1);
   bh7_w98_1_c0 <= tile_14_filtered_output_c0(2);
   bh7_w99_0_c0 <= tile_14_filtered_output_c0(3);
   bh7_w100_0_c0 <= tile_14_filtered_output_c0(4);
   tile_15_X_c0 <= X(52 downto 51);
   tile_15_Y_c0 <= Y(44 downto 42);
   tile_15_mult: IntMultiplierLUT_2x3_Freq800_uid66
      port map ( clk  => clk,
                 X => tile_15_X_c0,
                 Y => tile_15_Y_c0,
                 R => tile_15_output_c0);

   tile_15_filtered_output_c0 <= unsigned(tile_15_output_c0(4 downto 0));
   bh7_w93_1_c0 <= tile_15_filtered_output_c0(0);
   bh7_w94_1_c0 <= tile_15_filtered_output_c0(1);
   bh7_w95_1_c0 <= tile_15_filtered_output_c0(2);
   bh7_w96_2_c0 <= tile_15_filtered_output_c0(3);
   bh7_w97_2_c0 <= tile_15_filtered_output_c0(4);
   tile_16_X_c0 <= X(52 downto 51);
   tile_16_Y_c0 <= Y(41 downto 39);
   tile_16_mult: IntMultiplierLUT_2x3_Freq800_uid71
      port map ( clk  => clk,
                 X => tile_16_X_c0,
                 Y => tile_16_Y_c0,
                 R => tile_16_output_c0);

   tile_16_filtered_output_c0 <= unsigned(tile_16_output_c0(4 downto 0));
   bh7_w90_1_c0 <= tile_16_filtered_output_c0(0);
   bh7_w91_1_c0 <= tile_16_filtered_output_c0(1);
   bh7_w92_1_c0 <= tile_16_filtered_output_c0(2);
   bh7_w93_2_c0 <= tile_16_filtered_output_c0(3);
   bh7_w94_2_c0 <= tile_16_filtered_output_c0(4);
   tile_17_X_c0 <= X(52 downto 51);
   tile_17_Y_c0 <= Y(38 downto 36);
   tile_17_mult: IntMultiplierLUT_2x3_Freq800_uid76
      port map ( clk  => clk,
                 X => tile_17_X_c0,
                 Y => tile_17_Y_c0,
                 R => tile_17_output_c0);

   tile_17_filtered_output_c0 <= unsigned(tile_17_output_c0(4 downto 0));
   bh7_w87_1_c0 <= tile_17_filtered_output_c0(0);
   bh7_w88_1_c0 <= tile_17_filtered_output_c0(1);
   bh7_w89_1_c0 <= tile_17_filtered_output_c0(2);
   bh7_w90_2_c0 <= tile_17_filtered_output_c0(3);
   bh7_w91_2_c0 <= tile_17_filtered_output_c0(4);
   tile_18_X_c0 <= X(52 downto 51);
   tile_18_Y_c0 <= Y(35 downto 33);
   tile_18_mult: IntMultiplierLUT_2x3_Freq800_uid81
      port map ( clk  => clk,
                 X => tile_18_X_c0,
                 Y => tile_18_Y_c0,
                 R => tile_18_output_c0);

   tile_18_filtered_output_c0 <= unsigned(tile_18_output_c0(4 downto 0));
   bh7_w84_1_c0 <= tile_18_filtered_output_c0(0);
   bh7_w85_1_c0 <= tile_18_filtered_output_c0(1);
   bh7_w86_1_c0 <= tile_18_filtered_output_c0(2);
   bh7_w87_2_c0 <= tile_18_filtered_output_c0(3);
   bh7_w88_2_c0 <= tile_18_filtered_output_c0(4);
   tile_19_X_c0 <= X(52 downto 51);
   tile_19_Y_c0 <= Y(32 downto 30);
   tile_19_mult: IntMultiplierLUT_2x3_Freq800_uid86
      port map ( clk  => clk,
                 X => tile_19_X_c0,
                 Y => tile_19_Y_c0,
                 R => tile_19_output_c0);

   tile_19_filtered_output_c0 <= unsigned(tile_19_output_c0(4 downto 0));
   bh7_w81_2_c0 <= tile_19_filtered_output_c0(0);
   bh7_w82_1_c0 <= tile_19_filtered_output_c0(1);
   bh7_w83_1_c0 <= tile_19_filtered_output_c0(2);
   bh7_w84_2_c0 <= tile_19_filtered_output_c0(3);
   bh7_w85_2_c0 <= tile_19_filtered_output_c0(4);
   tile_20_X_c0 <= X(52 downto 51);
   tile_20_Y_c0 <= Y(29 downto 27);
   tile_20_mult: IntMultiplierLUT_2x3_Freq800_uid91
      port map ( clk  => clk,
                 X => tile_20_X_c0,
                 Y => tile_20_Y_c0,
                 R => tile_20_output_c0);

   tile_20_filtered_output_c0 <= unsigned(tile_20_output_c0(4 downto 0));
   bh7_w78_2_c0 <= tile_20_filtered_output_c0(0);
   bh7_w79_2_c0 <= tile_20_filtered_output_c0(1);
   bh7_w80_2_c0 <= tile_20_filtered_output_c0(2);
   bh7_w81_3_c0 <= tile_20_filtered_output_c0(3);
   bh7_w82_2_c0 <= tile_20_filtered_output_c0(4);
   tile_21_X_c0 <= X(52 downto 51);
   tile_21_Y_c0 <= Y(26 downto 24);
   tile_21_mult: IntMultiplierLUT_2x3_Freq800_uid96
      port map ( clk  => clk,
                 X => tile_21_X_c0,
                 Y => tile_21_Y_c0,
                 R => tile_21_output_c0);

   tile_21_filtered_output_c0 <= unsigned(tile_21_output_c0(4 downto 0));
   bh7_w75_3_c0 <= tile_21_filtered_output_c0(0);
   bh7_w76_3_c0 <= tile_21_filtered_output_c0(1);
   bh7_w77_2_c0 <= tile_21_filtered_output_c0(2);
   bh7_w78_3_c0 <= tile_21_filtered_output_c0(3);
   bh7_w79_3_c0 <= tile_21_filtered_output_c0(4);
   tile_22_X_c0 <= X(16 downto 16);
   tile_22_Y_c0 <= Y(52 downto 52);
   tile_22_mult: IntMultiplierLUT_1x1_Freq800_uid101
      port map ( clk  => clk,
                 X => tile_22_X_c0,
                 Y => tile_22_Y_c0,
                 R => tile_22_output_c0);

   tile_22_filtered_output_c0 <= unsigned(tile_22_output_c0(0 downto 0));
   bh7_w68_4_c0 <= tile_22_filtered_output_c0(0);
   tile_23_X_c0 <= X(15 downto 12);
   tile_23_Y_c0 <= Y(52 downto 52);
   tile_23_mult: IntMultiplierLUT_4x1_Freq800_uid103
      port map ( clk  => clk,
                 X => tile_23_X_c0,
                 Y => tile_23_Y_c0,
                 R => tile_23_output_c0);

   tile_23_filtered_output_c0 <= unsigned(tile_23_output_c0(3 downto 0));
   bh7_w64_6_c0 <= tile_23_filtered_output_c0(0);
   bh7_w65_4_c0 <= tile_23_filtered_output_c0(1);
   bh7_w66_5_c0 <= tile_23_filtered_output_c0(2);
   bh7_w67_5_c0 <= tile_23_filtered_output_c0(3);
   tile_24_X_c0 <= X(11 downto 8);
   tile_24_Y_c0 <= Y(52 downto 52);
   tile_24_mult: IntMultiplierLUT_4x1_Freq800_uid105
      port map ( clk  => clk,
                 X => tile_24_X_c0,
                 Y => tile_24_Y_c0,
                 R => tile_24_output_c0);

   tile_24_filtered_output_c0 <= unsigned(tile_24_output_c0(3 downto 0));
   bh7_w60_6_c0 <= tile_24_filtered_output_c0(0);
   bh7_w61_6_c0 <= tile_24_filtered_output_c0(1);
   bh7_w62_5_c0 <= tile_24_filtered_output_c0(2);
   bh7_w63_6_c0 <= tile_24_filtered_output_c0(3);
   tile_25_X_c0 <= X(7 downto 4);
   tile_25_Y_c0 <= Y(52 downto 52);
   tile_25_mult: IntMultiplierLUT_4x1_Freq800_uid107
      port map ( clk  => clk,
                 X => tile_25_X_c0,
                 Y => tile_25_Y_c0,
                 R => tile_25_output_c0);

   tile_25_filtered_output_c0 <= unsigned(tile_25_output_c0(3 downto 0));
   bh7_w56_5_c0 <= tile_25_filtered_output_c0(0);
   bh7_w57_6_c0 <= tile_25_filtered_output_c0(1);
   bh7_w58_6_c0 <= tile_25_filtered_output_c0(2);
   bh7_w59_5_c0 <= tile_25_filtered_output_c0(3);
   tile_26_X_c0 <= X(3 downto 0);
   tile_26_Y_c0 <= Y(52 downto 52);
   tile_26_mult: IntMultiplierLUT_4x1_Freq800_uid109
      port map ( clk  => clk,
                 X => tile_26_X_c0,
                 Y => tile_26_Y_c0,
                 R => tile_26_output_c0);

   tile_26_filtered_output_c0 <= unsigned(tile_26_output_c0(3 downto 0));
   bh7_w52_5_c0 <= tile_26_filtered_output_c0(0);
   bh7_w53_5_c0 <= tile_26_filtered_output_c0(1);
   bh7_w54_6_c0 <= tile_26_filtered_output_c0(2);
   bh7_w55_6_c0 <= tile_26_filtered_output_c0(3);
   tile_27_X_c0 <= X(16 downto 15);
   tile_27_Y_c0 <= Y(51 downto 50);
   tile_27_mult: IntMultiplierLUT_2x2_Freq800_uid111
      port map ( clk  => clk,
                 X => tile_27_X_c0,
                 Y => tile_27_Y_c0,
                 R => tile_27_output_c0);

   tile_27_filtered_output_c0 <= unsigned(tile_27_output_c0(3 downto 0));
   bh7_w65_5_c0 <= tile_27_filtered_output_c0(0);
   bh7_w66_6_c0 <= tile_27_filtered_output_c0(1);
   bh7_w67_6_c0 <= tile_27_filtered_output_c0(2);
   bh7_w68_5_c0 <= tile_27_filtered_output_c0(3);
   tile_28_X_c0 <= X(14 downto 12);
   tile_28_Y_c0 <= Y(51 downto 50);
   tile_28_mult: IntMultiplierLUT_3x2_Freq800_uid116
      port map ( clk  => clk,
                 X => tile_28_X_c0,
                 Y => tile_28_Y_c0,
                 R => tile_28_output_c0);

   tile_28_filtered_output_c0 <= unsigned(tile_28_output_c0(4 downto 0));
   bh7_w62_6_c0 <= tile_28_filtered_output_c0(0);
   bh7_w63_7_c0 <= tile_28_filtered_output_c0(1);
   bh7_w64_7_c0 <= tile_28_filtered_output_c0(2);
   bh7_w65_6_c0 <= tile_28_filtered_output_c0(3);
   bh7_w66_7_c0 <= tile_28_filtered_output_c0(4);
   tile_29_X_c0 <= X(11 downto 9);
   tile_29_Y_c0 <= Y(51 downto 50);
   tile_29_mult: IntMultiplierLUT_3x2_Freq800_uid121
      port map ( clk  => clk,
                 X => tile_29_X_c0,
                 Y => tile_29_Y_c0,
                 R => tile_29_output_c0);

   tile_29_filtered_output_c0 <= unsigned(tile_29_output_c0(4 downto 0));
   bh7_w59_6_c0 <= tile_29_filtered_output_c0(0);
   bh7_w60_7_c0 <= tile_29_filtered_output_c0(1);
   bh7_w61_7_c0 <= tile_29_filtered_output_c0(2);
   bh7_w62_7_c0 <= tile_29_filtered_output_c0(3);
   bh7_w63_8_c0 <= tile_29_filtered_output_c0(4);
   tile_30_X_c0 <= X(8 downto 6);
   tile_30_Y_c0 <= Y(51 downto 50);
   tile_30_mult: IntMultiplierLUT_3x2_Freq800_uid126
      port map ( clk  => clk,
                 X => tile_30_X_c0,
                 Y => tile_30_Y_c0,
                 R => tile_30_output_c0);

   tile_30_filtered_output_c0 <= unsigned(tile_30_output_c0(4 downto 0));
   bh7_w56_6_c0 <= tile_30_filtered_output_c0(0);
   bh7_w57_7_c0 <= tile_30_filtered_output_c0(1);
   bh7_w58_7_c0 <= tile_30_filtered_output_c0(2);
   bh7_w59_7_c0 <= tile_30_filtered_output_c0(3);
   bh7_w60_8_c0 <= tile_30_filtered_output_c0(4);
   tile_31_X_c0 <= X(5 downto 3);
   tile_31_Y_c0 <= Y(51 downto 50);
   tile_31_mult: IntMultiplierLUT_3x2_Freq800_uid131
      port map ( clk  => clk,
                 X => tile_31_X_c0,
                 Y => tile_31_Y_c0,
                 R => tile_31_output_c0);

   tile_31_filtered_output_c0 <= unsigned(tile_31_output_c0(4 downto 0));
   bh7_w53_6_c0 <= tile_31_filtered_output_c0(0);
   bh7_w54_7_c0 <= tile_31_filtered_output_c0(1);
   bh7_w55_7_c0 <= tile_31_filtered_output_c0(2);
   bh7_w56_7_c0 <= tile_31_filtered_output_c0(3);
   bh7_w57_8_c0 <= tile_31_filtered_output_c0(4);
   tile_32_X_c0 <= X(2 downto 0);
   tile_32_Y_c0 <= Y(51 downto 50);
   tile_32_mult: IntMultiplierLUT_3x2_Freq800_uid136
      port map ( clk  => clk,
                 X => tile_32_X_c0,
                 Y => tile_32_Y_c0,
                 R => tile_32_output_c0);

   tile_32_filtered_output_c0 <= unsigned(tile_32_output_c0(4 downto 0));
   bh7_w50_4_c0 <= tile_32_filtered_output_c0(0);
   bh7_w51_5_c0 <= tile_32_filtered_output_c0(1);
   bh7_w52_6_c0 <= tile_32_filtered_output_c0(2);
   bh7_w53_7_c0 <= tile_32_filtered_output_c0(3);
   bh7_w54_8_c0 <= tile_32_filtered_output_c0(4);
   tile_33_X_c0 <= X(16 downto 15);
   tile_33_Y_c0 <= Y(49 downto 48);
   tile_33_mult: IntMultiplierLUT_2x2_Freq800_uid141
      port map ( clk  => clk,
                 X => tile_33_X_c0,
                 Y => tile_33_Y_c0,
                 R => tile_33_output_c0);

   tile_33_filtered_output_c0 <= unsigned(tile_33_output_c0(3 downto 0));
   bh7_w63_9_c0 <= tile_33_filtered_output_c0(0);
   bh7_w64_8_c0 <= tile_33_filtered_output_c0(1);
   bh7_w65_7_c0 <= tile_33_filtered_output_c0(2);
   bh7_w66_8_c0 <= tile_33_filtered_output_c0(3);
   tile_34_X_c0 <= X(14 downto 12);
   tile_34_Y_c0 <= Y(49 downto 48);
   tile_34_mult: IntMultiplierLUT_3x2_Freq800_uid146
      port map ( clk  => clk,
                 X => tile_34_X_c0,
                 Y => tile_34_Y_c0,
                 R => tile_34_output_c0);

   tile_34_filtered_output_c0 <= unsigned(tile_34_output_c0(4 downto 0));
   bh7_w60_9_c0 <= tile_34_filtered_output_c0(0);
   bh7_w61_8_c0 <= tile_34_filtered_output_c0(1);
   bh7_w62_8_c0 <= tile_34_filtered_output_c0(2);
   bh7_w63_10_c0 <= tile_34_filtered_output_c0(3);
   bh7_w64_9_c0 <= tile_34_filtered_output_c0(4);
   tile_35_X_c0 <= X(11 downto 9);
   tile_35_Y_c0 <= Y(49 downto 48);
   tile_35_mult: IntMultiplierLUT_3x2_Freq800_uid151
      port map ( clk  => clk,
                 X => tile_35_X_c0,
                 Y => tile_35_Y_c0,
                 R => tile_35_output_c0);

   tile_35_filtered_output_c0 <= unsigned(tile_35_output_c0(4 downto 0));
   bh7_w57_9_c0 <= tile_35_filtered_output_c0(0);
   bh7_w58_8_c0 <= tile_35_filtered_output_c0(1);
   bh7_w59_8_c0 <= tile_35_filtered_output_c0(2);
   bh7_w60_10_c0 <= tile_35_filtered_output_c0(3);
   bh7_w61_9_c0 <= tile_35_filtered_output_c0(4);
   tile_36_X_c0 <= X(8 downto 6);
   tile_36_Y_c0 <= Y(49 downto 48);
   tile_36_mult: IntMultiplierLUT_3x2_Freq800_uid156
      port map ( clk  => clk,
                 X => tile_36_X_c0,
                 Y => tile_36_Y_c0,
                 R => tile_36_output_c0);

   tile_36_filtered_output_c0 <= unsigned(tile_36_output_c0(4 downto 0));
   bh7_w54_9_c0 <= tile_36_filtered_output_c0(0);
   bh7_w55_8_c0 <= tile_36_filtered_output_c0(1);
   bh7_w56_8_c0 <= tile_36_filtered_output_c0(2);
   bh7_w57_10_c0 <= tile_36_filtered_output_c0(3);
   bh7_w58_9_c0 <= tile_36_filtered_output_c0(4);
   tile_37_X_c0 <= X(5 downto 3);
   tile_37_Y_c0 <= Y(49 downto 48);
   tile_37_mult: IntMultiplierLUT_3x2_Freq800_uid161
      port map ( clk  => clk,
                 X => tile_37_X_c0,
                 Y => tile_37_Y_c0,
                 R => tile_37_output_c0);

   tile_37_filtered_output_c0 <= unsigned(tile_37_output_c0(4 downto 0));
   bh7_w51_6_c0 <= tile_37_filtered_output_c0(0);
   bh7_w52_7_c0 <= tile_37_filtered_output_c0(1);
   bh7_w53_8_c0 <= tile_37_filtered_output_c0(2);
   bh7_w54_10_c0 <= tile_37_filtered_output_c0(3);
   bh7_w55_9_c0 <= tile_37_filtered_output_c0(4);
   tile_38_X_c0 <= X(2 downto 0);
   tile_38_Y_c0 <= Y(49 downto 48);
   tile_38_mult: IntMultiplierLUT_3x2_Freq800_uid166
      port map ( clk  => clk,
                 X => tile_38_X_c0,
                 Y => tile_38_Y_c0,
                 R => tile_38_output_c0);

   tile_38_filtered_output_c0 <= unsigned(tile_38_output_c0(4 downto 0));
   bh7_w48_4_c0 <= tile_38_filtered_output_c0(0);
   bh7_w49_4_c0 <= tile_38_filtered_output_c0(1);
   bh7_w50_5_c0 <= tile_38_filtered_output_c0(2);
   bh7_w51_7_c0 <= tile_38_filtered_output_c0(3);
   bh7_w52_8_c0 <= tile_38_filtered_output_c0(4);
   tile_39_X_c0 <= X(33 downto 33);
   tile_39_Y_c0 <= Y(52 downto 52);
   tile_39_mult: IntMultiplierLUT_1x1_Freq800_uid171
      port map ( clk  => clk,
                 X => tile_39_X_c0,
                 Y => tile_39_Y_c0,
                 R => tile_39_output_c0);

   tile_39_filtered_output_c0 <= unsigned(tile_39_output_c0(0 downto 0));
   bh7_w85_3_c0 <= tile_39_filtered_output_c0(0);
   tile_40_X_c0 <= X(32 downto 29);
   tile_40_Y_c0 <= Y(52 downto 52);
   tile_40_mult: IntMultiplierLUT_4x1_Freq800_uid173
      port map ( clk  => clk,
                 X => tile_40_X_c0,
                 Y => tile_40_Y_c0,
                 R => tile_40_output_c0);

   tile_40_filtered_output_c0 <= unsigned(tile_40_output_c0(3 downto 0));
   bh7_w81_4_c0 <= tile_40_filtered_output_c0(0);
   bh7_w82_3_c0 <= tile_40_filtered_output_c0(1);
   bh7_w83_2_c0 <= tile_40_filtered_output_c0(2);
   bh7_w84_3_c0 <= tile_40_filtered_output_c0(3);
   tile_41_X_c0 <= X(28 downto 25);
   tile_41_Y_c0 <= Y(52 downto 52);
   tile_41_mult: IntMultiplierLUT_4x1_Freq800_uid175
      port map ( clk  => clk,
                 X => tile_41_X_c0,
                 Y => tile_41_Y_c0,
                 R => tile_41_output_c0);

   tile_41_filtered_output_c0 <= unsigned(tile_41_output_c0(3 downto 0));
   bh7_w77_3_c0 <= tile_41_filtered_output_c0(0);
   bh7_w78_4_c0 <= tile_41_filtered_output_c0(1);
   bh7_w79_4_c0 <= tile_41_filtered_output_c0(2);
   bh7_w80_3_c0 <= tile_41_filtered_output_c0(3);
   tile_42_X_c0 <= X(24 downto 21);
   tile_42_Y_c0 <= Y(52 downto 52);
   tile_42_mult: IntMultiplierLUT_4x1_Freq800_uid177
      port map ( clk  => clk,
                 X => tile_42_X_c0,
                 Y => tile_42_Y_c0,
                 R => tile_42_output_c0);

   tile_42_filtered_output_c0 <= unsigned(tile_42_output_c0(3 downto 0));
   bh7_w73_5_c0 <= tile_42_filtered_output_c0(0);
   bh7_w74_4_c0 <= tile_42_filtered_output_c0(1);
   bh7_w75_4_c0 <= tile_42_filtered_output_c0(2);
   bh7_w76_4_c0 <= tile_42_filtered_output_c0(3);
   tile_43_X_c0 <= X(20 downto 17);
   tile_43_Y_c0 <= Y(52 downto 52);
   tile_43_mult: IntMultiplierLUT_4x1_Freq800_uid179
      port map ( clk  => clk,
                 X => tile_43_X_c0,
                 Y => tile_43_Y_c0,
                 R => tile_43_output_c0);

   tile_43_filtered_output_c0 <= unsigned(tile_43_output_c0(3 downto 0));
   bh7_w69_5_c0 <= tile_43_filtered_output_c0(0);
   bh7_w70_5_c0 <= tile_43_filtered_output_c0(1);
   bh7_w71_4_c0 <= tile_43_filtered_output_c0(2);
   bh7_w72_5_c0 <= tile_43_filtered_output_c0(3);
   tile_44_X_c0 <= X(33 downto 32);
   tile_44_Y_c0 <= Y(51 downto 50);
   tile_44_mult: IntMultiplierLUT_2x2_Freq800_uid181
      port map ( clk  => clk,
                 X => tile_44_X_c0,
                 Y => tile_44_Y_c0,
                 R => tile_44_output_c0);

   tile_44_filtered_output_c0 <= unsigned(tile_44_output_c0(3 downto 0));
   bh7_w82_4_c0 <= tile_44_filtered_output_c0(0);
   bh7_w83_3_c0 <= tile_44_filtered_output_c0(1);
   bh7_w84_4_c0 <= tile_44_filtered_output_c0(2);
   bh7_w85_4_c0 <= tile_44_filtered_output_c0(3);
   tile_45_X_c0 <= X(31 downto 29);
   tile_45_Y_c0 <= Y(51 downto 50);
   tile_45_mult: IntMultiplierLUT_3x2_Freq800_uid186
      port map ( clk  => clk,
                 X => tile_45_X_c0,
                 Y => tile_45_Y_c0,
                 R => tile_45_output_c0);

   tile_45_filtered_output_c0 <= unsigned(tile_45_output_c0(4 downto 0));
   bh7_w79_5_c0 <= tile_45_filtered_output_c0(0);
   bh7_w80_4_c0 <= tile_45_filtered_output_c0(1);
   bh7_w81_5_c0 <= tile_45_filtered_output_c0(2);
   bh7_w82_5_c0 <= tile_45_filtered_output_c0(3);
   bh7_w83_4_c0 <= tile_45_filtered_output_c0(4);
   tile_46_X_c0 <= X(28 downto 26);
   tile_46_Y_c0 <= Y(51 downto 50);
   tile_46_mult: IntMultiplierLUT_3x2_Freq800_uid191
      port map ( clk  => clk,
                 X => tile_46_X_c0,
                 Y => tile_46_Y_c0,
                 R => tile_46_output_c0);

   tile_46_filtered_output_c0 <= unsigned(tile_46_output_c0(4 downto 0));
   bh7_w76_5_c0 <= tile_46_filtered_output_c0(0);
   bh7_w77_4_c0 <= tile_46_filtered_output_c0(1);
   bh7_w78_5_c0 <= tile_46_filtered_output_c0(2);
   bh7_w79_6_c0 <= tile_46_filtered_output_c0(3);
   bh7_w80_5_c0 <= tile_46_filtered_output_c0(4);
   tile_47_X_c0 <= X(25 downto 23);
   tile_47_Y_c0 <= Y(51 downto 50);
   tile_47_mult: IntMultiplierLUT_3x2_Freq800_uid196
      port map ( clk  => clk,
                 X => tile_47_X_c0,
                 Y => tile_47_Y_c0,
                 R => tile_47_output_c0);

   tile_47_filtered_output_c0 <= unsigned(tile_47_output_c0(4 downto 0));
   bh7_w73_6_c0 <= tile_47_filtered_output_c0(0);
   bh7_w74_5_c0 <= tile_47_filtered_output_c0(1);
   bh7_w75_5_c0 <= tile_47_filtered_output_c0(2);
   bh7_w76_6_c0 <= tile_47_filtered_output_c0(3);
   bh7_w77_5_c0 <= tile_47_filtered_output_c0(4);
   tile_48_X_c0 <= X(22 downto 20);
   tile_48_Y_c0 <= Y(51 downto 50);
   tile_48_mult: IntMultiplierLUT_3x2_Freq800_uid201
      port map ( clk  => clk,
                 X => tile_48_X_c0,
                 Y => tile_48_Y_c0,
                 R => tile_48_output_c0);

   tile_48_filtered_output_c0 <= unsigned(tile_48_output_c0(4 downto 0));
   bh7_w70_6_c0 <= tile_48_filtered_output_c0(0);
   bh7_w71_5_c0 <= tile_48_filtered_output_c0(1);
   bh7_w72_6_c0 <= tile_48_filtered_output_c0(2);
   bh7_w73_7_c0 <= tile_48_filtered_output_c0(3);
   bh7_w74_6_c0 <= tile_48_filtered_output_c0(4);
   tile_49_X_c0 <= X(19 downto 17);
   tile_49_Y_c0 <= Y(51 downto 50);
   tile_49_mult: IntMultiplierLUT_3x2_Freq800_uid206
      port map ( clk  => clk,
                 X => tile_49_X_c0,
                 Y => tile_49_Y_c0,
                 R => tile_49_output_c0);

   tile_49_filtered_output_c0 <= unsigned(tile_49_output_c0(4 downto 0));
   bh7_w67_7_c0 <= tile_49_filtered_output_c0(0);
   bh7_w68_6_c0 <= tile_49_filtered_output_c0(1);
   bh7_w69_6_c0 <= tile_49_filtered_output_c0(2);
   bh7_w70_7_c0 <= tile_49_filtered_output_c0(3);
   bh7_w71_6_c0 <= tile_49_filtered_output_c0(4);
   tile_50_X_c0 <= X(33 downto 32);
   tile_50_Y_c0 <= Y(49 downto 48);
   tile_50_mult: IntMultiplierLUT_2x2_Freq800_uid211
      port map ( clk  => clk,
                 X => tile_50_X_c0,
                 Y => tile_50_Y_c0,
                 R => tile_50_output_c0);

   tile_50_filtered_output_c0 <= unsigned(tile_50_output_c0(3 downto 0));
   bh7_w80_6_c0 <= tile_50_filtered_output_c0(0);
   bh7_w81_6_c0 <= tile_50_filtered_output_c0(1);
   bh7_w82_6_c0 <= tile_50_filtered_output_c0(2);
   bh7_w83_5_c0 <= tile_50_filtered_output_c0(3);
   tile_51_X_c0 <= X(31 downto 29);
   tile_51_Y_c0 <= Y(49 downto 48);
   tile_51_mult: IntMultiplierLUT_3x2_Freq800_uid216
      port map ( clk  => clk,
                 X => tile_51_X_c0,
                 Y => tile_51_Y_c0,
                 R => tile_51_output_c0);

   tile_51_filtered_output_c0 <= unsigned(tile_51_output_c0(4 downto 0));
   bh7_w77_6_c0 <= tile_51_filtered_output_c0(0);
   bh7_w78_6_c0 <= tile_51_filtered_output_c0(1);
   bh7_w79_7_c0 <= tile_51_filtered_output_c0(2);
   bh7_w80_7_c0 <= tile_51_filtered_output_c0(3);
   bh7_w81_7_c0 <= tile_51_filtered_output_c0(4);
   tile_52_X_c0 <= X(28 downto 26);
   tile_52_Y_c0 <= Y(49 downto 48);
   tile_52_mult: IntMultiplierLUT_3x2_Freq800_uid221
      port map ( clk  => clk,
                 X => tile_52_X_c0,
                 Y => tile_52_Y_c0,
                 R => tile_52_output_c0);

   tile_52_filtered_output_c0 <= unsigned(tile_52_output_c0(4 downto 0));
   bh7_w74_7_c0 <= tile_52_filtered_output_c0(0);
   bh7_w75_6_c0 <= tile_52_filtered_output_c0(1);
   bh7_w76_7_c0 <= tile_52_filtered_output_c0(2);
   bh7_w77_7_c0 <= tile_52_filtered_output_c0(3);
   bh7_w78_7_c0 <= tile_52_filtered_output_c0(4);
   tile_53_X_c0 <= X(25 downto 23);
   tile_53_Y_c0 <= Y(49 downto 48);
   tile_53_mult: IntMultiplierLUT_3x2_Freq800_uid226
      port map ( clk  => clk,
                 X => tile_53_X_c0,
                 Y => tile_53_Y_c0,
                 R => tile_53_output_c0);

   tile_53_filtered_output_c0 <= unsigned(tile_53_output_c0(4 downto 0));
   bh7_w71_7_c0 <= tile_53_filtered_output_c0(0);
   bh7_w72_7_c0 <= tile_53_filtered_output_c0(1);
   bh7_w73_8_c0 <= tile_53_filtered_output_c0(2);
   bh7_w74_8_c0 <= tile_53_filtered_output_c0(3);
   bh7_w75_7_c0 <= tile_53_filtered_output_c0(4);
   tile_54_X_c0 <= X(22 downto 20);
   tile_54_Y_c0 <= Y(49 downto 48);
   tile_54_mult: IntMultiplierLUT_3x2_Freq800_uid231
      port map ( clk  => clk,
                 X => tile_54_X_c0,
                 Y => tile_54_Y_c0,
                 R => tile_54_output_c0);

   tile_54_filtered_output_c0 <= unsigned(tile_54_output_c0(4 downto 0));
   bh7_w68_7_c0 <= tile_54_filtered_output_c0(0);
   bh7_w69_7_c0 <= tile_54_filtered_output_c0(1);
   bh7_w70_8_c0 <= tile_54_filtered_output_c0(2);
   bh7_w71_8_c0 <= tile_54_filtered_output_c0(3);
   bh7_w72_8_c0 <= tile_54_filtered_output_c0(4);
   tile_55_X_c0 <= X(19 downto 17);
   tile_55_Y_c0 <= Y(49 downto 48);
   tile_55_mult: IntMultiplierLUT_3x2_Freq800_uid236
      port map ( clk  => clk,
                 X => tile_55_X_c0,
                 Y => tile_55_Y_c0,
                 R => tile_55_output_c0);

   tile_55_filtered_output_c0 <= unsigned(tile_55_output_c0(4 downto 0));
   bh7_w65_8_c0 <= tile_55_filtered_output_c0(0);
   bh7_w66_9_c0 <= tile_55_filtered_output_c0(1);
   bh7_w67_8_c0 <= tile_55_filtered_output_c0(2);
   bh7_w68_8_c0 <= tile_55_filtered_output_c0(3);
   bh7_w69_8_c0 <= tile_55_filtered_output_c0(4);
   tile_56_X_c0 <= X(50 downto 50);
   tile_56_Y_c0 <= Y(52 downto 52);
   tile_56_mult: IntMultiplierLUT_1x1_Freq800_uid241
      port map ( clk  => clk,
                 X => tile_56_X_c0,
                 Y => tile_56_Y_c0,
                 R => tile_56_output_c0);

   tile_56_filtered_output_c0 <= unsigned(tile_56_output_c0(0 downto 0));
   bh7_w102_0_c0 <= tile_56_filtered_output_c0(0);
   tile_57_X_c0 <= X(49 downto 46);
   tile_57_Y_c0 <= Y(52 downto 52);
   tile_57_mult: IntMultiplierLUT_4x1_Freq800_uid243
      port map ( clk  => clk,
                 X => tile_57_X_c0,
                 Y => tile_57_Y_c0,
                 R => tile_57_output_c0);

   tile_57_filtered_output_c0 <= unsigned(tile_57_output_c0(3 downto 0));
   bh7_w98_2_c0 <= tile_57_filtered_output_c0(0);
   bh7_w99_1_c0 <= tile_57_filtered_output_c0(1);
   bh7_w100_1_c0 <= tile_57_filtered_output_c0(2);
   bh7_w101_0_c0 <= tile_57_filtered_output_c0(3);
   tile_58_X_c0 <= X(45 downto 42);
   tile_58_Y_c0 <= Y(52 downto 52);
   tile_58_mult: IntMultiplierLUT_4x1_Freq800_uid245
      port map ( clk  => clk,
                 X => tile_58_X_c0,
                 Y => tile_58_Y_c0,
                 R => tile_58_output_c0);

   tile_58_filtered_output_c0 <= unsigned(tile_58_output_c0(3 downto 0));
   bh7_w94_3_c0 <= tile_58_filtered_output_c0(0);
   bh7_w95_2_c0 <= tile_58_filtered_output_c0(1);
   bh7_w96_3_c0 <= tile_58_filtered_output_c0(2);
   bh7_w97_3_c0 <= tile_58_filtered_output_c0(3);
   tile_59_X_c0 <= X(41 downto 38);
   tile_59_Y_c0 <= Y(52 downto 52);
   tile_59_mult: IntMultiplierLUT_4x1_Freq800_uid247
      port map ( clk  => clk,
                 X => tile_59_X_c0,
                 Y => tile_59_Y_c0,
                 R => tile_59_output_c0);

   tile_59_filtered_output_c0 <= unsigned(tile_59_output_c0(3 downto 0));
   bh7_w90_3_c0 <= tile_59_filtered_output_c0(0);
   bh7_w91_3_c0 <= tile_59_filtered_output_c0(1);
   bh7_w92_2_c0 <= tile_59_filtered_output_c0(2);
   bh7_w93_3_c0 <= tile_59_filtered_output_c0(3);
   tile_60_X_c0 <= X(37 downto 34);
   tile_60_Y_c0 <= Y(52 downto 52);
   tile_60_mult: IntMultiplierLUT_4x1_Freq800_uid249
      port map ( clk  => clk,
                 X => tile_60_X_c0,
                 Y => tile_60_Y_c0,
                 R => tile_60_output_c0);

   tile_60_filtered_output_c0 <= unsigned(tile_60_output_c0(3 downto 0));
   bh7_w86_2_c0 <= tile_60_filtered_output_c0(0);
   bh7_w87_3_c0 <= tile_60_filtered_output_c0(1);
   bh7_w88_3_c0 <= tile_60_filtered_output_c0(2);
   bh7_w89_2_c0 <= tile_60_filtered_output_c0(3);
   tile_61_X_c0 <= X(50 downto 49);
   tile_61_Y_c0 <= Y(51 downto 50);
   tile_61_mult: IntMultiplierLUT_2x2_Freq800_uid251
      port map ( clk  => clk,
                 X => tile_61_X_c0,
                 Y => tile_61_Y_c0,
                 R => tile_61_output_c0);

   tile_61_filtered_output_c0 <= unsigned(tile_61_output_c0(3 downto 0));
   bh7_w99_2_c0 <= tile_61_filtered_output_c0(0);
   bh7_w100_2_c0 <= tile_61_filtered_output_c0(1);
   bh7_w101_1_c0 <= tile_61_filtered_output_c0(2);
   bh7_w102_1_c0 <= tile_61_filtered_output_c0(3);
   tile_62_X_c0 <= X(48 downto 46);
   tile_62_Y_c0 <= Y(51 downto 50);
   tile_62_mult: IntMultiplierLUT_3x2_Freq800_uid256
      port map ( clk  => clk,
                 X => tile_62_X_c0,
                 Y => tile_62_Y_c0,
                 R => tile_62_output_c0);

   tile_62_filtered_output_c0 <= unsigned(tile_62_output_c0(4 downto 0));
   bh7_w96_4_c0 <= tile_62_filtered_output_c0(0);
   bh7_w97_4_c0 <= tile_62_filtered_output_c0(1);
   bh7_w98_3_c0 <= tile_62_filtered_output_c0(2);
   bh7_w99_3_c0 <= tile_62_filtered_output_c0(3);
   bh7_w100_3_c0 <= tile_62_filtered_output_c0(4);
   tile_63_X_c0 <= X(45 downto 43);
   tile_63_Y_c0 <= Y(51 downto 50);
   tile_63_mult: IntMultiplierLUT_3x2_Freq800_uid261
      port map ( clk  => clk,
                 X => tile_63_X_c0,
                 Y => tile_63_Y_c0,
                 R => tile_63_output_c0);

   tile_63_filtered_output_c0 <= unsigned(tile_63_output_c0(4 downto 0));
   bh7_w93_4_c0 <= tile_63_filtered_output_c0(0);
   bh7_w94_4_c0 <= tile_63_filtered_output_c0(1);
   bh7_w95_3_c0 <= tile_63_filtered_output_c0(2);
   bh7_w96_5_c0 <= tile_63_filtered_output_c0(3);
   bh7_w97_5_c0 <= tile_63_filtered_output_c0(4);
   tile_64_X_c0 <= X(42 downto 40);
   tile_64_Y_c0 <= Y(51 downto 50);
   tile_64_mult: IntMultiplierLUT_3x2_Freq800_uid266
      port map ( clk  => clk,
                 X => tile_64_X_c0,
                 Y => tile_64_Y_c0,
                 R => tile_64_output_c0);

   tile_64_filtered_output_c0 <= unsigned(tile_64_output_c0(4 downto 0));
   bh7_w90_4_c0 <= tile_64_filtered_output_c0(0);
   bh7_w91_4_c0 <= tile_64_filtered_output_c0(1);
   bh7_w92_3_c0 <= tile_64_filtered_output_c0(2);
   bh7_w93_5_c0 <= tile_64_filtered_output_c0(3);
   bh7_w94_5_c0 <= tile_64_filtered_output_c0(4);
   tile_65_X_c0 <= X(39 downto 37);
   tile_65_Y_c0 <= Y(51 downto 50);
   tile_65_mult: IntMultiplierLUT_3x2_Freq800_uid271
      port map ( clk  => clk,
                 X => tile_65_X_c0,
                 Y => tile_65_Y_c0,
                 R => tile_65_output_c0);

   tile_65_filtered_output_c0 <= unsigned(tile_65_output_c0(4 downto 0));
   bh7_w87_4_c0 <= tile_65_filtered_output_c0(0);
   bh7_w88_4_c0 <= tile_65_filtered_output_c0(1);
   bh7_w89_3_c0 <= tile_65_filtered_output_c0(2);
   bh7_w90_5_c0 <= tile_65_filtered_output_c0(3);
   bh7_w91_5_c0 <= tile_65_filtered_output_c0(4);
   tile_66_X_c0 <= X(36 downto 34);
   tile_66_Y_c0 <= Y(51 downto 50);
   tile_66_mult: IntMultiplierLUT_3x2_Freq800_uid276
      port map ( clk  => clk,
                 X => tile_66_X_c0,
                 Y => tile_66_Y_c0,
                 R => tile_66_output_c0);

   tile_66_filtered_output_c0 <= unsigned(tile_66_output_c0(4 downto 0));
   bh7_w84_5_c0 <= tile_66_filtered_output_c0(0);
   bh7_w85_5_c0 <= tile_66_filtered_output_c0(1);
   bh7_w86_3_c0 <= tile_66_filtered_output_c0(2);
   bh7_w87_5_c0 <= tile_66_filtered_output_c0(3);
   bh7_w88_5_c0 <= tile_66_filtered_output_c0(4);
   tile_67_X_c0 <= X(50 downto 49);
   tile_67_Y_c0 <= Y(49 downto 48);
   tile_67_mult: IntMultiplierLUT_2x2_Freq800_uid281
      port map ( clk  => clk,
                 X => tile_67_X_c0,
                 Y => tile_67_Y_c0,
                 R => tile_67_output_c0);

   tile_67_filtered_output_c0 <= unsigned(tile_67_output_c0(3 downto 0));
   bh7_w97_6_c0 <= tile_67_filtered_output_c0(0);
   bh7_w98_4_c0 <= tile_67_filtered_output_c0(1);
   bh7_w99_4_c0 <= tile_67_filtered_output_c0(2);
   bh7_w100_4_c0 <= tile_67_filtered_output_c0(3);
   tile_68_X_c0 <= X(48 downto 46);
   tile_68_Y_c0 <= Y(49 downto 48);
   tile_68_mult: IntMultiplierLUT_3x2_Freq800_uid286
      port map ( clk  => clk,
                 X => tile_68_X_c0,
                 Y => tile_68_Y_c0,
                 R => tile_68_output_c0);

   tile_68_filtered_output_c0 <= unsigned(tile_68_output_c0(4 downto 0));
   bh7_w94_6_c0 <= tile_68_filtered_output_c0(0);
   bh7_w95_4_c0 <= tile_68_filtered_output_c0(1);
   bh7_w96_6_c0 <= tile_68_filtered_output_c0(2);
   bh7_w97_7_c0 <= tile_68_filtered_output_c0(3);
   bh7_w98_5_c0 <= tile_68_filtered_output_c0(4);
   tile_69_X_c0 <= X(45 downto 43);
   tile_69_Y_c0 <= Y(49 downto 48);
   tile_69_mult: IntMultiplierLUT_3x2_Freq800_uid291
      port map ( clk  => clk,
                 X => tile_69_X_c0,
                 Y => tile_69_Y_c0,
                 R => tile_69_output_c0);

   tile_69_filtered_output_c0 <= unsigned(tile_69_output_c0(4 downto 0));
   bh7_w91_6_c0 <= tile_69_filtered_output_c0(0);
   bh7_w92_4_c0 <= tile_69_filtered_output_c0(1);
   bh7_w93_6_c0 <= tile_69_filtered_output_c0(2);
   bh7_w94_7_c0 <= tile_69_filtered_output_c0(3);
   bh7_w95_5_c0 <= tile_69_filtered_output_c0(4);
   tile_70_X_c0 <= X(42 downto 40);
   tile_70_Y_c0 <= Y(49 downto 48);
   tile_70_mult: IntMultiplierLUT_3x2_Freq800_uid296
      port map ( clk  => clk,
                 X => tile_70_X_c0,
                 Y => tile_70_Y_c0,
                 R => tile_70_output_c0);

   tile_70_filtered_output_c0 <= unsigned(tile_70_output_c0(4 downto 0));
   bh7_w88_6_c0 <= tile_70_filtered_output_c0(0);
   bh7_w89_4_c0 <= tile_70_filtered_output_c0(1);
   bh7_w90_6_c0 <= tile_70_filtered_output_c0(2);
   bh7_w91_7_c0 <= tile_70_filtered_output_c0(3);
   bh7_w92_5_c0 <= tile_70_filtered_output_c0(4);
   tile_71_X_c0 <= X(39 downto 37);
   tile_71_Y_c0 <= Y(49 downto 48);
   tile_71_mult: IntMultiplierLUT_3x2_Freq800_uid301
      port map ( clk  => clk,
                 X => tile_71_X_c0,
                 Y => tile_71_Y_c0,
                 R => tile_71_output_c0);

   tile_71_filtered_output_c0 <= unsigned(tile_71_output_c0(4 downto 0));
   bh7_w85_6_c0 <= tile_71_filtered_output_c0(0);
   bh7_w86_4_c0 <= tile_71_filtered_output_c0(1);
   bh7_w87_6_c0 <= tile_71_filtered_output_c0(2);
   bh7_w88_7_c0 <= tile_71_filtered_output_c0(3);
   bh7_w89_5_c0 <= tile_71_filtered_output_c0(4);
   tile_72_X_c0 <= X(36 downto 34);
   tile_72_Y_c0 <= Y(49 downto 48);
   tile_72_mult: IntMultiplierLUT_3x2_Freq800_uid306
      port map ( clk  => clk,
                 X => tile_72_X_c0,
                 Y => tile_72_Y_c0,
                 R => tile_72_output_c0);

   tile_72_filtered_output_c0 <= unsigned(tile_72_output_c0(4 downto 0));
   bh7_w82_7_c0 <= tile_72_filtered_output_c0(0);
   bh7_w83_6_c0 <= tile_72_filtered_output_c0(1);
   bh7_w84_6_c0 <= tile_72_filtered_output_c0(2);
   bh7_w85_7_c0 <= tile_72_filtered_output_c0(3);
   bh7_w86_5_c0 <= tile_72_filtered_output_c0(4);
   tile_73_X_c0 <= X(52 downto 51);
   tile_73_Y_c0 <= Y(52 downto 51);
   tile_73_mult: IntMultiplierLUT_2x2_Freq800_uid311
      port map ( clk  => clk,
                 X => tile_73_X_c0,
                 Y => tile_73_Y_c0,
                 R => tile_73_output_c0);

   tile_73_filtered_output_c0 <= unsigned(tile_73_output_c0(3 downto 0));
   bh7_w102_2_c0 <= tile_73_filtered_output_c0(0);
   bh7_w103_0_c0 <= tile_73_filtered_output_c0(1);
   bh7_w104_0_c0 <= tile_73_filtered_output_c0(2);
   bh7_w105_0_c0 <= tile_73_filtered_output_c0(3);
   tile_74_X_c0 <= X(52 downto 51);
   tile_74_Y_c0 <= Y(50 downto 48);
   tile_74_mult: IntMultiplierLUT_2x3_Freq800_uid316
      port map ( clk  => clk,
                 X => tile_74_X_c0,
                 Y => tile_74_Y_c0,
                 R => tile_74_output_c0);

   tile_74_filtered_output_c0 <= unsigned(tile_74_output_c0(4 downto 0));
   bh7_w99_5_c0 <= tile_74_filtered_output_c0(0);
   bh7_w100_5_c0 <= tile_74_filtered_output_c0(1);
   bh7_w101_2_c0 <= tile_74_filtered_output_c0(2);
   bh7_w102_3_c0 <= tile_74_filtered_output_c0(3);
   bh7_w103_1_c0 <= tile_74_filtered_output_c0(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq800_uid322_bh7_uid323_In0_c0 <= "" & bh7_w49_4_c0 & "0" & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid323_In1_c0 <= "" & bh7_w50_4_c0 & bh7_w50_5_c0;
   bh7_w49_5_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1(0);
   bh7_w50_6_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1(1);
   bh7_w51_8_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid323: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid323_In0_c0,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid323_In1_c0,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c0);
   Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid323_Out0_copy324_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid327_In0_c0 <= "" & bh7_w51_2_c0 & bh7_w51_5_c0 & bh7_w51_6_c0 & bh7_w51_7_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid327_In1_c0 <= "" & bh7_w52_2_c0;
   bh7_w51_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1(0);
   bh7_w52_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1(1);
   bh7_w53_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid327: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid327_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid327_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid327_Out0_copy328_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid329_In0_c0 <= "" & bh7_w52_5_c0 & bh7_w52_6_c0 & bh7_w52_7_c0 & bh7_w52_8_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid329_In1_c0 <= "" & bh7_w53_2_c0;
   bh7_w52_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1(0);
   bh7_w53_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1(1);
   bh7_w54_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid329: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid329_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid329_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid329_Out0_copy330_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid331_In0_c0 <= "" & bh7_w53_5_c0 & bh7_w53_6_c0 & bh7_w53_7_c0 & bh7_w53_8_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid331_In1_c0 <= "" & bh7_w54_2_c0;
   bh7_w53_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1(0);
   bh7_w54_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1(1);
   bh7_w55_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid331: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid331_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid331_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid331_Out0_copy332_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid335_In0_c0 <= "" & bh7_w54_3_c0 & bh7_w54_6_c0 & bh7_w54_7_c0 & bh7_w54_8_c0 & bh7_w54_9_c0 & bh7_w54_10_c0;
   bh7_w54_13_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1(0);
   bh7_w55_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1(1);
   bh7_w56_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid335: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid335_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid335_Out0_copy336_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid337_In0_c0 <= "" & bh7_w55_2_c0 & bh7_w55_3_c0 & bh7_w55_6_c0 & bh7_w55_7_c0 & bh7_w55_8_c0 & bh7_w55_9_c0;
   bh7_w55_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1(0);
   bh7_w56_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1(1);
   bh7_w57_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid337: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid337_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid337_Out0_copy338_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid339_In0_c0 <= "" & bh7_w56_2_c0 & bh7_w56_5_c0 & bh7_w56_6_c0 & bh7_w56_7_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid339_In1_c0 <= "" & bh7_w57_2_c0;
   bh7_w56_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1(0);
   bh7_w57_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1(1);
   bh7_w58_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid339: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid339_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid339_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid339_Out0_copy340_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid341_In0_c0 <= "" & bh7_w57_3_c0 & bh7_w57_6_c0 & bh7_w57_7_c0 & bh7_w57_8_c0 & bh7_w57_9_c0 & bh7_w57_10_c0;
   bh7_w57_13_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1(0);
   bh7_w58_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1(1);
   bh7_w59_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid341: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid341_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid341_Out0_copy342_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid343_In0_c0 <= "" & bh7_w58_1_c0 & bh7_w58_2_c0 & bh7_w58_6_c0 & bh7_w58_7_c0 & bh7_w58_8_c0 & bh7_w58_9_c0;
   bh7_w58_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1(0);
   bh7_w59_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1(1);
   bh7_w60_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid343: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid343_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid343_Out0_copy344_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid345_In0_c0 <= "" & bh7_w59_1_c0 & bh7_w59_5_c0 & bh7_w59_6_c0 & bh7_w59_7_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid345_In1_c0 <= "" & bh7_w60_1_c0;
   bh7_w59_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1(0);
   bh7_w60_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1(1);
   bh7_w61_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid345: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid345_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid345_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid345_Out0_copy346_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid347_In0_c0 <= "" & bh7_w60_2_c0 & bh7_w60_6_c0 & bh7_w60_7_c0 & bh7_w60_8_c0 & bh7_w60_9_c0 & bh7_w60_10_c0;
   bh7_w60_13_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1(0);
   bh7_w61_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1(1);
   bh7_w62_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid347: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid347_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid347_Out0_copy348_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid349_In0_c0 <= "" & bh7_w61_1_c0 & bh7_w61_2_c0 & bh7_w61_6_c0 & bh7_w61_7_c0 & bh7_w61_8_c0 & bh7_w61_9_c0;
   bh7_w61_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1(0);
   bh7_w62_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1(1);
   bh7_w63_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid349: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid349_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid349_Out0_copy350_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid351_In0_c0 <= "" & bh7_w62_1_c0 & bh7_w62_5_c0 & bh7_w62_6_c0 & bh7_w62_7_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid351_In1_c0 <= "" & bh7_w63_1_c0;
   bh7_w62_11_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1(0);
   bh7_w63_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1(1);
   bh7_w64_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid351: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid351_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid351_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid351_Out0_copy352_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid353_In0_c0 <= "" & bh7_w63_2_c0 & bh7_w63_6_c0 & bh7_w63_7_c0 & bh7_w63_8_c0 & bh7_w63_9_c0 & bh7_w63_10_c0;
   bh7_w63_13_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1(0);
   bh7_w64_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1(1);
   bh7_w65_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid353: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid353_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid353_Out0_copy354_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid355_In0_c0 <= "" & bh7_w64_1_c0 & bh7_w64_2_c0 & bh7_w64_6_c0 & bh7_w64_7_c0 & bh7_w64_8_c0 & bh7_w64_9_c0;
   bh7_w64_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1(0);
   bh7_w65_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1(1);
   bh7_w66_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid355: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid355_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid355_Out0_copy356_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid357_In0_c0 <= "" & bh7_w65_1_c0 & bh7_w65_4_c0 & bh7_w65_5_c0 & bh7_w65_6_c0 & bh7_w65_7_c0 & bh7_w65_8_c0;
   bh7_w65_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1(0);
   bh7_w66_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1(1);
   bh7_w67_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid357: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid357_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid357_Out0_copy358_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid359_In0_c0 <= "" & bh7_w66_1_c0 & bh7_w66_2_c0 & bh7_w66_5_c0 & bh7_w66_6_c0 & bh7_w66_7_c0 & bh7_w66_8_c0;
   bh7_w66_12_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1(0);
   bh7_w67_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1(1);
   bh7_w68_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid359: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid359_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid359_Out0_copy360_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid361_In0_c0 <= "" & bh7_w67_1_c0 & bh7_w67_2_c0 & bh7_w67_5_c0 & bh7_w67_6_c0 & bh7_w67_7_c0 & bh7_w67_8_c0;
   bh7_w67_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1(0);
   bh7_w68_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1(1);
   bh7_w69_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid361: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid361_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid361_Out0_copy362_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid363_In0_c0 <= "" & bh7_w68_1_c0 & bh7_w68_4_c0 & bh7_w68_5_c0 & bh7_w68_6_c0 & bh7_w68_7_c0 & bh7_w68_8_c0;
   bh7_w68_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1(0);
   bh7_w69_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1(1);
   bh7_w70_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid363: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid363_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid363_Out0_copy364_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid365_In0_c0 <= "" & bh7_w69_1_c0 & bh7_w69_2_c0 & bh7_w69_5_c0 & bh7_w69_6_c0 & bh7_w69_7_c0 & bh7_w69_8_c0;
   bh7_w69_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1(0);
   bh7_w70_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1(1);
   bh7_w71_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid365: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid365_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid365_Out0_copy366_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid367_In0_c0 <= "" & bh7_w70_1_c0 & bh7_w70_2_c0 & bh7_w70_5_c0 & bh7_w70_6_c0 & bh7_w70_7_c0 & bh7_w70_8_c0;
   bh7_w70_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1(0);
   bh7_w71_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1(1);
   bh7_w72_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid367: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid367_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid367_Out0_copy368_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid369_In0_c0 <= "" & bh7_w71_1_c0 & bh7_w71_4_c0 & bh7_w71_5_c0 & bh7_w71_6_c0 & bh7_w71_7_c0 & bh7_w71_8_c0;
   bh7_w71_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1(0);
   bh7_w72_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1(1);
   bh7_w73_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid369: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid369_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid369_Out0_copy370_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid371_In0_c0 <= "" & bh7_w72_1_c0 & bh7_w72_2_c0 & bh7_w72_5_c0 & bh7_w72_6_c0 & bh7_w72_7_c0 & bh7_w72_8_c0;
   bh7_w72_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1(0);
   bh7_w73_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1(1);
   bh7_w74_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid371: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid371_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid371_Out0_copy372_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid373_In0_c0 <= "" & bh7_w73_1_c0 & bh7_w73_2_c0 & bh7_w73_5_c0 & bh7_w73_6_c0 & bh7_w73_7_c0 & bh7_w73_8_c0;
   bh7_w73_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1(0);
   bh7_w74_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1(1);
   bh7_w75_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid373: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid373_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid373_Out0_copy374_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid375_In0_c0 <= "" & bh7_w74_1_c0 & bh7_w74_4_c0 & bh7_w74_5_c0 & bh7_w74_6_c0 & bh7_w74_7_c0 & bh7_w74_8_c0;
   bh7_w74_11_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1(0);
   bh7_w75_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1(1);
   bh7_w76_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid375: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid375_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid375_Out0_copy376_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid377_In0_c0 <= "" & bh7_w75_0_c0 & bh7_w75_3_c0 & bh7_w75_4_c0 & bh7_w75_5_c0 & bh7_w75_6_c0 & bh7_w75_7_c0;
   bh7_w75_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1(0);
   bh7_w76_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1(1);
   bh7_w77_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid377: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid377_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid377_Out0_copy378_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid379_In0_c0 <= "" & bh7_w76_0_c0 & bh7_w76_3_c0 & bh7_w76_4_c0 & bh7_w76_5_c0 & bh7_w76_6_c0 & bh7_w76_7_c0;
   bh7_w76_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1(0);
   bh7_w77_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1(1);
   bh7_w78_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid379: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid379_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid379_Out0_copy380_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid381_In0_c0 <= "" & bh7_w77_2_c0 & bh7_w77_3_c0 & bh7_w77_4_c0 & bh7_w77_5_c0 & bh7_w77_6_c0 & bh7_w77_7_c0;
   bh7_w77_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1(0);
   bh7_w78_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1(1);
   bh7_w79_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid381: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid381_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid381_Out0_copy382_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid383_In0_c0 <= "" & bh7_w78_2_c0 & bh7_w78_3_c0 & bh7_w78_4_c0 & bh7_w78_5_c0 & bh7_w78_6_c0 & bh7_w78_7_c0;
   bh7_w78_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1(0);
   bh7_w79_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1(1);
   bh7_w80_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid383: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid383_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid383_Out0_copy384_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid385_In0_c0 <= "" & bh7_w79_2_c0 & bh7_w79_3_c0 & bh7_w79_4_c0 & bh7_w79_5_c0 & bh7_w79_6_c0 & bh7_w79_7_c0;
   bh7_w79_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1(0);
   bh7_w80_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1(1);
   bh7_w81_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid385: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid385_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid385_Out0_copy386_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid387_In0_c0 <= "" & bh7_w80_2_c0 & bh7_w80_3_c0 & bh7_w80_4_c0 & bh7_w80_5_c0 & bh7_w80_6_c0 & bh7_w80_7_c0;
   bh7_w80_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1(0);
   bh7_w81_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1(1);
   bh7_w82_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid387: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid387_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid387_Out0_copy388_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid389_In0_c0 <= "" & bh7_w81_2_c0 & bh7_w81_3_c0 & bh7_w81_4_c0 & bh7_w81_5_c0 & bh7_w81_6_c0 & bh7_w81_7_c0;
   bh7_w81_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1(0);
   bh7_w82_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1(1);
   bh7_w83_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid389: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid389_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid389_Out0_copy390_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid391_In0_c0 <= "" & bh7_w82_1_c0 & bh7_w82_2_c0 & bh7_w82_3_c0 & bh7_w82_4_c0 & bh7_w82_5_c0 & bh7_w82_6_c0;
   bh7_w82_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1(0);
   bh7_w83_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1(1);
   bh7_w84_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid391: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid391_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid391_Out0_copy392_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid393_In0_c0 <= "" & bh7_w83_1_c0 & bh7_w83_2_c0 & bh7_w83_3_c0 & bh7_w83_4_c0 & bh7_w83_5_c0 & bh7_w83_6_c0;
   bh7_w83_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1(0);
   bh7_w84_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1(1);
   bh7_w85_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid393: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid393_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid393_Out0_copy394_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid395_In0_c0 <= "" & bh7_w84_1_c0 & bh7_w84_2_c0 & bh7_w84_3_c0 & bh7_w84_4_c0 & bh7_w84_5_c0 & bh7_w84_6_c0;
   bh7_w84_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1(0);
   bh7_w85_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1(1);
   bh7_w86_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid395: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid395_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid395_Out0_copy396_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid397_In0_c0 <= "" & bh7_w85_1_c0 & bh7_w85_2_c0 & bh7_w85_3_c0 & bh7_w85_4_c0 & bh7_w85_5_c0 & bh7_w85_6_c0;
   bh7_w85_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1(0);
   bh7_w86_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1(1);
   bh7_w87_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid397: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid397_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid397_Out0_copy398_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid401_In0_c0 <= "" & bh7_w86_1_c0 & bh7_w86_2_c0 & bh7_w86_3_c0 & bh7_w86_4_c0 & bh7_w86_5_c0;
   bh7_w86_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1(0);
   bh7_w87_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1(1);
   bh7_w88_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid401: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid401_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid401_Out0_copy402_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid403_In0_c0 <= "" & bh7_w87_1_c0 & bh7_w87_2_c0 & bh7_w87_3_c0 & bh7_w87_4_c0 & bh7_w87_5_c0 & bh7_w87_6_c0;
   bh7_w87_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1(0);
   bh7_w88_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1(1);
   bh7_w89_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid403: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid403_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid403_Out0_copy404_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid405_In0_c0 <= "" & bh7_w88_1_c0 & bh7_w88_2_c0 & bh7_w88_3_c0 & bh7_w88_4_c0 & bh7_w88_5_c0 & bh7_w88_6_c0;
   bh7_w88_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1(0);
   bh7_w89_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1(1);
   bh7_w90_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid405: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid405_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid405_Out0_copy406_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid407_In0_c0 <= "" & bh7_w89_1_c0 & bh7_w89_2_c0 & bh7_w89_3_c0 & bh7_w89_4_c0 & bh7_w89_5_c0;
   bh7_w89_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1(0);
   bh7_w90_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1(1);
   bh7_w91_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid407: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid407_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid407_Out0_copy408_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid409_In0_c0 <= "" & bh7_w90_1_c0 & bh7_w90_2_c0 & bh7_w90_3_c0 & bh7_w90_4_c0 & bh7_w90_5_c0 & bh7_w90_6_c0;
   bh7_w90_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1(0);
   bh7_w91_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1(1);
   bh7_w92_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid409: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid409_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid409_Out0_copy410_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid411_In0_c0 <= "" & bh7_w91_1_c0 & bh7_w91_2_c0 & bh7_w91_3_c0 & bh7_w91_4_c0 & bh7_w91_5_c0 & bh7_w91_6_c0;
   bh7_w91_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1(0);
   bh7_w92_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1(1);
   bh7_w93_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid411: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid411_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid411_Out0_copy412_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid413_In0_c0 <= "" & bh7_w92_1_c0 & bh7_w92_2_c0 & bh7_w92_3_c0 & bh7_w92_4_c0 & bh7_w92_5_c0;
   bh7_w92_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1(0);
   bh7_w93_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1(1);
   bh7_w94_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid413: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid413_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid413_Out0_copy414_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid415_In0_c0 <= "" & bh7_w93_1_c0 & bh7_w93_2_c0 & bh7_w93_3_c0 & bh7_w93_4_c0 & bh7_w93_5_c0 & bh7_w93_6_c0;
   bh7_w93_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1(0);
   bh7_w94_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1(1);
   bh7_w95_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid415: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid415_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid415_Out0_copy416_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid417_In0_c0 <= "" & bh7_w94_1_c0 & bh7_w94_2_c0 & bh7_w94_3_c0 & bh7_w94_4_c0 & bh7_w94_5_c0 & bh7_w94_6_c0;
   bh7_w94_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1(0);
   bh7_w95_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1(1);
   bh7_w96_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid417: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid417_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid417_Out0_copy418_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid419_In0_c0 <= "" & bh7_w95_1_c0 & bh7_w95_2_c0 & bh7_w95_3_c0 & bh7_w95_4_c0 & bh7_w95_5_c0;
   bh7_w95_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1(0);
   bh7_w96_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1(1);
   bh7_w97_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid419: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid419_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid419_Out0_copy420_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid421_In0_c0 <= "" & bh7_w96_1_c0 & bh7_w96_2_c0 & bh7_w96_3_c0 & bh7_w96_4_c0 & bh7_w96_5_c0 & bh7_w96_6_c0;
   bh7_w96_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1(0);
   bh7_w97_9_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1(1);
   bh7_w98_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid421: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid421_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid421_Out0_copy422_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid423_In0_c0 <= "" & bh7_w97_1_c0 & bh7_w97_2_c0 & bh7_w97_3_c0 & bh7_w97_4_c0 & bh7_w97_5_c0 & bh7_w97_6_c0;
   bh7_w97_10_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1(0);
   bh7_w98_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1(1);
   bh7_w99_6_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid423: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid423_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid423_Out0_copy424_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid425_In0_c0 <= "" & bh7_w98_1_c0 & bh7_w98_2_c0 & bh7_w98_3_c0 & bh7_w98_4_c0 & bh7_w98_5_c0;
   bh7_w98_8_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1(0);
   bh7_w99_7_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1(1);
   bh7_w100_6_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1(2);
   Compressor_5_3_Freq800_uid400_uid425: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid425_In0_c0,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c0);
   Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_c1 <= Compressor_5_3_Freq800_uid400_bh7_uid425_Out0_copy426_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid427_In0_c0 <= "" & bh7_w99_0_c0 & bh7_w99_1_c0 & bh7_w99_2_c0 & bh7_w99_3_c0 & bh7_w99_4_c0 & bh7_w99_5_c0;
   bh7_w99_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1(0);
   bh7_w100_7_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1(1);
   bh7_w101_3_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid427: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid427_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid427_Out0_copy428_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid429_In0_c0 <= "" & bh7_w100_0_c0 & bh7_w100_1_c0 & bh7_w100_2_c0 & bh7_w100_3_c0 & bh7_w100_4_c0 & bh7_w100_5_c0;
   bh7_w100_8_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1(0);
   bh7_w101_4_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1(1);
   bh7_w102_4_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1(2);
   Compressor_6_3_Freq800_uid334_uid429: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid429_In0_c0,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c0);
   Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_c1 <= Compressor_6_3_Freq800_uid334_bh7_uid429_Out0_copy430_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid433_In0_c0 <= "" & bh7_w101_0_c0 & bh7_w101_1_c0 & bh7_w101_2_c0;
   bh7_w101_5_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_c1(0);
   bh7_w102_5_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid433: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid433_In0_c0,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c0);
   Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid433_Out0_copy434_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid435_In0_c0 <= "" & bh7_w102_0_c0 & bh7_w102_1_c0 & bh7_w102_2_c0 & bh7_w102_3_c0;
   Compressor_14_3_Freq800_uid326_bh7_uid435_In1_c0 <= "" & bh7_w103_0_c0;
   bh7_w102_6_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1(0);
   bh7_w103_2_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1(1);
   bh7_w104_1_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid435: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid435_In0_c0,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid435_In1_c0,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c0);
   Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid435_Out0_copy436_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid437_In0_c1 <= "" & bh7_w51_9_c1 & bh7_w51_8_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid437_In1_c1 <= "" & bh7_w52_10_c1 & bh7_w52_9_c1;
   bh7_w51_10_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1(0);
   bh7_w52_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1(1);
   bh7_w53_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid437: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid437_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid437_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_copy438_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid437_Out0_copy438_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid439_In0_c1 <= "" & bh7_w53_11_c1 & bh7_w53_10_c1 & bh7_w53_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid439_In1_c1 <= "" & bh7_w54_12_c1 & bh7_w54_11_c1;
   bh7_w53_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1(0);
   bh7_w54_14_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1(1);
   bh7_w55_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid439: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid439_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid439_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_copy440_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid439_Out0_copy440_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid441_In0_c1 <= "" & bh7_w55_10_c1 & bh7_w55_12_c1 & bh7_w55_11_c1;
   bh7_w55_14_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_c1(0);
   bh7_w56_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid441: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid441_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_copy442_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid441_Out0_copy442_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid443_In0_c1 <= "" & bh7_w56_8_c1 & bh7_w56_11_c1 & bh7_w56_10_c1 & bh7_w56_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c0 <= "" & "0";
   bh7_w56_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1(0);
   bh7_w57_14_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1(1);
   bh7_w58_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid443: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid443_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid443_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_copy444_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid443_Out0_copy444_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid445_In0_c1 <= "" & bh7_w57_12_c1 & bh7_w57_13_c1 & bh7_w57_11_c1;
   bh7_w57_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_c1(0);
   bh7_w58_14_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid445: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid445_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_copy446_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid445_Out0_copy446_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid447_In0_c1 <= "" & bh7_w58_10_c1 & bh7_w58_12_c1 & bh7_w58_11_c1;
   bh7_w58_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_c1(0);
   bh7_w59_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid447: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid447_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_copy448_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid447_Out0_copy448_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid449_In0_c1 <= "" & bh7_w59_8_c1 & bh7_w59_11_c1 & bh7_w59_10_c1 & bh7_w59_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c0 <= "" & "0";
   bh7_w59_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1(0);
   bh7_w60_14_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1(1);
   bh7_w61_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid449: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid449_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid449_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_copy450_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid449_Out0_copy450_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid451_In0_c1 <= "" & bh7_w60_12_c1 & bh7_w60_13_c1 & bh7_w60_11_c1;
   bh7_w60_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_c1(0);
   bh7_w61_14_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid451: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid451_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_copy452_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid451_Out0_copy452_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid453_In0_c1 <= "" & bh7_w61_10_c1 & bh7_w61_12_c1 & bh7_w61_11_c1;
   bh7_w61_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_c1(0);
   bh7_w62_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid453: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid453_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_copy454_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid453_Out0_copy454_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid455_In0_c1 <= "" & bh7_w62_8_c1 & bh7_w62_11_c1 & bh7_w62_10_c1 & bh7_w62_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c0 <= "" & "0";
   bh7_w62_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1(0);
   bh7_w63_14_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1(1);
   bh7_w64_13_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid455: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid455_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid455_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_copy456_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid455_Out0_copy456_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid457_In0_c1 <= "" & bh7_w63_12_c1 & bh7_w63_13_c1 & bh7_w63_11_c1;
   bh7_w63_15_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_c1(0);
   bh7_w64_14_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid457: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid457_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_copy458_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid457_Out0_copy458_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid459_In0_c1 <= "" & bh7_w64_10_c1 & bh7_w64_12_c1 & bh7_w64_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid459_In1_c1 <= "" & bh7_w65_11_c1 & bh7_w65_10_c1;
   bh7_w64_15_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1(0);
   bh7_w65_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1(1);
   bh7_w66_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid459: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid459_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid459_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_copy460_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid459_Out0_copy460_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid461_In0_c1 <= "" & bh7_w66_9_c1 & bh7_w66_12_c1 & bh7_w66_11_c1 & bh7_w66_10_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c0 <= "" & "0";
   bh7_w66_14_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1(0);
   bh7_w67_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1(1);
   bh7_w68_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid461: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid461_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid461_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_copy462_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid461_Out0_copy462_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid463_In0_c1 <= "" & bh7_w67_11_c1 & bh7_w67_10_c1 & bh7_w67_9_c1;
   bh7_w67_13_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_c1(0);
   bh7_w68_13_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid463: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid463_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_copy464_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid463_Out0_copy464_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid465_In0_c1 <= "" & bh7_w68_11_c1 & bh7_w68_10_c1 & bh7_w68_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid465_In1_c1 <= "" & bh7_w69_11_c1 & bh7_w69_10_c1;
   bh7_w68_14_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1(0);
   bh7_w69_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1(1);
   bh7_w70_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid465: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid465_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid465_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_copy466_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid465_Out0_copy466_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid467_In0_c1 <= "" & bh7_w70_11_c1 & bh7_w70_10_c1 & bh7_w70_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid467_In1_c1 <= "" & bh7_w71_11_c1 & bh7_w71_10_c1;
   bh7_w70_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1(0);
   bh7_w71_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1(1);
   bh7_w72_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid467: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid467_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid467_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_copy468_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid467_Out0_copy468_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid469_In0_c1 <= "" & bh7_w72_11_c1 & bh7_w72_10_c1 & bh7_w72_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid469_In1_c1 <= "" & bh7_w73_11_c1 & bh7_w73_10_c1;
   bh7_w72_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1(0);
   bh7_w73_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1(1);
   bh7_w74_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid469: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid469_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid469_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_copy470_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid469_Out0_copy470_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid471_In0_c1 <= "" & bh7_w74_11_c1 & bh7_w74_10_c1 & bh7_w74_9_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid471_In1_c1 <= "" & bh7_w75_10_c1 & bh7_w75_9_c1;
   bh7_w74_13_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1(0);
   bh7_w75_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1(1);
   bh7_w76_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid471: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid471_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid471_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_copy472_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid471_Out0_copy472_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid473_In0_c1 <= "" & bh7_w76_10_c1 & bh7_w76_9_c1 & bh7_w76_8_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid473_In1_c1 <= "" & bh7_w77_10_c1 & bh7_w77_9_c1;
   bh7_w76_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1(0);
   bh7_w77_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1(1);
   bh7_w78_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid473: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid473_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid473_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_copy474_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid473_Out0_copy474_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid475_In0_c1 <= "" & bh7_w78_10_c1 & bh7_w78_9_c1 & bh7_w78_8_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid475_In1_c1 <= "" & bh7_w79_10_c1 & bh7_w79_9_c1;
   bh7_w78_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1(0);
   bh7_w79_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1(1);
   bh7_w80_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid475: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid475_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid475_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_copy476_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid475_Out0_copy476_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid477_In0_c1 <= "" & bh7_w80_10_c1 & bh7_w80_9_c1 & bh7_w80_8_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid477_In1_c1 <= "" & bh7_w81_10_c1 & bh7_w81_9_c1;
   bh7_w80_12_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1(0);
   bh7_w81_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1(1);
   bh7_w82_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid477: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid477_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid477_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_copy478_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid477_Out0_copy478_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid479_In0_c1 <= "" & bh7_w82_7_c1 & bh7_w82_10_c1 & bh7_w82_9_c1 & bh7_w82_8_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c0 <= "" & "0";
   bh7_w82_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1(0);
   bh7_w83_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1(1);
   bh7_w84_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid479: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid479_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid479_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_copy480_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid479_Out0_copy480_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid481_In0_c1 <= "" & bh7_w83_9_c1 & bh7_w83_8_c1 & bh7_w83_7_c1;
   bh7_w83_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_c1(0);
   bh7_w84_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid481: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid481_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_copy482_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid481_Out0_copy482_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid483_In0_c1 <= "" & bh7_w84_9_c1 & bh7_w84_8_c1 & bh7_w84_7_c1;
   bh7_w84_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_c1(0);
   bh7_w85_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid483: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid483_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_copy484_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid483_Out0_copy484_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid485_In0_c1 <= "" & bh7_w85_7_c1 & bh7_w85_10_c1 & bh7_w85_9_c1 & bh7_w85_8_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c0 <= "" & "0";
   bh7_w85_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1(0);
   bh7_w86_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1(1);
   bh7_w87_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid485: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid485_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid485_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_copy486_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid485_Out0_copy486_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid487_In0_c1 <= "" & bh7_w86_8_c1 & bh7_w86_7_c1 & bh7_w86_6_c1;
   bh7_w86_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_c1(0);
   bh7_w87_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid487: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid487_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_copy488_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid487_Out0_copy488_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid489_In0_c1 <= "" & bh7_w87_8_c1 & bh7_w87_9_c1 & bh7_w87_7_c1;
   bh7_w87_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_c1(0);
   bh7_w88_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid489: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid489_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_copy490_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid489_Out0_copy490_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid491_In0_c1 <= "" & bh7_w88_7_c1 & bh7_w88_8_c1 & bh7_w88_10_c1 & bh7_w88_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c0 <= "" & "0";
   bh7_w88_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1(0);
   bh7_w89_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1(1);
   bh7_w90_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid491: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid491_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid491_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_copy492_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid491_Out0_copy492_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid493_In0_c1 <= "" & bh7_w89_8_c1 & bh7_w89_7_c1 & bh7_w89_6_c1;
   bh7_w89_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_c1(0);
   bh7_w90_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid493: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid493_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_copy494_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid493_Out0_copy494_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid495_In0_c1 <= "" & bh7_w90_8_c1 & bh7_w90_9_c1 & bh7_w90_7_c1;
   bh7_w90_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_c1(0);
   bh7_w91_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid495: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid495_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_copy496_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid495_Out0_copy496_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid497_In0_c1 <= "" & bh7_w91_7_c1 & bh7_w91_8_c1 & bh7_w91_10_c1 & bh7_w91_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c0 <= "" & "0";
   bh7_w91_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1(0);
   bh7_w92_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1(1);
   bh7_w93_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid497: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid497_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid497_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_copy498_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid497_Out0_copy498_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid499_In0_c1 <= "" & bh7_w92_8_c1 & bh7_w92_7_c1 & bh7_w92_6_c1;
   bh7_w92_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_c1(0);
   bh7_w93_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid499: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid499_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_copy500_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid499_Out0_copy500_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid501_In0_c1 <= "" & bh7_w93_8_c1 & bh7_w93_9_c1 & bh7_w93_7_c1;
   bh7_w93_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_c1(0);
   bh7_w94_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid501: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid501_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_copy502_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid501_Out0_copy502_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid503_In0_c1 <= "" & bh7_w94_7_c1 & bh7_w94_8_c1 & bh7_w94_10_c1 & bh7_w94_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c0 <= "" & "0";
   bh7_w94_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1(0);
   bh7_w95_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1(1);
   bh7_w96_10_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid503: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid503_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid503_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_copy504_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid503_Out0_copy504_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid505_In0_c1 <= "" & bh7_w95_8_c1 & bh7_w95_7_c1 & bh7_w95_6_c1;
   bh7_w95_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_c1(0);
   bh7_w96_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid505: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid505_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_copy506_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid505_Out0_copy506_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid507_In0_c1 <= "" & bh7_w96_8_c1 & bh7_w96_9_c1 & bh7_w96_7_c1;
   bh7_w96_12_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_c1(0);
   bh7_w97_11_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid507: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid507_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_copy508_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid507_Out0_copy508_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid509_In0_c1 <= "" & bh7_w97_7_c1 & bh7_w97_8_c1 & bh7_w97_10_c1 & bh7_w97_9_c1;
   Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c0 <= "" & "0";
   bh7_w97_12_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1(0);
   bh7_w98_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1(1);
   bh7_w99_9_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1(2);
   Compressor_14_3_Freq800_uid326_uid509: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid509_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid509_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_copy510_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_c1 <= Compressor_14_3_Freq800_uid326_bh7_uid509_Out0_copy510_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid511_In0_c1 <= "" & bh7_w98_8_c1 & bh7_w98_7_c1 & bh7_w98_6_c1;
   bh7_w98_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_c1(0);
   bh7_w99_10_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_c1(1);
   Compressor_3_2_Freq800_uid432_uid511: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid511_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_copy512_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_c1 <= Compressor_3_2_Freq800_uid432_bh7_uid511_Out0_copy512_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid513_In0_c1 <= "" & bh7_w99_7_c1 & bh7_w99_8_c1 & bh7_w99_6_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid513_In1_c1 <= "" & bh7_w100_6_c1 & bh7_w100_8_c1;
   bh7_w99_11_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1(0);
   bh7_w100_9_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1(1);
   bh7_w101_6_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid513: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid513_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid513_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_copy514_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid513_Out0_copy514_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid515_In0_c1 <= "" & bh7_w101_5_c1 & bh7_w101_4_c1 & bh7_w101_3_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid515_In1_c1 <= "" & bh7_w102_6_c1 & bh7_w102_5_c1;
   bh7_w101_7_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1(0);
   bh7_w102_7_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1(1);
   bh7_w103_3_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid515: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid515_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid515_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_copy516_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid515_Out0_copy516_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid517_In0_c1 <= "" & bh7_w103_1_c1 & bh7_w103_2_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid517_In1_c1 <= "" & bh7_w104_0_c1 & bh7_w104_1_c1;
   bh7_w103_4_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1(0);
   bh7_w104_2_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1(1);
   bh7_w105_1_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1(2);
   Compressor_23_3_Freq800_uid322_uid517: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid517_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid517_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_copy518_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_c1 <= Compressor_23_3_Freq800_uid322_bh7_uid517_Out0_copy518_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid519_In0_c1 <= "" & bh7_w53_13_c1 & bh7_w53_12_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid519_In1_c1 <= "" & bh7_w54_13_c1 & bh7_w54_14_c1;
   bh7_w53_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2(0);
   bh7_w54_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2(1);
   bh7_w55_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid519: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid519_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid519_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid519_Out0_copy520_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid521_In0_c1 <= "" & bh7_w55_13_c1 & bh7_w55_14_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid521_In1_c1 <= "" & bh7_w56_13_c1 & bh7_w56_12_c1;
   bh7_w55_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2(0);
   bh7_w56_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2(1);
   bh7_w57_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid521: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid521_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid521_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid521_Out0_copy522_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid523_In0_c1 <= "" & bh7_w57_14_c1 & bh7_w57_15_c1 & "0";
   bh7_w57_17_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_c2(0);
   bh7_w58_16_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid523: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid523_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid523_Out0_copy524_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid525_In0_c1 <= "" & bh7_w58_13_c1 & bh7_w58_15_c1 & bh7_w58_14_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid525_In1_c1 <= "" & bh7_w59_13_c1 & bh7_w59_12_c1;
   bh7_w58_17_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2(0);
   bh7_w59_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2(1);
   bh7_w60_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid525: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid525_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid525_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid525_Out0_copy526_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid527_In0_c1 <= "" & bh7_w60_14_c1 & bh7_w60_15_c1 & "0";
   bh7_w60_17_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_c2(0);
   bh7_w61_16_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid527: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid527_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid527_Out0_copy528_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid529_In0_c1 <= "" & bh7_w61_13_c1 & bh7_w61_15_c1 & bh7_w61_14_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid529_In1_c1 <= "" & bh7_w62_13_c1 & bh7_w62_12_c1;
   bh7_w61_17_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2(0);
   bh7_w62_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2(1);
   bh7_w63_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid529: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid529_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid529_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid529_Out0_copy530_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid531_In0_c1 <= "" & bh7_w63_14_c1 & bh7_w63_15_c1 & "0";
   bh7_w63_17_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_c2(0);
   bh7_w64_16_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid531: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid531_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid531_Out0_copy532_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid533_In0_c1 <= "" & bh7_w64_13_c1 & bh7_w64_15_c1 & bh7_w64_14_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid533_In1_c1 <= "" & bh7_w65_9_c1 & bh7_w65_12_c1;
   bh7_w64_17_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2(0);
   bh7_w65_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2(1);
   bh7_w66_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid533: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid533_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid533_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid533_Out0_copy534_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid535_In0_c1 <= "" & bh7_w66_14_c1 & bh7_w66_13_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid535_In1_c1 <= "" & bh7_w67_12_c1 & bh7_w67_13_c1;
   bh7_w66_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2(0);
   bh7_w67_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2(1);
   bh7_w68_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid535: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid535_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid535_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid535_Out0_copy536_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid537_In0_c1 <= "" & bh7_w68_12_c1 & bh7_w68_14_c1 & bh7_w68_13_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid537_In1_c1 <= "" & bh7_w69_9_c1 & bh7_w69_12_c1;
   bh7_w68_16_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2(0);
   bh7_w69_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2(1);
   bh7_w70_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid537: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid537_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid537_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid537_Out0_copy538_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid539_In0_c1 <= "" & bh7_w70_13_c1 & bh7_w70_12_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid539_In1_c1 <= "" & bh7_w71_9_c1 & bh7_w71_12_c1;
   bh7_w70_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2(0);
   bh7_w71_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2(1);
   bh7_w72_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid539: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid539_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid539_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid539_Out0_copy540_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid541_In0_c1 <= "" & bh7_w72_13_c1 & bh7_w72_12_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid541_In1_c1 <= "" & bh7_w73_9_c1 & bh7_w73_12_c1;
   bh7_w72_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2(0);
   bh7_w73_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2(1);
   bh7_w74_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid541: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid541_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid541_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid541_Out0_copy542_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid543_In0_c1 <= "" & bh7_w74_13_c1 & bh7_w74_12_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid543_In1_c1 <= "" & bh7_w75_8_c1 & bh7_w75_11_c1;
   bh7_w74_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2(0);
   bh7_w75_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2(1);
   bh7_w76_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid543: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid543_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid543_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid543_Out0_copy544_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid545_In0_c1 <= "" & bh7_w76_12_c1 & bh7_w76_11_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid545_In1_c1 <= "" & bh7_w77_8_c1 & bh7_w77_11_c1;
   bh7_w76_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2(0);
   bh7_w77_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2(1);
   bh7_w78_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid545: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid545_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid545_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid545_Out0_copy546_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid547_In0_c1 <= "" & bh7_w78_12_c1 & bh7_w78_11_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid547_In1_c1 <= "" & bh7_w79_8_c1 & bh7_w79_11_c1;
   bh7_w78_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2(0);
   bh7_w79_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2(1);
   bh7_w80_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid547: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid547_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid547_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid547_Out0_copy548_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid549_In0_c1 <= "" & bh7_w80_12_c1 & bh7_w80_11_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid549_In1_c1 <= "" & bh7_w81_8_c1 & bh7_w81_11_c1;
   bh7_w80_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2(0);
   bh7_w81_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2(1);
   bh7_w82_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid549: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid549_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid549_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid549_Out0_copy550_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid551_In0_c1 <= "" & bh7_w82_12_c1 & bh7_w82_11_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid551_In1_c1 <= "" & bh7_w83_10_c1 & bh7_w83_11_c1;
   bh7_w82_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2(0);
   bh7_w83_12_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2(1);
   bh7_w84_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid551: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid551_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid551_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid551_Out0_copy552_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid553_In0_c1 <= "" & bh7_w84_10_c1 & bh7_w84_12_c1 & bh7_w84_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid553_In1_c1 <= "" & bh7_w85_12_c1 & bh7_w85_11_c1;
   bh7_w84_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2(0);
   bh7_w85_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2(1);
   bh7_w86_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid553: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid553_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid553_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid553_Out0_copy554_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid555_In0_c1 <= "" & bh7_w86_9_c1 & bh7_w86_10_c1 & "0";
   bh7_w86_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_c2(0);
   bh7_w87_13_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid555: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid555_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid555_Out0_copy556_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid557_In0_c1 <= "" & bh7_w87_10_c1 & bh7_w87_12_c1 & bh7_w87_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid557_In1_c1 <= "" & bh7_w88_12_c1 & bh7_w88_11_c1;
   bh7_w87_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2(0);
   bh7_w88_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2(1);
   bh7_w89_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid557: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid557_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid557_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid557_Out0_copy558_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid559_In0_c1 <= "" & bh7_w89_9_c1 & bh7_w89_10_c1 & "0";
   bh7_w89_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_c2(0);
   bh7_w90_13_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid559: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid559_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid559_Out0_copy560_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid561_In0_c1 <= "" & bh7_w90_10_c1 & bh7_w90_12_c1 & bh7_w90_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid561_In1_c1 <= "" & bh7_w91_12_c1 & bh7_w91_11_c1;
   bh7_w90_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2(0);
   bh7_w91_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2(1);
   bh7_w92_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid561: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid561_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid561_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid561_Out0_copy562_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid563_In0_c1 <= "" & bh7_w92_9_c1 & bh7_w92_10_c1 & "0";
   bh7_w92_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_c2(0);
   bh7_w93_13_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid563: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid563_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid563_Out0_copy564_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid565_In0_c1 <= "" & bh7_w93_10_c1 & bh7_w93_12_c1 & bh7_w93_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid565_In1_c1 <= "" & bh7_w94_12_c1 & bh7_w94_11_c1;
   bh7_w93_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2(0);
   bh7_w94_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2(1);
   bh7_w95_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid565: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid565_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid565_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid565_Out0_copy566_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid567_In0_c1 <= "" & bh7_w95_9_c1 & bh7_w95_10_c1 & "0";
   bh7_w95_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_c2(0);
   bh7_w96_13_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid567: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid567_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid567_Out0_copy568_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid569_In0_c1 <= "" & bh7_w96_10_c1 & bh7_w96_12_c1 & bh7_w96_11_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid569_In1_c1 <= "" & bh7_w97_12_c1 & bh7_w97_11_c1;
   bh7_w96_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2(0);
   bh7_w97_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2(1);
   bh7_w98_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid569: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid569_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid569_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid569_Out0_copy570_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid571_In0_c1 <= "" & bh7_w98_9_c1 & bh7_w98_10_c1 & "0";
   bh7_w98_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_c2(0);
   bh7_w99_12_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_c2(1);
   Compressor_3_2_Freq800_uid432_uid571: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid571_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid571_Out0_copy572_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid573_In0_c1 <= "" & bh7_w99_9_c1 & bh7_w99_11_c1 & bh7_w99_10_c1;
   Compressor_23_3_Freq800_uid322_bh7_uid573_In1_c1 <= "" & bh7_w100_7_c1 & bh7_w100_9_c1;
   bh7_w99_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2(0);
   bh7_w100_10_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2(1);
   bh7_w101_8_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid573: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid573_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid573_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid573_Out0_copy574_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid575_In0_c1 <= "" & bh7_w101_7_c1 & bh7_w101_6_c1 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid575_In1_c1 <= "" & bh7_w102_4_c1 & bh7_w102_7_c1;
   bh7_w101_9_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2(0);
   bh7_w102_8_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2(1);
   bh7_w103_5_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid575: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid575_In0_c1,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid575_In1_c1,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c1);
   Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid575_Out0_copy576_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid577_In0_c1 <= "" & bh7_w103_4_c1 & bh7_w103_3_c1 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid577_In1_c1 <= "" & bh7_w104_2_c1;
   bh7_w103_6_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2(0);
   bh7_w104_3_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2(1);
   bh7_w105_2_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid577: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid577_In0_c1,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid577_In1_c1,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c1);
   Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid577_Out0_copy578_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid579_In0_c1 <= "" & bh7_w105_0_c1 & bh7_w105_1_c1 & "0";
   bh7_w105_3_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_c2(0);
   Compressor_3_2_Freq800_uid432_uid579: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid579_In0_c1,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c1);
   Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_c2 <= Compressor_3_2_Freq800_uid432_bh7_uid579_Out0_copy580_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid581_In0_c2 <= "" & bh7_w55_16_c2 & bh7_w55_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid581_In1_c2 <= "" & bh7_w56_14_c2;
   bh7_w55_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2(0);
   bh7_w56_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2(1);
   bh7_w57_18_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid581: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid581_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid581_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_copy582_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid581_Out0_copy582_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid583_In0_c2 <= "" & bh7_w57_16_c2 & bh7_w57_17_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid583_In1_c2 <= "" & bh7_w58_16_c2 & bh7_w58_17_c2;
   bh7_w57_19_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2(0);
   bh7_w58_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2(1);
   bh7_w59_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid583: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid583_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid583_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_copy584_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid583_Out0_copy584_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid585_In0_c2 <= "" & bh7_w60_16_c2 & bh7_w60_17_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid585_In1_c2 <= "" & bh7_w61_16_c2 & bh7_w61_17_c2;
   bh7_w60_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2(0);
   bh7_w61_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2(1);
   bh7_w62_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid585: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid585_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid585_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_copy586_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid585_Out0_copy586_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid587_In0_c2 <= "" & bh7_w63_16_c2 & bh7_w63_17_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid587_In1_c2 <= "" & bh7_w64_16_c2 & bh7_w64_17_c2;
   bh7_w63_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2(0);
   bh7_w64_18_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2(1);
   bh7_w65_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid587: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid587_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid587_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_copy588_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid587_Out0_copy588_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid589_In0_c2 <= "" & bh7_w66_15_c2 & bh7_w66_16_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid589_In1_c2 <= "" & bh7_w67_14_c2;
   bh7_w66_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2(0);
   bh7_w67_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2(1);
   bh7_w68_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid589: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid589_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid589_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_copy590_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid589_Out0_copy590_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid591_In0_c2 <= "" & bh7_w68_15_c2 & bh7_w68_16_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid591_In1_c2 <= "" & bh7_w69_13_c2;
   bh7_w68_18_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2(0);
   bh7_w69_14_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2(1);
   bh7_w70_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid591: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid591_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid591_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_copy592_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid591_Out0_copy592_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid593_In0_c2 <= "" & bh7_w70_14_c2 & bh7_w70_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid593_In1_c2 <= "" & bh7_w71_13_c2;
   bh7_w70_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2(0);
   bh7_w71_14_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2(1);
   bh7_w72_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid593: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid593_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid593_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_copy594_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid593_Out0_copy594_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid595_In0_c2 <= "" & bh7_w72_15_c2 & bh7_w72_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid595_In1_c2 <= "" & bh7_w73_13_c2;
   bh7_w72_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2(0);
   bh7_w73_14_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2(1);
   bh7_w74_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid595: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid595_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid595_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_copy596_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid595_Out0_copy596_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid597_In0_c2 <= "" & bh7_w74_15_c2 & bh7_w74_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid597_In1_c2 <= "" & bh7_w75_12_c2;
   bh7_w74_17_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2(0);
   bh7_w75_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2(1);
   bh7_w76_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid597: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid597_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid597_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_copy598_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid597_Out0_copy598_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid599_In0_c2 <= "" & bh7_w76_14_c2 & bh7_w76_13_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid599_In1_c2 <= "" & bh7_w77_12_c2;
   bh7_w76_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2(0);
   bh7_w77_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2(1);
   bh7_w78_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid599: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid599_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid599_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_copy600_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid599_Out0_copy600_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid601_In0_c2 <= "" & bh7_w78_14_c2 & bh7_w78_13_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid601_In1_c2 <= "" & bh7_w79_12_c2;
   bh7_w78_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2(0);
   bh7_w79_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2(1);
   bh7_w80_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid601: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid601_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid601_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_copy602_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid601_Out0_copy602_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid603_In0_c2 <= "" & bh7_w80_14_c2 & bh7_w80_13_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid603_In1_c2 <= "" & bh7_w81_12_c2;
   bh7_w80_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2(0);
   bh7_w81_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2(1);
   bh7_w82_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid603: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid603_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid603_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_copy604_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid603_Out0_copy604_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid605_In0_c2 <= "" & bh7_w82_14_c2 & bh7_w82_13_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid605_In1_c2 <= "" & bh7_w83_12_c2;
   bh7_w82_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2(0);
   bh7_w83_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2(1);
   bh7_w84_15_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid605: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid605_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid605_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_copy606_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid605_Out0_copy606_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid607_In0_c2 <= "" & bh7_w84_13_c2 & bh7_w84_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid607_In1_c2 <= "" & bh7_w85_13_c2;
   bh7_w84_16_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2(0);
   bh7_w85_14_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2(1);
   bh7_w86_13_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid607: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid607_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid607_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_copy608_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid607_Out0_copy608_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid609_In0_c2 <= "" & bh7_w86_11_c2 & bh7_w86_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid609_In1_c2 <= "" & bh7_w87_13_c2 & bh7_w87_14_c2;
   bh7_w86_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2(0);
   bh7_w87_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2(1);
   bh7_w88_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid609: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid609_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid609_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_copy610_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid609_Out0_copy610_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid611_In0_c2 <= "" & bh7_w89_11_c2 & bh7_w89_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid611_In1_c2 <= "" & bh7_w90_13_c2 & bh7_w90_14_c2;
   bh7_w89_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2(0);
   bh7_w90_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2(1);
   bh7_w91_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid611: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid611_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid611_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_copy612_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid611_Out0_copy612_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid613_In0_c2 <= "" & bh7_w92_11_c2 & bh7_w92_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid613_In1_c2 <= "" & bh7_w93_13_c2 & bh7_w93_14_c2;
   bh7_w92_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2(0);
   bh7_w93_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2(1);
   bh7_w94_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid613: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid613_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid613_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_copy614_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid613_Out0_copy614_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid615_In0_c2 <= "" & bh7_w95_11_c2 & bh7_w95_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid615_In1_c2 <= "" & bh7_w96_13_c2 & bh7_w96_14_c2;
   bh7_w95_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2(0);
   bh7_w96_15_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2(1);
   bh7_w97_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid615: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid615_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid615_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_copy616_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid615_Out0_copy616_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid617_In0_c2 <= "" & bh7_w98_11_c2 & bh7_w98_12_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid617_In1_c2 <= "" & bh7_w99_12_c2 & bh7_w99_13_c2;
   bh7_w98_13_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2(0);
   bh7_w99_14_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2(1);
   bh7_w100_11_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2(2);
   Compressor_23_3_Freq800_uid322_uid617: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid617_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid617_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_copy618_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_c2 <= Compressor_23_3_Freq800_uid322_bh7_uid617_Out0_copy618_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid619_In0_c2 <= "" & bh7_w101_8_c2 & bh7_w101_9_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid619_In1_c2 <= "" & bh7_w102_8_c2;
   bh7_w101_10_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2(0);
   bh7_w102_9_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2(1);
   bh7_w103_7_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid619: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid619_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid619_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_copy620_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid619_Out0_copy620_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid621_In0_c2 <= "" & bh7_w103_6_c2 & bh7_w103_5_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid621_In1_c2 <= "" & bh7_w104_3_c2;
   bh7_w103_8_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2(0);
   bh7_w104_4_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2(1);
   bh7_w105_4_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2(2);
   Compressor_14_3_Freq800_uid326_uid621: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid621_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid621_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_copy622_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid621_Out0_copy622_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid623_In0_c2 <= "" & bh7_w105_3_c2 & bh7_w105_2_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c0 <= "" & "0";
   bh7_w105_5_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_c2(0);
   Compressor_14_3_Freq800_uid326_uid623: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid623_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid623_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_copy624_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_c2 <= Compressor_14_3_Freq800_uid326_bh7_uid623_Out0_copy624_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid625_In0_c2 <= "" & bh7_w57_18_c2 & bh7_w57_19_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid625_In1_c2 <= "" & bh7_w58_18_c2;
   bh7_w57_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3(0);
   bh7_w58_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3(1);
   bh7_w59_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid625: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid625_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid625_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid625_Out0_copy626_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid627_In0_c2 <= "" & bh7_w59_14_c2 & bh7_w59_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid627_In1_c2 <= "" & bh7_w60_18_c2;
   bh7_w59_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3(0);
   bh7_w60_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3(1);
   bh7_w61_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid627: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid627_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid627_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid627_Out0_copy628_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid629_In0_c2 <= "" & bh7_w62_14_c2 & bh7_w62_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid629_In1_c2 <= "" & bh7_w63_18_c2;
   bh7_w62_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3(0);
   bh7_w63_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3(1);
   bh7_w64_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid629: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid629_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid629_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid629_Out0_copy630_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid631_In0_c2 <= "" & bh7_w65_13_c2 & bh7_w65_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid631_In1_c2 <= "" & bh7_w66_17_c2;
   bh7_w65_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3(0);
   bh7_w66_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3(1);
   bh7_w67_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid631: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid631_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid631_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid631_Out0_copy632_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid633_In0_c2 <= "" & bh7_w68_17_c2 & bh7_w68_18_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid633_In1_c2 <= "" & bh7_w69_14_c2;
   bh7_w68_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3(0);
   bh7_w69_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3(1);
   bh7_w70_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid633: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid633_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid633_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid633_Out0_copy634_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid635_In0_c2 <= "" & bh7_w70_16_c2 & bh7_w70_17_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid635_In1_c2 <= "" & bh7_w71_14_c2;
   bh7_w70_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3(0);
   bh7_w71_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3(1);
   bh7_w72_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid635: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid635_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid635_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid635_Out0_copy636_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid637_In0_c2 <= "" & bh7_w72_16_c2 & bh7_w72_17_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid637_In1_c2 <= "" & bh7_w73_14_c2;
   bh7_w72_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3(0);
   bh7_w73_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3(1);
   bh7_w74_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid637: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid637_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid637_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid637_Out0_copy638_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid639_In0_c2 <= "" & bh7_w74_17_c2 & bh7_w74_16_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid639_In1_c2 <= "" & bh7_w75_13_c2;
   bh7_w74_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3(0);
   bh7_w75_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3(1);
   bh7_w76_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid639: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid639_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid639_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid639_Out0_copy640_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid641_In0_c2 <= "" & bh7_w76_16_c2 & bh7_w76_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid641_In1_c2 <= "" & bh7_w77_13_c2;
   bh7_w76_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3(0);
   bh7_w77_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3(1);
   bh7_w78_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid641: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid641_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid641_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid641_Out0_copy642_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid643_In0_c2 <= "" & bh7_w78_16_c2 & bh7_w78_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid643_In1_c2 <= "" & bh7_w79_13_c2;
   bh7_w78_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3(0);
   bh7_w79_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3(1);
   bh7_w80_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid643: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid643_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid643_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid643_Out0_copy644_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid645_In0_c2 <= "" & bh7_w80_16_c2 & bh7_w80_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid645_In1_c2 <= "" & bh7_w81_13_c2;
   bh7_w80_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3(0);
   bh7_w81_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3(1);
   bh7_w82_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid645: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid645_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid645_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid645_Out0_copy646_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid647_In0_c2 <= "" & bh7_w82_16_c2 & bh7_w82_15_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid647_In1_c2 <= "" & bh7_w83_13_c2;
   bh7_w82_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3(0);
   bh7_w83_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3(1);
   bh7_w84_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid647: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid647_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid647_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid647_Out0_copy648_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid649_In0_c2 <= "" & bh7_w84_15_c2 & bh7_w84_16_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid649_In1_c2 <= "" & bh7_w85_14_c2;
   bh7_w84_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3(0);
   bh7_w85_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3(1);
   bh7_w86_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid649: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid649_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid649_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid649_Out0_copy650_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid651_In0_c2 <= "" & bh7_w86_13_c2 & bh7_w86_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid651_In1_c2 <= "" & bh7_w87_15_c2;
   bh7_w86_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3(0);
   bh7_w87_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3(1);
   bh7_w88_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid651: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid651_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid651_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid651_Out0_copy652_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid653_In0_c2 <= "" & bh7_w88_13_c2 & bh7_w88_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid653_In1_c2 <= "" & bh7_w89_13_c2;
   bh7_w88_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3(0);
   bh7_w89_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3(1);
   bh7_w90_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid653: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid653_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid653_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid653_Out0_copy654_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid655_In0_c2 <= "" & bh7_w91_13_c2 & bh7_w91_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid655_In1_c2 <= "" & bh7_w92_13_c2;
   bh7_w91_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3(0);
   bh7_w92_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3(1);
   bh7_w93_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid655: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid655_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid655_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid655_Out0_copy656_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid657_In0_c2 <= "" & bh7_w94_13_c2 & bh7_w94_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid657_In1_c2 <= "" & bh7_w95_13_c2;
   bh7_w94_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3(0);
   bh7_w95_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3(1);
   bh7_w96_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid657: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid657_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid657_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid657_Out0_copy658_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid659_In0_c2 <= "" & bh7_w97_13_c2 & bh7_w97_14_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid659_In1_c2 <= "" & bh7_w98_13_c2;
   bh7_w97_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3(0);
   bh7_w98_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3(1);
   bh7_w99_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid659: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid659_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid659_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid659_Out0_copy660_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid661_In0_c2 <= "" & bh7_w100_10_c2 & bh7_w100_11_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid661_In1_c2 <= "" & bh7_w101_10_c2;
   bh7_w100_12_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3(0);
   bh7_w101_11_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3(1);
   bh7_w102_10_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid661: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid661_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid661_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid661_Out0_copy662_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid663_In0_c2 <= "" & bh7_w103_7_c2 & bh7_w103_8_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid663_In1_c2 <= "" & bh7_w104_4_c2;
   bh7_w103_9_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3(0);
   bh7_w104_5_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3(1);
   bh7_w105_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid663: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid663_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid663_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid663_Out0_copy664_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid665_In0_c2 <= "" & bh7_w105_5_c2 & bh7_w105_4_c2 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c0 <= "" & "0";
   bh7_w105_7_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_c3(0);
   Compressor_14_3_Freq800_uid326_uid665: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid665_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid665_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid665_Out0_copy666_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid667_In0_c2 <= "" & bh7_w17_0_c2 & bh7_w17_1_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid667_In1_c2 <= "" & bh7_w18_0_c2 & bh7_w18_1_c2;
   bh7_w17_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3(0);
   bh7_w18_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3(1);
   bh7_w19_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid667: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid667_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid667_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid667_Out0_copy668_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid669_In0_c2 <= "" & bh7_w19_0_c2 & bh7_w19_1_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid669_In1_c2 <= "" & bh7_w20_0_c2 & bh7_w20_1_c2;
   bh7_w19_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3(0);
   bh7_w20_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3(1);
   bh7_w21_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid669: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid669_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid669_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid669_Out0_copy670_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid671_In0_c2 <= "" & bh7_w21_0_c2 & bh7_w21_1_c2 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid671_In1_c2 <= "" & bh7_w22_0_c2 & bh7_w22_1_c2;
   bh7_w21_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3(0);
   bh7_w22_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3(1);
   bh7_w23_2_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid671: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid671_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid671_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid671_Out0_copy672_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid673_In0_c2 <= "" & bh7_w23_0_c2 & bh7_w23_1_c2 & "0";
   bh7_w23_3_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_c3(0);
   bh7_w24_3_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid673: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid673_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid673_Out0_copy674_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid675_In0_c2 <= "" & bh7_w24_0_c2 & bh7_w24_1_c2 & bh7_w24_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid675_In1_c2 <= "" & bh7_w25_0_c2 & bh7_w25_1_c2;
   bh7_w24_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3(0);
   bh7_w25_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3(1);
   bh7_w26_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid675: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid675_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid675_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid675_Out0_copy676_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid677_In0_c2 <= "" & bh7_w26_0_c2 & bh7_w26_1_c2 & bh7_w26_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid677_In1_c2 <= "" & bh7_w27_0_c2 & bh7_w27_1_c2;
   bh7_w26_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3(0);
   bh7_w27_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3(1);
   bh7_w28_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid677: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid677_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid677_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid677_Out0_copy678_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid679_In0_c2 <= "" & bh7_w28_0_c2 & bh7_w28_1_c2 & bh7_w28_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid679_In1_c2 <= "" & bh7_w29_0_c2 & bh7_w29_1_c2;
   bh7_w28_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3(0);
   bh7_w29_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3(1);
   bh7_w30_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid679: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid679_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid679_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid679_Out0_copy680_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid681_In0_c2 <= "" & bh7_w30_0_c2 & bh7_w30_1_c2 & bh7_w30_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid681_In1_c2 <= "" & bh7_w31_0_c2 & bh7_w31_1_c2;
   bh7_w30_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3(0);
   bh7_w31_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3(1);
   bh7_w32_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid681: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid681_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid681_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid681_Out0_copy682_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid683_In0_c2 <= "" & bh7_w32_0_c2 & bh7_w32_1_c2 & bh7_w32_2_c2;
   Compressor_23_3_Freq800_uid322_bh7_uid683_In1_c2 <= "" & bh7_w33_0_c2 & bh7_w33_1_c2;
   bh7_w32_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3(0);
   bh7_w33_3_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3(1);
   bh7_w34_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid683: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid683_In0_c2,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid683_In1_c2,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c2);
   Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid683_Out0_copy684_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid685_In0_c2 <= "" & bh7_w34_0_c2 & bh7_w34_1_c2 & bh7_w34_2_c2 & bh7_w34_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid685_In1_c2 <= "" & bh7_w35_0_c2;
   bh7_w34_5_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3(0);
   bh7_w35_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3(1);
   bh7_w36_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid685: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid685_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid685_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid685_Out0_copy686_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid687_In0_c2 <= "" & bh7_w35_1_c2 & bh7_w35_2_c2 & bh7_w35_3_c2;
   bh7_w35_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_c3(0);
   bh7_w36_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid687: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid687_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid687_Out0_copy688_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid689_In0_c2 <= "" & bh7_w36_0_c2 & bh7_w36_1_c2 & bh7_w36_2_c2 & bh7_w36_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid689_In1_c2 <= "" & bh7_w37_0_c2;
   bh7_w36_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3(0);
   bh7_w37_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3(1);
   bh7_w38_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid689: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid689_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid689_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid689_Out0_copy690_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid691_In0_c2 <= "" & bh7_w37_1_c2 & bh7_w37_2_c2 & bh7_w37_3_c2;
   bh7_w37_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_c3(0);
   bh7_w38_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid691: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid691_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid691_Out0_copy692_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid693_In0_c2 <= "" & bh7_w38_0_c2 & bh7_w38_1_c2 & bh7_w38_2_c2 & bh7_w38_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid693_In1_c2 <= "" & bh7_w39_0_c2;
   bh7_w38_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3(0);
   bh7_w39_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3(1);
   bh7_w40_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid693: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid693_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid693_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid693_Out0_copy694_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid695_In0_c2 <= "" & bh7_w39_1_c2 & bh7_w39_2_c2 & bh7_w39_3_c2;
   bh7_w39_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_c3(0);
   bh7_w40_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid695: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid695_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid695_Out0_copy696_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid697_In0_c2 <= "" & bh7_w40_0_c2 & bh7_w40_1_c2 & bh7_w40_2_c2 & bh7_w40_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid697_In1_c2 <= "" & bh7_w41_0_c2;
   bh7_w40_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3(0);
   bh7_w41_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3(1);
   bh7_w42_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid697: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid697_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid697_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid697_Out0_copy698_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid699_In0_c2 <= "" & bh7_w41_1_c2 & bh7_w41_2_c2 & bh7_w41_3_c2;
   bh7_w41_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_c3(0);
   bh7_w42_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid699: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid699_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid699_Out0_copy700_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid701_In0_c2 <= "" & bh7_w42_0_c2 & bh7_w42_1_c2 & bh7_w42_2_c2 & bh7_w42_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid701_In1_c2 <= "" & bh7_w43_0_c2;
   bh7_w42_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3(0);
   bh7_w43_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3(1);
   bh7_w44_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid701: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid701_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid701_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid701_Out0_copy702_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid703_In0_c2 <= "" & bh7_w43_1_c2 & bh7_w43_2_c2 & bh7_w43_3_c2;
   bh7_w43_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_c3(0);
   bh7_w44_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid703: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid703_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid703_Out0_copy704_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid705_In0_c2 <= "" & bh7_w44_0_c2 & bh7_w44_1_c2 & bh7_w44_2_c2 & bh7_w44_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid705_In1_c2 <= "" & bh7_w45_0_c2;
   bh7_w44_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3(0);
   bh7_w45_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3(1);
   bh7_w46_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid705: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid705_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid705_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid705_Out0_copy706_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid707_In0_c2 <= "" & bh7_w45_1_c2 & bh7_w45_2_c2 & bh7_w45_3_c2;
   bh7_w45_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_c3(0);
   bh7_w46_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid707: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid707_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid707_Out0_copy708_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid709_In0_c2 <= "" & bh7_w46_0_c2 & bh7_w46_1_c2 & bh7_w46_2_c2 & bh7_w46_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid709_In1_c2 <= "" & bh7_w47_0_c2;
   bh7_w46_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3(0);
   bh7_w47_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3(1);
   bh7_w48_5_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid709: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid709_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid709_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid709_Out0_copy710_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid711_In0_c2 <= "" & bh7_w47_1_c2 & bh7_w47_2_c2 & bh7_w47_3_c2;
   bh7_w47_5_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_c3(0);
   bh7_w48_6_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid711: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid711_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid711_Out0_copy712_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid713_In0_c2 <= "" & bh7_w48_4_c2 & bh7_w48_0_c2 & bh7_w48_1_c2 & bh7_w48_2_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c1 <= "" & bh7_w49_5_c1;
   bh7_w48_7_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3(0);
   bh7_w49_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3(1);
   bh7_w50_7_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid713: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid713_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid713_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid713_Out0_copy714_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid715_In0_c2 <= "" & bh7_w49_0_c2 & bh7_w49_1_c2 & bh7_w49_2_c2 & bh7_w49_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c1 <= "" & bh7_w50_6_c1;
   bh7_w49_7_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3(0);
   bh7_w50_8_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3(1);
   bh7_w51_11_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid715: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid715_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid715_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid715_Out0_copy716_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid717_In0_c2 <= "" & bh7_w50_0_c2 & bh7_w50_1_c2 & bh7_w50_2_c2 & bh7_w50_3_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c1 <= "" & bh7_w51_10_c1;
   bh7_w50_9_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3(0);
   bh7_w51_12_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3(1);
   bh7_w52_12_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid717: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid717_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid717_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid717_Out0_copy718_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid719_In0_c2 <= "" & bh7_w51_0_c2 & bh7_w51_1_c2 & bh7_w51_3_c2 & bh7_w51_4_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c1 <= "" & bh7_w52_11_c1;
   bh7_w51_13_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3(0);
   bh7_w52_13_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3(1);
   bh7_w53_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid719: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid719_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid719_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid719_Out0_copy720_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid721_In0_c2 <= "" & bh7_w52_0_c2 & bh7_w52_1_c2 & bh7_w52_3_c2 & bh7_w52_4_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid721_In1_c2 <= "" & bh7_w53_14_c2;
   bh7_w52_14_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3(0);
   bh7_w53_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3(1);
   bh7_w54_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid721: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid721_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid721_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid721_Out0_copy722_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid723_In0_c2 <= "" & bh7_w53_0_c2 & bh7_w53_1_c2 & bh7_w53_3_c2 & bh7_w53_4_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid723_In1_c2 <= "" & bh7_w54_15_c2;
   bh7_w53_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3(0);
   bh7_w54_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3(1);
   bh7_w55_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid723: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid723_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid723_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid723_Out0_copy724_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid725_In0_c2 <= "" & bh7_w54_0_c2 & bh7_w54_1_c2 & bh7_w54_4_c2 & bh7_w54_5_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid725_In1_c2 <= "" & bh7_w55_17_c2;
   bh7_w54_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3(0);
   bh7_w55_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3(1);
   bh7_w56_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid725: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid725_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid725_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid725_Out0_copy726_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid727_In0_c2 <= "" & bh7_w55_0_c2 & bh7_w55_1_c2 & bh7_w55_4_c2 & bh7_w55_5_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid727_In1_c2 <= "" & bh7_w56_15_c2;
   bh7_w55_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3(0);
   bh7_w56_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3(1);
   bh7_w57_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid727: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid727_In0_c2,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid727_In1_c2,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c2);
   Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid727_Out0_copy728_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c2 <= "" & bh7_w56_0_c2 & bh7_w56_1_c2 & bh7_w56_3_c2 & bh7_w56_4_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid729_In1_c3 <= "" & bh7_w57_20_c3;
   bh7_w56_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3(0);
   bh7_w57_22_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3(1);
   bh7_w58_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid729: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid729_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid729_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_copy730_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid729_Out0_copy730_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c2 <= "" & bh7_w57_0_c2 & bh7_w57_1_c2 & bh7_w57_4_c2 & bh7_w57_5_c2;
   Compressor_14_3_Freq800_uid326_bh7_uid731_In1_c3 <= "" & bh7_w58_19_c3;
   bh7_w57_23_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3(0);
   bh7_w58_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3(1);
   bh7_w59_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid731: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid731_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid731_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_copy732_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid731_Out0_copy732_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid733_In0_c2 <= "" & bh7_w58_0_c2 & bh7_w58_3_c2 & bh7_w58_4_c2;
   bh7_w58_22_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_c3(0);
   bh7_w59_19_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid733: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid733_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid733_Out0_copy734_c3; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid735_In0_c3 <= "" & bh7_w59_16_c3 & bh7_w59_17_c3 & bh7_w59_0_c3 & bh7_w59_2_c3 & bh7_w59_3_c3 & bh7_w59_4_c3;
   bh7_w59_20_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3(0);
   bh7_w60_20_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3(1);
   bh7_w61_20_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3(2);
   Compressor_6_3_Freq800_uid334_uid735: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid735_In0_c3,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_copy736_c3);
   Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid735_Out0_copy736_c3; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq800_uid400_bh7_uid737_In0_c3 <= "" & bh7_w60_19_c3 & bh7_w60_0_c3 & bh7_w60_3_c3 & bh7_w60_4_c3 & bh7_w60_5_c3;
   bh7_w60_21_c3 <= Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3(0);
   bh7_w61_21_c3 <= Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3(1);
   bh7_w62_17_c3 <= Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3(2);
   Compressor_5_3_Freq800_uid400_uid737: Compressor_5_3_Freq800_uid400
      port map ( X0 => Compressor_5_3_Freq800_uid400_bh7_uid737_In0_c3,
                 R => Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_copy738_c3);
   Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_c3 <= Compressor_5_3_Freq800_uid400_bh7_uid737_Out0_copy738_c3; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid739_In0_c3 <= "" & bh7_w61_18_c3 & bh7_w61_19_c3 & bh7_w61_0_c3 & bh7_w61_3_c3 & bh7_w61_4_c3 & bh7_w61_5_c3;
   bh7_w61_22_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3(0);
   bh7_w62_18_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3(1);
   bh7_w63_20_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3(2);
   Compressor_6_3_Freq800_uid334_uid739: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid739_In0_c3,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_copy740_c3);
   Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid739_Out0_copy740_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid741_In0_c3 <= "" & bh7_w62_16_c3 & bh7_w62_0_c3 & bh7_w62_2_c3 & bh7_w62_3_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid741_In1_c3 <= "" & bh7_w63_19_c3;
   bh7_w62_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3(0);
   bh7_w63_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3(1);
   bh7_w64_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid741: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid741_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid741_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_copy742_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid741_Out0_copy742_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid743_In0_c2 <= "" & bh7_w63_0_c2 & bh7_w63_3_c2 & bh7_w63_4_c2;
   bh7_w63_22_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_c3(0);
   bh7_w64_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid743: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid743_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid743_Out0_copy744_c3; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq800_uid334_bh7_uid745_In0_c3 <= "" & bh7_w64_18_c3 & bh7_w64_19_c3 & bh7_w64_0_c3 & bh7_w64_3_c3 & bh7_w64_4_c3 & bh7_w64_5_c3;
   bh7_w64_22_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3(0);
   bh7_w65_16_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3(1);
   bh7_w66_19_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3(2);
   Compressor_6_3_Freq800_uid334_uid745: Compressor_6_3_Freq800_uid334
      port map ( X0 => Compressor_6_3_Freq800_uid334_bh7_uid745_In0_c3,
                 R => Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_copy746_c3);
   Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_c3 <= Compressor_6_3_Freq800_uid334_bh7_uid745_Out0_copy746_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid747_In0_c3 <= "" & bh7_w65_15_c3 & bh7_w65_0_c3 & bh7_w65_2_c3 & bh7_w65_3_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid747_In1_c3 <= "" & bh7_w66_18_c3;
   bh7_w65_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3(0);
   bh7_w66_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3(1);
   bh7_w67_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid747: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid747_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid747_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_copy748_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid747_Out0_copy748_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid749_In0_c2 <= "" & bh7_w66_0_c2 & bh7_w66_3_c2 & bh7_w66_4_c2;
   bh7_w66_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_c3(0);
   bh7_w67_18_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid749: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid749_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid749_Out0_copy750_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid751_In0_c3 <= "" & bh7_w67_15_c3 & bh7_w67_16_c3 & bh7_w67_0_c3 & bh7_w67_3_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid751_In1_c3 <= "" & bh7_w68_19_c3;
   bh7_w67_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3(0);
   bh7_w68_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3(1);
   bh7_w69_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid751: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid751_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid751_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_copy752_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid751_Out0_copy752_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid753_In0_c2 <= "" & bh7_w68_0_c2 & bh7_w68_2_c2 & bh7_w68_3_c2;
   bh7_w68_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_c3(0);
   bh7_w69_17_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid753: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid753_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid753_Out0_copy754_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid755_In0_c3 <= "" & bh7_w69_15_c3 & bh7_w69_0_c3 & bh7_w69_3_c3 & bh7_w69_4_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid755_In1_c3 <= "" & bh7_w70_18_c3;
   bh7_w69_18_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3(0);
   bh7_w70_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3(1);
   bh7_w71_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid755: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid755_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid755_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_copy756_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid755_Out0_copy756_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid757_In0_c3 <= "" & bh7_w70_19_c3 & bh7_w70_0_c3 & bh7_w70_3_c3 & bh7_w70_4_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid757_In1_c3 <= "" & bh7_w71_15_c3;
   bh7_w70_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3(0);
   bh7_w71_17_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3(1);
   bh7_w72_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid757: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid757_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid757_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_copy758_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid757_Out0_copy758_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid759_In0_c2 <= "" & bh7_w71_0_c2 & bh7_w71_2_c2 & bh7_w71_3_c2;
   bh7_w71_18_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_c3(0);
   bh7_w72_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid759: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid759_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid759_Out0_copy760_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid761_In0_c3 <= "" & bh7_w72_18_c3 & bh7_w72_19_c3 & bh7_w72_0_c3 & bh7_w72_3_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid761_In1_c3 <= "" & bh7_w73_15_c3;
   bh7_w72_22_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3(0);
   bh7_w73_16_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3(1);
   bh7_w74_20_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid761: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid761_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid761_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_copy762_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid761_Out0_copy762_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid763_In0_c2 <= "" & bh7_w73_0_c2 & bh7_w73_3_c2 & bh7_w73_4_c2;
   bh7_w73_17_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_c3(0);
   bh7_w74_21_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid763: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid763_In0_c2,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c2);
   Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid763_Out0_copy764_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid765_In0_c3 <= "" & bh7_w74_18_c3 & bh7_w74_0_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c2 <= "" & bh7_w75_1_c2;
   bh7_w74_22_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3(0);
   bh7_w75_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3(1);
   bh7_w76_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid765: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid765_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid765_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_copy766_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid765_Out0_copy766_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid767_In0_c3 <= "" & bh7_w74_2_c3 & bh7_w74_3_c3 & bh7_w74_19_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid767_In1_c3 <= "" & bh7_w75_2_c3 & bh7_w75_14_c3;
   bh7_w74_23_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3(0);
   bh7_w75_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3(1);
   bh7_w76_20_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid767: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid767_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid767_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_copy768_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid767_Out0_copy768_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid769_In0_c3 <= "" & bh7_w76_1_c3 & bh7_w76_2_c3 & bh7_w76_18_c3 & bh7_w76_17_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c0 <= "" & "0";
   bh7_w76_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3(0);
   bh7_w77_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3(1);
   bh7_w78_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid769: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid769_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid769_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_copy770_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid769_Out0_copy770_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid771_In0_c3 <= "" & bh7_w77_0_c3 & bh7_w77_1_c3 & bh7_w77_14_c3;
   bh7_w77_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_c3(0);
   bh7_w78_20_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid771: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid771_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_copy772_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid771_Out0_copy772_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid773_In0_c3 <= "" & bh7_w78_0_c3 & bh7_w78_1_c3 & bh7_w78_18_c3 & bh7_w78_17_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c0 <= "" & "0";
   bh7_w78_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3(0);
   bh7_w79_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3(1);
   bh7_w80_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid773: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid773_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid773_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_copy774_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid773_Out0_copy774_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid775_In0_c3 <= "" & bh7_w79_0_c3 & bh7_w79_1_c3 & bh7_w79_14_c3;
   bh7_w79_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_c3(0);
   bh7_w80_20_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid775: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid775_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_copy776_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid775_Out0_copy776_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid777_In0_c3 <= "" & bh7_w80_0_c3 & bh7_w80_1_c3 & bh7_w80_18_c3 & bh7_w80_17_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c0 <= "" & "0";
   bh7_w80_21_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3(0);
   bh7_w81_15_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3(1);
   bh7_w82_19_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid777: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid777_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid777_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_copy778_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid777_Out0_copy778_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid779_In0_c3 <= "" & bh7_w81_0_c3 & bh7_w81_1_c3 & bh7_w81_14_c3;
   bh7_w81_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_c3(0);
   bh7_w82_20_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid779: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid779_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_copy780_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid779_Out0_copy780_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid781_In0_c3 <= "" & bh7_w82_18_c3 & bh7_w82_0_c3 & bh7_w82_17_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid781_In1_c3 <= "" & bh7_w83_14_c3 & bh7_w83_0_c3;
   bh7_w82_21_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3(0);
   bh7_w83_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3(1);
   bh7_w84_19_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid781: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid781_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid781_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_copy782_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid781_Out0_copy782_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid783_In0_c3 <= "" & bh7_w84_17_c3 & bh7_w84_18_c3 & bh7_w84_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid783_In1_c3 <= "" & bh7_w85_15_c3 & bh7_w85_0_c3;
   bh7_w84_20_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3(0);
   bh7_w85_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3(1);
   bh7_w86_17_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid783: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid783_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid783_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_copy784_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid783_Out0_copy784_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid785_In0_c3 <= "" & bh7_w86_15_c3 & bh7_w86_16_c3 & bh7_w86_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid785_In1_c3 <= "" & bh7_w87_16_c3 & bh7_w87_0_c3;
   bh7_w86_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3(0);
   bh7_w87_17_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3(1);
   bh7_w88_17_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid785: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid785_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid785_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_copy786_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid785_Out0_copy786_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid787_In0_c3 <= "" & bh7_w88_15_c3 & bh7_w88_16_c3 & bh7_w88_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid787_In1_c3 <= "" & bh7_w89_14_c3 & bh7_w89_0_c3;
   bh7_w88_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3(0);
   bh7_w89_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3(1);
   bh7_w90_17_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid787: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid787_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid787_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_copy788_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid787_Out0_copy788_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid789_In0_c3 <= "" & bh7_w90_15_c3 & bh7_w90_16_c3 & bh7_w90_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid789_In1_c3 <= "" & bh7_w91_15_c3 & bh7_w91_0_c3;
   bh7_w90_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3(0);
   bh7_w91_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3(1);
   bh7_w92_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid789: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid789_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid789_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_copy790_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid789_Out0_copy790_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid791_In0_c3 <= "" & bh7_w92_14_c3 & bh7_w92_0_c3 & "0";
   bh7_w92_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_c3(0);
   bh7_w93_17_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid791: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid791_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_copy792_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid791_Out0_copy792_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid793_In0_c3 <= "" & bh7_w93_15_c3 & bh7_w93_16_c3 & bh7_w93_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid793_In1_c3 <= "" & bh7_w94_15_c3 & bh7_w94_0_c3;
   bh7_w93_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3(0);
   bh7_w94_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3(1);
   bh7_w95_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid793: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid793_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid793_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_copy794_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid793_Out0_copy794_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid795_In0_c3 <= "" & bh7_w95_14_c3 & bh7_w95_0_c3 & "0";
   bh7_w95_16_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_c3(0);
   bh7_w96_17_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid795: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid795_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_copy796_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid795_Out0_copy796_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid797_In0_c3 <= "" & bh7_w96_15_c3 & bh7_w96_16_c3 & bh7_w96_0_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid797_In1_c3 <= "" & bh7_w97_15_c3 & bh7_w97_0_c3;
   bh7_w96_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3(0);
   bh7_w97_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3(1);
   bh7_w98_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid797: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid797_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid797_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_copy798_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid797_Out0_copy798_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid799_In0_c3 <= "" & bh7_w98_14_c3 & bh7_w98_0_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid799_In1_c3 <= "" & bh7_w99_14_c3 & bh7_w99_15_c3;
   bh7_w98_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3(0);
   bh7_w99_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3(1);
   bh7_w100_13_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid799: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid799_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid799_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_copy800_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid799_Out0_copy800_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid801_In0_c3 <= "" & bh7_w102_9_c3 & bh7_w102_10_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid801_In1_c3 <= "" & bh7_w103_9_c3;
   bh7_w102_11_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3(0);
   bh7_w103_10_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3(1);
   bh7_w104_6_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid801: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid801_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid801_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_copy802_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid801_Out0_copy802_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid803_In0_c3 <= "" & bh7_w105_6_c3 & bh7_w105_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c0 <= "" & "0";
   bh7_w105_8_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_c3(0);
   Compressor_14_3_Freq800_uid326_uid803: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid803_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid803_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_copy804_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid803_Out0_copy804_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid805_In0_c3 <= "" & bh7_w19_3_c3 & bh7_w19_2_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid805_In1_c3 <= "" & bh7_w20_2_c3;
   bh7_w19_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3(0);
   bh7_w20_3_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3(1);
   bh7_w21_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid805: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid805_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid805_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_copy806_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid805_Out0_copy806_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid807_In0_c3 <= "" & bh7_w21_3_c3 & bh7_w21_2_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid807_In1_c3 <= "" & bh7_w22_2_c3;
   bh7_w21_5_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3(0);
   bh7_w22_3_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3(1);
   bh7_w23_4_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid807: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid807_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid807_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_copy808_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid807_Out0_copy808_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid809_In0_c3 <= "" & bh7_w23_3_c3 & bh7_w23_2_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid809_In1_c3 <= "" & bh7_w24_4_c3 & bh7_w24_3_c3;
   bh7_w23_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3(0);
   bh7_w24_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3(1);
   bh7_w25_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid809: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid809_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid809_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_copy810_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid809_Out0_copy810_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid811_In0_c3 <= "" & bh7_w25_2_c3 & bh7_w25_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid811_In1_c3 <= "" & bh7_w26_4_c3 & bh7_w26_3_c3;
   bh7_w25_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3(0);
   bh7_w26_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3(1);
   bh7_w27_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid811: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid811_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid811_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_copy812_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid811_Out0_copy812_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid813_In0_c3 <= "" & bh7_w27_2_c3 & bh7_w27_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid813_In1_c3 <= "" & bh7_w28_4_c3 & bh7_w28_3_c3;
   bh7_w27_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3(0);
   bh7_w28_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3(1);
   bh7_w29_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid813: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid813_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid813_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_copy814_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid813_Out0_copy814_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid815_In0_c3 <= "" & bh7_w29_2_c3 & bh7_w29_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid815_In1_c3 <= "" & bh7_w30_4_c3 & bh7_w30_3_c3;
   bh7_w29_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3(0);
   bh7_w30_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3(1);
   bh7_w31_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid815: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid815_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid815_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_copy816_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid815_Out0_copy816_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid817_In0_c3 <= "" & bh7_w31_2_c3 & bh7_w31_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid817_In1_c3 <= "" & bh7_w32_4_c3 & bh7_w32_3_c3;
   bh7_w31_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3(0);
   bh7_w32_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3(1);
   bh7_w33_4_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid817: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid817_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid817_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_copy818_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid817_Out0_copy818_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid819_In0_c3 <= "" & bh7_w33_2_c3 & bh7_w33_3_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid819_In1_c3 <= "" & bh7_w34_5_c3 & bh7_w34_4_c3;
   bh7_w33_5_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3(0);
   bh7_w34_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3(1);
   bh7_w35_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid819: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid819_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid819_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_copy820_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid819_Out0_copy820_c3; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid821_In0_c3 <= "" & bh7_w35_5_c3 & bh7_w35_4_c3 & "0";
   bh7_w35_7_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_c3(0);
   bh7_w36_7_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_c3(1);
   Compressor_3_2_Freq800_uid432_uid821: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid821_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_copy822_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_c3 <= Compressor_3_2_Freq800_uid432_bh7_uid821_Out0_copy822_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid823_In0_c3 <= "" & bh7_w36_6_c3 & bh7_w36_5_c3 & bh7_w36_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid823_In1_c3 <= "" & bh7_w37_5_c3 & bh7_w37_4_c3;
   bh7_w36_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3(0);
   bh7_w37_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3(1);
   bh7_w38_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid823: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid823_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid823_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_copy824_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid823_Out0_copy824_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid825_In0_c3 <= "" & bh7_w38_6_c3 & bh7_w38_5_c3 & bh7_w38_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid825_In1_c3 <= "" & bh7_w39_5_c3 & bh7_w39_4_c3;
   bh7_w38_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3(0);
   bh7_w39_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3(1);
   bh7_w40_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid825: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid825_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid825_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_copy826_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid825_Out0_copy826_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid827_In0_c3 <= "" & bh7_w40_6_c3 & bh7_w40_5_c3 & bh7_w40_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid827_In1_c3 <= "" & bh7_w41_5_c3 & bh7_w41_4_c3;
   bh7_w40_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3(0);
   bh7_w41_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3(1);
   bh7_w42_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid827: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid827_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid827_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_copy828_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid827_Out0_copy828_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid829_In0_c3 <= "" & bh7_w42_6_c3 & bh7_w42_5_c3 & bh7_w42_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid829_In1_c3 <= "" & bh7_w43_5_c3 & bh7_w43_4_c3;
   bh7_w42_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3(0);
   bh7_w43_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3(1);
   bh7_w44_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid829: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid829_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid829_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_copy830_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid829_Out0_copy830_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid831_In0_c3 <= "" & bh7_w44_6_c3 & bh7_w44_5_c3 & bh7_w44_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid831_In1_c3 <= "" & bh7_w45_5_c3 & bh7_w45_4_c3;
   bh7_w44_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3(0);
   bh7_w45_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3(1);
   bh7_w46_7_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid831: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid831_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid831_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_copy832_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid831_Out0_copy832_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid833_In0_c3 <= "" & bh7_w46_6_c3 & bh7_w46_5_c3 & bh7_w46_4_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid833_In1_c3 <= "" & bh7_w47_5_c3 & bh7_w47_4_c3;
   bh7_w46_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3(0);
   bh7_w47_6_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3(1);
   bh7_w48_8_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid833: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid833_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid833_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_copy834_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid833_Out0_copy834_c3; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid835_In0_c3 <= "" & bh7_w48_3_c3 & bh7_w48_7_c3 & bh7_w48_6_c3 & bh7_w48_5_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid835_In1_c3 <= "" & bh7_w49_7_c3;
   bh7_w48_9_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3(0);
   bh7_w49_8_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3(1);
   bh7_w50_10_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3(2);
   Compressor_14_3_Freq800_uid326_uid835: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid835_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid835_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_copy836_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_c3 <= Compressor_14_3_Freq800_uid326_bh7_uid835_Out0_copy836_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid837_In0_c3 <= "" & bh7_w50_9_c3 & bh7_w50_8_c3 & bh7_w50_7_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid837_In1_c3 <= "" & bh7_w51_13_c3 & bh7_w51_12_c3;
   bh7_w50_11_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3(0);
   bh7_w51_14_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3(1);
   bh7_w52_15_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid837: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid837_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid837_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_copy838_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid837_Out0_copy838_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid839_In0_c3 <= "" & bh7_w52_14_c3 & bh7_w52_13_c3 & bh7_w52_12_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid839_In1_c3 <= "" & bh7_w53_17_c3 & bh7_w53_16_c3;
   bh7_w52_16_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3(0);
   bh7_w53_18_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3(1);
   bh7_w54_19_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid839: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid839_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid839_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_copy840_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid839_Out0_copy840_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid841_In0_c3 <= "" & bh7_w54_18_c3 & bh7_w54_17_c3 & bh7_w54_16_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid841_In1_c3 <= "" & bh7_w55_19_c3 & bh7_w55_20_c3;
   bh7_w54_20_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3(0);
   bh7_w55_21_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3(1);
   bh7_w56_19_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3(2);
   Compressor_23_3_Freq800_uid322_uid841: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid841_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid841_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_copy842_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_c3 <= Compressor_23_3_Freq800_uid322_bh7_uid841_Out0_copy842_c3; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid843_In0_c3 <= "" & bh7_w56_16_c3 & bh7_w56_17_c3 & bh7_w56_18_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid843_In1_c3 <= "" & bh7_w57_21_c3 & bh7_w57_22_c3;
   bh7_w56_20_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4(0);
   bh7_w57_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4(1);
   bh7_w58_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid843: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid843_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid843_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid843_Out0_copy844_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid845_In0_c3 <= "" & bh7_w58_20_c3 & bh7_w58_21_c3 & bh7_w58_5_c3 & bh7_w58_22_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c0 <= "" & "0";
   bh7_w58_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4(0);
   bh7_w59_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4(1);
   bh7_w60_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid845: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid845_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid845_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid845_Out0_copy846_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid847_In0_c3 <= "" & bh7_w59_18_c3 & bh7_w59_20_c3 & bh7_w59_19_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid847_In1_c3 <= "" & bh7_w60_20_c3 & bh7_w60_21_c3;
   bh7_w59_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4(0);
   bh7_w60_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4(1);
   bh7_w61_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid847: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid847_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid847_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid847_Out0_copy848_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid849_In0_c3 <= "" & bh7_w61_20_c3 & bh7_w61_21_c3 & bh7_w61_22_c3;
   bh7_w61_24_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_c4(0);
   bh7_w62_20_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_c4(1);
   Compressor_3_2_Freq800_uid432_uid849: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid849_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid849_Out0_copy850_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid851_In0_c3 <= "" & bh7_w62_17_c3 & bh7_w62_18_c3 & bh7_w62_19_c3 & bh7_w62_4_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid851_In1_c3 <= "" & bh7_w63_20_c3;
   bh7_w62_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4(0);
   bh7_w63_23_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4(1);
   bh7_w64_23_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid851: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid851_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid851_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid851_Out0_copy852_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid853_In0_c3 <= "" & bh7_w63_21_c3 & bh7_w63_5_c3 & bh7_w63_22_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c0 <= "" & "0" & "0";
   bh7_w63_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4(0);
   bh7_w64_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4(1);
   bh7_w65_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid853: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid853_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid853_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid853_Out0_copy854_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid855_In0_c3 <= "" & bh7_w64_20_c3 & bh7_w64_22_c3 & bh7_w64_21_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid855_In1_c3 <= "" & bh7_w65_16_c3 & bh7_w65_17_c3;
   bh7_w64_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4(0);
   bh7_w65_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4(1);
   bh7_w66_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid855: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid855_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid855_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid855_Out0_copy856_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid857_In0_c3 <= "" & bh7_w66_19_c3 & bh7_w66_20_c3 & bh7_w66_21_c3;
   bh7_w66_23_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_c4(0);
   bh7_w67_20_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_c4(1);
   Compressor_3_2_Freq800_uid432_uid857: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid857_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid857_Out0_copy858_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid859_In0_c3 <= "" & bh7_w67_17_c3 & bh7_w67_19_c3 & bh7_w67_4_c3 & bh7_w67_18_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid859_In1_c3 <= "" & bh7_w68_20_c3;
   bh7_w67_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4(0);
   bh7_w68_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4(1);
   bh7_w69_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid859: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid859_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid859_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid859_Out0_copy860_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid861_In0_c3 <= "" & bh7_w69_16_c3 & bh7_w69_18_c3 & bh7_w69_17_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid861_In1_c3 <= "" & bh7_w70_20_c3 & bh7_w70_21_c3;
   bh7_w69_20_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4(0);
   bh7_w70_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4(1);
   bh7_w71_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid861: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid861_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid861_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid861_Out0_copy862_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid863_In0_c3 <= "" & bh7_w71_16_c3 & bh7_w71_17_c3 & bh7_w71_18_c3;
   bh7_w71_20_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_c4(0);
   bh7_w72_23_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_c4(1);
   Compressor_3_2_Freq800_uid432_uid863: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid863_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid863_Out0_copy864_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid865_In0_c3 <= "" & bh7_w72_20_c3 & bh7_w72_22_c3 & bh7_w72_4_c3 & bh7_w72_21_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid865_In1_c3 <= "" & bh7_w73_16_c3;
   bh7_w72_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4(0);
   bh7_w73_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4(1);
   bh7_w74_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid865: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid865_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid865_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid865_Out0_copy866_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid867_In0_c3 <= "" & bh7_w74_20_c3 & bh7_w74_22_c3 & bh7_w74_21_c3 & bh7_w74_23_c3;
   Compressor_14_3_Freq800_uid326_bh7_uid867_In1_c3 <= "" & bh7_w75_15_c3;
   bh7_w74_25_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4(0);
   bh7_w75_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4(1);
   bh7_w76_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid867: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid867_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid867_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid867_Out0_copy868_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid869_In0_c3 <= "" & bh7_w76_19_c3 & bh7_w76_21_c3 & bh7_w76_20_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid869_In1_c3 <= "" & bh7_w77_15_c3 & bh7_w77_16_c3;
   bh7_w76_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4(0);
   bh7_w77_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4(1);
   bh7_w78_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid869: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid869_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid869_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid869_Out0_copy870_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid871_In0_c3 <= "" & bh7_w78_19_c3 & bh7_w78_21_c3 & bh7_w78_20_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid871_In1_c3 <= "" & bh7_w79_15_c3 & bh7_w79_16_c3;
   bh7_w78_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4(0);
   bh7_w79_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4(1);
   bh7_w80_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid871: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid871_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid871_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid871_Out0_copy872_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid873_In0_c3 <= "" & bh7_w80_19_c3 & bh7_w80_21_c3 & bh7_w80_20_c3;
   Compressor_23_3_Freq800_uid322_bh7_uid873_In1_c3 <= "" & bh7_w81_15_c3 & bh7_w81_16_c3;
   bh7_w80_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4(0);
   bh7_w81_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4(1);
   bh7_w82_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid873: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid873_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid873_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid873_Out0_copy874_c4; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq800_uid432_bh7_uid875_In0_c3 <= "" & bh7_w82_19_c3 & bh7_w82_21_c3 & bh7_w82_20_c3;
   bh7_w82_23_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_c4(0);
   bh7_w83_16_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_c4(1);
   Compressor_3_2_Freq800_uid432_uid875: Compressor_3_2_Freq800_uid432
      port map ( X0 => Compressor_3_2_Freq800_uid432_bh7_uid875_In0_c3,
                 R => Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c3);
   Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_c4 <= Compressor_3_2_Freq800_uid432_bh7_uid875_Out0_copy876_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid877_In0_c3 <= "" & bh7_w84_19_c3 & bh7_w84_20_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid877_In1_c3 <= "" & bh7_w85_16_c3;
   bh7_w84_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4(0);
   bh7_w85_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4(1);
   bh7_w86_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid877: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid877_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid877_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid877_Out0_copy878_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid879_In0_c3 <= "" & bh7_w86_17_c3 & bh7_w86_18_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid879_In1_c3 <= "" & bh7_w87_17_c3;
   bh7_w86_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4(0);
   bh7_w87_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4(1);
   bh7_w88_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid879: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid879_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid879_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid879_Out0_copy880_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid881_In0_c3 <= "" & bh7_w88_17_c3 & bh7_w88_18_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid881_In1_c3 <= "" & bh7_w89_15_c3;
   bh7_w88_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4(0);
   bh7_w89_16_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4(1);
   bh7_w90_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid881: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid881_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid881_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid881_Out0_copy882_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid883_In0_c3 <= "" & bh7_w90_17_c3 & bh7_w90_18_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid883_In1_c3 <= "" & bh7_w91_16_c3;
   bh7_w90_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4(0);
   bh7_w91_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4(1);
   bh7_w92_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid883: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid883_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid883_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid883_Out0_copy884_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid885_In0_c3 <= "" & bh7_w92_15_c3 & bh7_w92_16_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid885_In1_c3 <= "" & bh7_w93_17_c3 & bh7_w93_18_c3;
   bh7_w92_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4(0);
   bh7_w93_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4(1);
   bh7_w94_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid885: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid885_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid885_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid885_Out0_copy886_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid887_In0_c3 <= "" & bh7_w95_15_c3 & bh7_w95_16_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid887_In1_c3 <= "" & bh7_w96_17_c3 & bh7_w96_18_c3;
   bh7_w95_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4(0);
   bh7_w96_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4(1);
   bh7_w97_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid887: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid887_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid887_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid887_Out0_copy888_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid889_In0_c3 <= "" & bh7_w98_15_c3 & bh7_w98_16_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid889_In1_c3 <= "" & bh7_w99_16_c3;
   bh7_w98_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4(0);
   bh7_w99_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4(1);
   bh7_w100_14_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid889: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid889_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid889_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid889_Out0_copy890_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid891_In0_c3 <= "" & bh7_w100_12_c3 & bh7_w100_13_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid891_In1_c3 <= "" & bh7_w101_11_c3;
   bh7_w100_15_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4(0);
   bh7_w101_12_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4(1);
   bh7_w102_12_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid891: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid891_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid891_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid891_Out0_copy892_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid893_In0_c3 <= "" & bh7_w104_5_c3 & bh7_w104_6_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid893_In1_c3 <= "" & bh7_w105_8_c3;
   bh7_w104_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_c4(0);
   bh7_w105_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_c4(1);
   Compressor_14_3_Freq800_uid326_uid893: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid893_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid893_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid893_Out0_copy894_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid895_In0_c3 <= "" & bh7_w21_5_c3 & bh7_w21_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid895_In1_c3 <= "" & bh7_w22_3_c3;
   bh7_w21_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4(0);
   bh7_w22_4_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4(1);
   bh7_w23_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid895: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid895_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid895_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid895_Out0_copy896_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid897_In0_c3 <= "" & bh7_w23_5_c3 & bh7_w23_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid897_In1_c3 <= "" & bh7_w24_5_c3;
   bh7_w23_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4(0);
   bh7_w24_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4(1);
   bh7_w25_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid897: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid897_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid897_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid897_Out0_copy898_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid899_In0_c3 <= "" & bh7_w25_5_c3 & bh7_w25_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid899_In1_c3 <= "" & bh7_w26_5_c3;
   bh7_w25_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4(0);
   bh7_w26_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4(1);
   bh7_w27_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid899: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid899_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid899_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid899_Out0_copy900_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid901_In0_c3 <= "" & bh7_w27_5_c3 & bh7_w27_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid901_In1_c3 <= "" & bh7_w28_5_c3;
   bh7_w27_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4(0);
   bh7_w28_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4(1);
   bh7_w29_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid901: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid901_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid901_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid901_Out0_copy902_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid903_In0_c3 <= "" & bh7_w29_5_c3 & bh7_w29_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid903_In1_c3 <= "" & bh7_w30_5_c3;
   bh7_w29_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4(0);
   bh7_w30_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4(1);
   bh7_w31_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid903: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid903_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid903_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid903_Out0_copy904_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid905_In0_c3 <= "" & bh7_w31_5_c3 & bh7_w31_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid905_In1_c3 <= "" & bh7_w32_5_c3;
   bh7_w31_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4(0);
   bh7_w32_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4(1);
   bh7_w33_6_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid905: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid905_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid905_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid905_Out0_copy906_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid907_In0_c3 <= "" & bh7_w33_5_c3 & bh7_w33_4_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid907_In1_c3 <= "" & bh7_w34_6_c3;
   bh7_w33_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4(0);
   bh7_w34_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4(1);
   bh7_w35_8_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid907: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid907_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid907_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid907_Out0_copy908_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid909_In0_c3 <= "" & bh7_w35_7_c3 & bh7_w35_6_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid909_In1_c3 <= "" & bh7_w36_8_c3 & bh7_w36_7_c3;
   bh7_w35_9_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4(0);
   bh7_w36_9_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4(1);
   bh7_w37_7_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid909: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid909_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid909_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid909_Out0_copy910_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid911_In0_c3 <= "" & bh7_w38_8_c3 & bh7_w38_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid911_In1_c3 <= "" & bh7_w39_6_c3;
   bh7_w38_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4(0);
   bh7_w39_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4(1);
   bh7_w40_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid911: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid911_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid911_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid911_Out0_copy912_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid913_In0_c3 <= "" & bh7_w40_8_c3 & bh7_w40_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid913_In1_c3 <= "" & bh7_w41_6_c3;
   bh7_w40_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4(0);
   bh7_w41_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4(1);
   bh7_w42_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid913: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid913_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid913_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid913_Out0_copy914_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid915_In0_c3 <= "" & bh7_w42_8_c3 & bh7_w42_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid915_In1_c3 <= "" & bh7_w43_6_c3;
   bh7_w42_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4(0);
   bh7_w43_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4(1);
   bh7_w44_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid915: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid915_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid915_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid915_Out0_copy916_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid917_In0_c3 <= "" & bh7_w44_8_c3 & bh7_w44_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid917_In1_c3 <= "" & bh7_w45_6_c3;
   bh7_w44_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4(0);
   bh7_w45_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4(1);
   bh7_w46_9_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid917: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid917_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid917_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid917_Out0_copy918_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid919_In0_c3 <= "" & bh7_w46_8_c3 & bh7_w46_7_c3 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid919_In1_c3 <= "" & bh7_w47_6_c3;
   bh7_w46_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4(0);
   bh7_w47_7_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4(1);
   bh7_w48_10_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid919: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid919_In0_c3,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid919_In1_c3,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c3);
   Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid919_Out0_copy920_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid921_In0_c3 <= "" & bh7_w48_9_c3 & bh7_w48_8_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid921_In1_c3 <= "" & bh7_w49_6_c3 & bh7_w49_8_c3;
   bh7_w48_11_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4(0);
   bh7_w49_9_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4(1);
   bh7_w50_12_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid921: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid921_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid921_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid921_Out0_copy922_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid923_In0_c3 <= "" & bh7_w50_11_c3 & bh7_w50_10_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid923_In1_c3 <= "" & bh7_w51_11_c3 & bh7_w51_14_c3;
   bh7_w50_13_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4(0);
   bh7_w51_15_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4(1);
   bh7_w52_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid923: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid923_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid923_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid923_Out0_copy924_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid925_In0_c3 <= "" & bh7_w52_16_c3 & bh7_w52_15_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid925_In1_c3 <= "" & bh7_w53_15_c3 & bh7_w53_18_c3;
   bh7_w52_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4(0);
   bh7_w53_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4(1);
   bh7_w54_21_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid925: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid925_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid925_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid925_Out0_copy926_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid927_In0_c3 <= "" & bh7_w54_20_c3 & bh7_w54_19_c3 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid927_In1_c3 <= "" & bh7_w55_21_c3 & bh7_w55_18_c3;
   bh7_w54_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4(0);
   bh7_w55_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4(1);
   bh7_w56_21_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid927: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid927_In0_c3,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid927_In1_c3,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c3);
   Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid927_Out0_copy928_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid929_In0_c4 <= "" & bh7_w56_19_c4 & bh7_w56_20_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid929_In1_c4 <= "" & bh7_w57_23_c4 & bh7_w57_24_c4;
   bh7_w56_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4(0);
   bh7_w57_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4(1);
   bh7_w58_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid929: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid929_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid929_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_copy930_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid929_Out0_copy930_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid931_In0_c4 <= "" & bh7_w58_23_c4 & bh7_w58_24_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid931_In1_c4 <= "" & bh7_w59_21_c4 & bh7_w59_22_c4;
   bh7_w58_26_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4(0);
   bh7_w59_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4(1);
   bh7_w60_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid931: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid931_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid931_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_copy932_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid931_Out0_copy932_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid933_In0_c4 <= "" & bh7_w60_22_c4 & bh7_w60_23_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid933_In1_c4 <= "" & bh7_w61_23_c4 & bh7_w61_24_c4;
   bh7_w60_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4(0);
   bh7_w61_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4(1);
   bh7_w62_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid933: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid933_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid933_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_copy934_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid933_Out0_copy934_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid935_In0_c4 <= "" & bh7_w62_20_c4 & bh7_w62_21_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid935_In1_c4 <= "" & bh7_w63_23_c4 & bh7_w63_24_c4;
   bh7_w62_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4(0);
   bh7_w63_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4(1);
   bh7_w64_26_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid935: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid935_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid935_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_copy936_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid935_Out0_copy936_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid937_In0_c4 <= "" & bh7_w64_23_c4 & bh7_w64_24_c4 & bh7_w64_25_c4;
   Compressor_23_3_Freq800_uid322_bh7_uid937_In1_c4 <= "" & bh7_w65_18_c4 & bh7_w65_19_c4;
   bh7_w64_27_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4(0);
   bh7_w65_20_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4(1);
   bh7_w66_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid937: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid937_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid937_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_copy938_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid937_Out0_copy938_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid939_In0_c4 <= "" & bh7_w66_22_c4 & bh7_w66_23_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid939_In1_c4 <= "" & bh7_w67_20_c4 & bh7_w67_21_c4;
   bh7_w66_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4(0);
   bh7_w67_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4(1);
   bh7_w68_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid939: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid939_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid939_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_copy940_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid939_Out0_copy940_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid941_In0_c4 <= "" & bh7_w68_22_c4 & bh7_w68_21_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid941_In1_c4 <= "" & bh7_w69_19_c4 & bh7_w69_20_c4;
   bh7_w68_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4(0);
   bh7_w69_21_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4(1);
   bh7_w70_23_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid941: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid941_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid941_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_copy942_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid941_Out0_copy942_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid943_In0_c4 <= "" & bh7_w71_19_c4 & bh7_w71_20_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid943_In1_c4 <= "" & bh7_w72_23_c4 & bh7_w72_24_c4;
   bh7_w71_21_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4(0);
   bh7_w72_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4(1);
   bh7_w73_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid943: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid943_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid943_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_copy944_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid943_Out0_copy944_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid945_In0_c4 <= "" & bh7_w73_18_c4 & bh7_w73_17_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid945_In1_c4 <= "" & bh7_w74_24_c4 & bh7_w74_25_c4;
   bh7_w73_20_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4(0);
   bh7_w74_26_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4(1);
   bh7_w75_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid945: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid945_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid945_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_copy946_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid945_Out0_copy946_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid947_In0_c4 <= "" & bh7_w75_17_c4 & bh7_w75_16_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid947_In1_c4 <= "" & bh7_w76_22_c4 & bh7_w76_23_c4;
   bh7_w75_19_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4(0);
   bh7_w76_24_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4(1);
   bh7_w77_18_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid947: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid947_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid947_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_copy948_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid947_Out0_copy948_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid949_In0_c4 <= "" & bh7_w78_22_c4 & bh7_w78_23_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid949_In1_c4 <= "" & bh7_w79_17_c4;
   bh7_w78_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4(0);
   bh7_w79_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4(1);
   bh7_w80_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid949: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid949_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid949_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_copy950_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid949_Out0_copy950_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid951_In0_c4 <= "" & bh7_w80_22_c4 & bh7_w80_23_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid951_In1_c4 <= "" & bh7_w81_17_c4;
   bh7_w80_25_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4(0);
   bh7_w81_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4(1);
   bh7_w82_24_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid951: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid951_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid951_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_copy952_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid951_Out0_copy952_c4; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq800_uid322_bh7_uid953_In0_c4 <= "" & bh7_w82_22_c4 & bh7_w82_23_c4 & "0";
   Compressor_23_3_Freq800_uid322_bh7_uid953_In1_c4 <= "" & bh7_w83_15_c4 & bh7_w83_16_c4;
   bh7_w82_25_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4(0);
   bh7_w83_17_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4(1);
   bh7_w84_22_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4(2);
   Compressor_23_3_Freq800_uid322_uid953: Compressor_23_3_Freq800_uid322
      port map ( X0 => Compressor_23_3_Freq800_uid322_bh7_uid953_In0_c4,
                 X1 => Compressor_23_3_Freq800_uid322_bh7_uid953_In1_c4,
                 R => Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_copy954_c4);
   Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_c4 <= Compressor_23_3_Freq800_uid322_bh7_uid953_Out0_copy954_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid955_In0_c4 <= "" & bh7_w86_19_c4 & bh7_w86_20_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid955_In1_c4 <= "" & bh7_w87_18_c4;
   bh7_w86_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4(0);
   bh7_w87_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4(1);
   bh7_w88_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid955: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid955_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid955_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_copy956_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid955_Out0_copy956_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid957_In0_c4 <= "" & bh7_w88_19_c4 & bh7_w88_20_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid957_In1_c4 <= "" & bh7_w89_16_c4;
   bh7_w88_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4(0);
   bh7_w89_17_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4(1);
   bh7_w90_21_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid957: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid957_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid957_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_copy958_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid957_Out0_copy958_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid959_In0_c4 <= "" & bh7_w90_19_c4 & bh7_w90_20_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid959_In1_c4 <= "" & bh7_w91_17_c4;
   bh7_w90_22_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4(0);
   bh7_w91_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4(1);
   bh7_w92_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid959: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid959_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid959_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_copy960_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid959_Out0_copy960_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid961_In0_c4 <= "" & bh7_w92_17_c4 & bh7_w92_18_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid961_In1_c4 <= "" & bh7_w93_19_c4;
   bh7_w92_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4(0);
   bh7_w93_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4(1);
   bh7_w94_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid961: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid961_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid961_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_copy962_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid961_Out0_copy962_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid963_In0_c4 <= "" & bh7_w94_16_c4 & bh7_w94_17_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid963_In1_c4 <= "" & bh7_w95_17_c4;
   bh7_w94_19_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4(0);
   bh7_w95_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4(1);
   bh7_w96_20_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid963: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid963_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid963_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_copy964_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid963_Out0_copy964_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid965_In0_c4 <= "" & bh7_w97_16_c4 & bh7_w97_17_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid965_In1_c4 <= "" & bh7_w98_17_c4;
   bh7_w97_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4(0);
   bh7_w98_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4(1);
   bh7_w99_18_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid965: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid965_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid965_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_copy966_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid965_Out0_copy966_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid967_In0_c4 <= "" & bh7_w100_14_c4 & bh7_w100_15_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid967_In1_c4 <= "" & bh7_w101_12_c4;
   bh7_w100_16_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4(0);
   bh7_w101_13_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4(1);
   bh7_w102_13_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid967: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid967_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid967_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_copy968_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid967_Out0_copy968_c4; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq800_uid326_bh7_uid969_In0_c4 <= "" & bh7_w102_11_c4 & bh7_w102_12_c4 & "0" & "0";
   Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c3 <= "" & bh7_w103_10_c3;
   bh7_w102_14_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4(0);
   bh7_w103_11_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4(1);
   bh7_w104_8_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4(2);
   Compressor_14_3_Freq800_uid326_uid969: Compressor_14_3_Freq800_uid326
      port map ( X0 => Compressor_14_3_Freq800_uid326_bh7_uid969_In0_c4,
                 X1 => Compressor_14_3_Freq800_uid326_bh7_uid969_In1_c4,
                 R => Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_copy970_c4);
   Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_c4 <= Compressor_14_3_Freq800_uid326_bh7_uid969_Out0_copy970_c4; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh7_22_c4 <= bh7_w22_4_c4 & bh7_w21_6_c4 & bh7_w20_3_c4 & bh7_w19_4_c4 & bh7_w18_2_c4 & bh7_w17_2_c4 & bh7_w16_0_c4 & bh7_w15_0_c4 & bh7_w14_0_c4 & bh7_w13_0_c4 & bh7_w12_0_c4 & bh7_w11_0_c4 & bh7_w10_0_c4 & bh7_w9_0_c4 & bh7_w8_0_c4 & bh7_w7_0_c4 & bh7_w6_0_c4 & bh7_w5_0_c4 & bh7_w4_0_c4 & bh7_w3_0_c4 & bh7_w2_0_c4 & bh7_w1_0_c4 & bh7_w0_0_c4;

   bitheapFinalAdd_bh7_In0_c4 <= "0" & bh7_w105_9_c4 & bh7_w104_7_c4 & bh7_w103_11_c4 & bh7_w102_13_c4 & bh7_w101_13_c4 & bh7_w100_16_c4 & bh7_w99_17_c4 & bh7_w98_18_c4 & bh7_w97_18_c4 & bh7_w96_19_c4 & bh7_w95_18_c4 & bh7_w94_18_c4 & bh7_w93_20_c4 & bh7_w92_19_c4 & bh7_w91_18_c4 & bh7_w90_21_c4 & bh7_w89_17_c4 & bh7_w88_21_c4 & bh7_w87_19_c4 & bh7_w86_21_c4 & bh7_w85_17_c4 & bh7_w84_21_c4 & bh7_w83_17_c4 & bh7_w82_24_c4 & bh7_w81_18_c4 & bh7_w80_24_c4 & bh7_w79_18_c4 & bh7_w78_24_c4 & bh7_w77_17_c4 & bh7_w76_24_c4 & bh7_w75_18_c4 & bh7_w74_26_c4 & bh7_w73_19_c4 & bh7_w72_25_c4 & bh7_w71_21_c4 & bh7_w70_22_c4 & bh7_w69_21_c4 & bh7_w68_23_c4 & bh7_w67_22_c4 & bh7_w66_24_c4 & bh7_w65_20_c4 & bh7_w64_26_c4 & bh7_w63_25_c4 & bh7_w62_22_c4 & bh7_w61_25_c4 & bh7_w60_24_c4 & bh7_w59_23_c4 & bh7_w58_25_c4 & bh7_w57_25_c4 & bh7_w56_21_c4 & bh7_w55_22_c4 & bh7_w54_22_c4 & bh7_w53_19_c4 & bh7_w52_18_c4 & bh7_w51_15_c4 & bh7_w50_13_c4 & bh7_w49_9_c4 & bh7_w48_11_c4 & bh7_w47_7_c4 & bh7_w46_10_c4 & bh7_w45_7_c4 & bh7_w44_10_c4 & bh7_w43_7_c4 & bh7_w42_10_c4 & bh7_w41_7_c4 & bh7_w40_10_c4 & bh7_w39_7_c4 & bh7_w38_9_c4 & bh7_w37_6_c4 & bh7_w36_9_c4 & bh7_w35_9_c4 & bh7_w34_7_c4 & bh7_w33_7_c4 & bh7_w32_6_c4 & bh7_w31_7_c4 & bh7_w30_6_c4 & bh7_w29_7_c4 & bh7_w28_6_c4 & bh7_w27_7_c4 & bh7_w26_6_c4 & bh7_w25_7_c4 & bh7_w24_6_c4 & bh7_w23_7_c4;
   bitheapFinalAdd_bh7_In1_c4 <= "0" & "0" & bh7_w104_8_c4 & "0" & bh7_w102_14_c4 & "0" & "0" & bh7_w99_18_c4 & "0" & "0" & bh7_w96_20_c4 & "0" & bh7_w94_19_c4 & "0" & bh7_w92_20_c4 & "0" & bh7_w90_22_c4 & "0" & bh7_w88_22_c4 & "0" & "0" & "0" & bh7_w84_22_c4 & "0" & bh7_w82_25_c4 & "0" & bh7_w80_25_c4 & "0" & "0" & bh7_w77_18_c4 & "0" & bh7_w75_19_c4 & "0" & bh7_w73_20_c4 & "0" & "0" & bh7_w70_23_c4 & "0" & bh7_w68_24_c4 & "0" & bh7_w66_25_c4 & "0" & bh7_w64_27_c4 & "0" & bh7_w62_23_c4 & "0" & bh7_w60_25_c4 & "0" & bh7_w58_26_c4 & "0" & bh7_w56_22_c4 & "0" & bh7_w54_21_c4 & "0" & bh7_w52_17_c4 & "0" & bh7_w50_12_c4 & "0" & bh7_w48_10_c4 & "0" & bh7_w46_9_c4 & "0" & bh7_w44_9_c4 & "0" & bh7_w42_9_c4 & "0" & bh7_w40_9_c4 & "0" & "0" & bh7_w37_7_c4 & "0" & bh7_w35_8_c4 & "0" & bh7_w33_6_c4 & "0" & bh7_w31_6_c4 & "0" & bh7_w29_6_c4 & "0" & bh7_w27_6_c4 & "0" & bh7_w25_6_c4 & "0" & bh7_w23_6_c4;
   bitheapFinalAdd_bh7_Cin_c0 <= '0';

   bitheapFinalAdd_bh7: IntAdder_84_Freq800_uid972
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 Cin => bitheapFinalAdd_bh7_Cin_c0,
                 X => bitheapFinalAdd_bh7_In0_c4,
                 Y => bitheapFinalAdd_bh7_In1_c4,
                 R => bitheapFinalAdd_bh7_Out_c33);
   bitheapResult_bh7_c33 <= bitheapFinalAdd_bh7_Out_c33(82 downto 0) & tmp_bitheapResult_bh7_22_c33;
   R <= bitheapResult_bh7_c33(105 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_65_Freq800_uid975
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 56 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_65_Freq800_uid975 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56 : in std_logic;
          X : in  std_logic_vector(64 downto 0);
          Y : in  std_logic_vector(64 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(64 downto 0)   );
end entity;

architecture arch of IntAdder_65_Freq800_uid975 is
signal Cin_1_c34, Cin_1_c35 :  std_logic;
signal X_1_c33, X_1_c34, X_1_c35 :  std_logic_vector(3 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3, Y_1_c4, Y_1_c5, Y_1_c6, Y_1_c7, Y_1_c8, Y_1_c9, Y_1_c10, Y_1_c11, Y_1_c12, Y_1_c13, Y_1_c14, Y_1_c15, Y_1_c16, Y_1_c17, Y_1_c18, Y_1_c19, Y_1_c20, Y_1_c21, Y_1_c22, Y_1_c23, Y_1_c24, Y_1_c25, Y_1_c26, Y_1_c27, Y_1_c28, Y_1_c29, Y_1_c30, Y_1_c31, Y_1_c32, Y_1_c33, Y_1_c34, Y_1_c35 :  std_logic_vector(3 downto 0);
signal S_1_c35 :  std_logic_vector(3 downto 0);
signal R_1_c35, R_1_c36, R_1_c37, R_1_c38, R_1_c39, R_1_c40, R_1_c41, R_1_c42, R_1_c43, R_1_c44, R_1_c45, R_1_c46, R_1_c47, R_1_c48, R_1_c49, R_1_c50, R_1_c51, R_1_c52, R_1_c53, R_1_c54, R_1_c55, R_1_c56 :  std_logic_vector(2 downto 0);
signal Cin_2_c35, Cin_2_c36 :  std_logic;
signal X_2_c33, X_2_c34, X_2_c35, X_2_c36 :  std_logic_vector(3 downto 0);
signal Y_2_c0, Y_2_c1, Y_2_c2, Y_2_c3, Y_2_c4, Y_2_c5, Y_2_c6, Y_2_c7, Y_2_c8, Y_2_c9, Y_2_c10, Y_2_c11, Y_2_c12, Y_2_c13, Y_2_c14, Y_2_c15, Y_2_c16, Y_2_c17, Y_2_c18, Y_2_c19, Y_2_c20, Y_2_c21, Y_2_c22, Y_2_c23, Y_2_c24, Y_2_c25, Y_2_c26, Y_2_c27, Y_2_c28, Y_2_c29, Y_2_c30, Y_2_c31, Y_2_c32, Y_2_c33, Y_2_c34, Y_2_c35, Y_2_c36 :  std_logic_vector(3 downto 0);
signal S_2_c36 :  std_logic_vector(3 downto 0);
signal R_2_c36, R_2_c37, R_2_c38, R_2_c39, R_2_c40, R_2_c41, R_2_c42, R_2_c43, R_2_c44, R_2_c45, R_2_c46, R_2_c47, R_2_c48, R_2_c49, R_2_c50, R_2_c51, R_2_c52, R_2_c53, R_2_c54, R_2_c55, R_2_c56 :  std_logic_vector(2 downto 0);
signal Cin_3_c36, Cin_3_c37 :  std_logic;
signal X_3_c33, X_3_c34, X_3_c35, X_3_c36, X_3_c37 :  std_logic_vector(3 downto 0);
signal Y_3_c0, Y_3_c1, Y_3_c2, Y_3_c3, Y_3_c4, Y_3_c5, Y_3_c6, Y_3_c7, Y_3_c8, Y_3_c9, Y_3_c10, Y_3_c11, Y_3_c12, Y_3_c13, Y_3_c14, Y_3_c15, Y_3_c16, Y_3_c17, Y_3_c18, Y_3_c19, Y_3_c20, Y_3_c21, Y_3_c22, Y_3_c23, Y_3_c24, Y_3_c25, Y_3_c26, Y_3_c27, Y_3_c28, Y_3_c29, Y_3_c30, Y_3_c31, Y_3_c32, Y_3_c33, Y_3_c34, Y_3_c35, Y_3_c36, Y_3_c37 :  std_logic_vector(3 downto 0);
signal S_3_c37 :  std_logic_vector(3 downto 0);
signal R_3_c37, R_3_c38, R_3_c39, R_3_c40, R_3_c41, R_3_c42, R_3_c43, R_3_c44, R_3_c45, R_3_c46, R_3_c47, R_3_c48, R_3_c49, R_3_c50, R_3_c51, R_3_c52, R_3_c53, R_3_c54, R_3_c55, R_3_c56 :  std_logic_vector(2 downto 0);
signal Cin_4_c37, Cin_4_c38 :  std_logic;
signal X_4_c33, X_4_c34, X_4_c35, X_4_c36, X_4_c37, X_4_c38 :  std_logic_vector(3 downto 0);
signal Y_4_c0, Y_4_c1, Y_4_c2, Y_4_c3, Y_4_c4, Y_4_c5, Y_4_c6, Y_4_c7, Y_4_c8, Y_4_c9, Y_4_c10, Y_4_c11, Y_4_c12, Y_4_c13, Y_4_c14, Y_4_c15, Y_4_c16, Y_4_c17, Y_4_c18, Y_4_c19, Y_4_c20, Y_4_c21, Y_4_c22, Y_4_c23, Y_4_c24, Y_4_c25, Y_4_c26, Y_4_c27, Y_4_c28, Y_4_c29, Y_4_c30, Y_4_c31, Y_4_c32, Y_4_c33, Y_4_c34, Y_4_c35, Y_4_c36, Y_4_c37, Y_4_c38 :  std_logic_vector(3 downto 0);
signal S_4_c38 :  std_logic_vector(3 downto 0);
signal R_4_c38, R_4_c39, R_4_c40, R_4_c41, R_4_c42, R_4_c43, R_4_c44, R_4_c45, R_4_c46, R_4_c47, R_4_c48, R_4_c49, R_4_c50, R_4_c51, R_4_c52, R_4_c53, R_4_c54, R_4_c55, R_4_c56 :  std_logic_vector(2 downto 0);
signal Cin_5_c38, Cin_5_c39 :  std_logic;
signal X_5_c33, X_5_c34, X_5_c35, X_5_c36, X_5_c37, X_5_c38, X_5_c39 :  std_logic_vector(3 downto 0);
signal Y_5_c0, Y_5_c1, Y_5_c2, Y_5_c3, Y_5_c4, Y_5_c5, Y_5_c6, Y_5_c7, Y_5_c8, Y_5_c9, Y_5_c10, Y_5_c11, Y_5_c12, Y_5_c13, Y_5_c14, Y_5_c15, Y_5_c16, Y_5_c17, Y_5_c18, Y_5_c19, Y_5_c20, Y_5_c21, Y_5_c22, Y_5_c23, Y_5_c24, Y_5_c25, Y_5_c26, Y_5_c27, Y_5_c28, Y_5_c29, Y_5_c30, Y_5_c31, Y_5_c32, Y_5_c33, Y_5_c34, Y_5_c35, Y_5_c36, Y_5_c37, Y_5_c38, Y_5_c39 :  std_logic_vector(3 downto 0);
signal S_5_c39 :  std_logic_vector(3 downto 0);
signal R_5_c39, R_5_c40, R_5_c41, R_5_c42, R_5_c43, R_5_c44, R_5_c45, R_5_c46, R_5_c47, R_5_c48, R_5_c49, R_5_c50, R_5_c51, R_5_c52, R_5_c53, R_5_c54, R_5_c55, R_5_c56 :  std_logic_vector(2 downto 0);
signal Cin_6_c39, Cin_6_c40 :  std_logic;
signal X_6_c33, X_6_c34, X_6_c35, X_6_c36, X_6_c37, X_6_c38, X_6_c39, X_6_c40 :  std_logic_vector(3 downto 0);
signal Y_6_c0, Y_6_c1, Y_6_c2, Y_6_c3, Y_6_c4, Y_6_c5, Y_6_c6, Y_6_c7, Y_6_c8, Y_6_c9, Y_6_c10, Y_6_c11, Y_6_c12, Y_6_c13, Y_6_c14, Y_6_c15, Y_6_c16, Y_6_c17, Y_6_c18, Y_6_c19, Y_6_c20, Y_6_c21, Y_6_c22, Y_6_c23, Y_6_c24, Y_6_c25, Y_6_c26, Y_6_c27, Y_6_c28, Y_6_c29, Y_6_c30, Y_6_c31, Y_6_c32, Y_6_c33, Y_6_c34, Y_6_c35, Y_6_c36, Y_6_c37, Y_6_c38, Y_6_c39, Y_6_c40 :  std_logic_vector(3 downto 0);
signal S_6_c40 :  std_logic_vector(3 downto 0);
signal R_6_c40, R_6_c41, R_6_c42, R_6_c43, R_6_c44, R_6_c45, R_6_c46, R_6_c47, R_6_c48, R_6_c49, R_6_c50, R_6_c51, R_6_c52, R_6_c53, R_6_c54, R_6_c55, R_6_c56 :  std_logic_vector(2 downto 0);
signal Cin_7_c40, Cin_7_c41 :  std_logic;
signal X_7_c33, X_7_c34, X_7_c35, X_7_c36, X_7_c37, X_7_c38, X_7_c39, X_7_c40, X_7_c41 :  std_logic_vector(3 downto 0);
signal Y_7_c0, Y_7_c1, Y_7_c2, Y_7_c3, Y_7_c4, Y_7_c5, Y_7_c6, Y_7_c7, Y_7_c8, Y_7_c9, Y_7_c10, Y_7_c11, Y_7_c12, Y_7_c13, Y_7_c14, Y_7_c15, Y_7_c16, Y_7_c17, Y_7_c18, Y_7_c19, Y_7_c20, Y_7_c21, Y_7_c22, Y_7_c23, Y_7_c24, Y_7_c25, Y_7_c26, Y_7_c27, Y_7_c28, Y_7_c29, Y_7_c30, Y_7_c31, Y_7_c32, Y_7_c33, Y_7_c34, Y_7_c35, Y_7_c36, Y_7_c37, Y_7_c38, Y_7_c39, Y_7_c40, Y_7_c41 :  std_logic_vector(3 downto 0);
signal S_7_c41 :  std_logic_vector(3 downto 0);
signal R_7_c41, R_7_c42, R_7_c43, R_7_c44, R_7_c45, R_7_c46, R_7_c47, R_7_c48, R_7_c49, R_7_c50, R_7_c51, R_7_c52, R_7_c53, R_7_c54, R_7_c55, R_7_c56 :  std_logic_vector(2 downto 0);
signal Cin_8_c41, Cin_8_c42 :  std_logic;
signal X_8_c33, X_8_c34, X_8_c35, X_8_c36, X_8_c37, X_8_c38, X_8_c39, X_8_c40, X_8_c41, X_8_c42 :  std_logic_vector(3 downto 0);
signal Y_8_c0, Y_8_c1, Y_8_c2, Y_8_c3, Y_8_c4, Y_8_c5, Y_8_c6, Y_8_c7, Y_8_c8, Y_8_c9, Y_8_c10, Y_8_c11, Y_8_c12, Y_8_c13, Y_8_c14, Y_8_c15, Y_8_c16, Y_8_c17, Y_8_c18, Y_8_c19, Y_8_c20, Y_8_c21, Y_8_c22, Y_8_c23, Y_8_c24, Y_8_c25, Y_8_c26, Y_8_c27, Y_8_c28, Y_8_c29, Y_8_c30, Y_8_c31, Y_8_c32, Y_8_c33, Y_8_c34, Y_8_c35, Y_8_c36, Y_8_c37, Y_8_c38, Y_8_c39, Y_8_c40, Y_8_c41, Y_8_c42 :  std_logic_vector(3 downto 0);
signal S_8_c42 :  std_logic_vector(3 downto 0);
signal R_8_c42, R_8_c43, R_8_c44, R_8_c45, R_8_c46, R_8_c47, R_8_c48, R_8_c49, R_8_c50, R_8_c51, R_8_c52, R_8_c53, R_8_c54, R_8_c55, R_8_c56 :  std_logic_vector(2 downto 0);
signal Cin_9_c42, Cin_9_c43 :  std_logic;
signal X_9_c33, X_9_c34, X_9_c35, X_9_c36, X_9_c37, X_9_c38, X_9_c39, X_9_c40, X_9_c41, X_9_c42, X_9_c43 :  std_logic_vector(3 downto 0);
signal Y_9_c0, Y_9_c1, Y_9_c2, Y_9_c3, Y_9_c4, Y_9_c5, Y_9_c6, Y_9_c7, Y_9_c8, Y_9_c9, Y_9_c10, Y_9_c11, Y_9_c12, Y_9_c13, Y_9_c14, Y_9_c15, Y_9_c16, Y_9_c17, Y_9_c18, Y_9_c19, Y_9_c20, Y_9_c21, Y_9_c22, Y_9_c23, Y_9_c24, Y_9_c25, Y_9_c26, Y_9_c27, Y_9_c28, Y_9_c29, Y_9_c30, Y_9_c31, Y_9_c32, Y_9_c33, Y_9_c34, Y_9_c35, Y_9_c36, Y_9_c37, Y_9_c38, Y_9_c39, Y_9_c40, Y_9_c41, Y_9_c42, Y_9_c43 :  std_logic_vector(3 downto 0);
signal S_9_c43 :  std_logic_vector(3 downto 0);
signal R_9_c43, R_9_c44, R_9_c45, R_9_c46, R_9_c47, R_9_c48, R_9_c49, R_9_c50, R_9_c51, R_9_c52, R_9_c53, R_9_c54, R_9_c55, R_9_c56 :  std_logic_vector(2 downto 0);
signal Cin_10_c43, Cin_10_c44 :  std_logic;
signal X_10_c33, X_10_c34, X_10_c35, X_10_c36, X_10_c37, X_10_c38, X_10_c39, X_10_c40, X_10_c41, X_10_c42, X_10_c43, X_10_c44 :  std_logic_vector(3 downto 0);
signal Y_10_c0, Y_10_c1, Y_10_c2, Y_10_c3, Y_10_c4, Y_10_c5, Y_10_c6, Y_10_c7, Y_10_c8, Y_10_c9, Y_10_c10, Y_10_c11, Y_10_c12, Y_10_c13, Y_10_c14, Y_10_c15, Y_10_c16, Y_10_c17, Y_10_c18, Y_10_c19, Y_10_c20, Y_10_c21, Y_10_c22, Y_10_c23, Y_10_c24, Y_10_c25, Y_10_c26, Y_10_c27, Y_10_c28, Y_10_c29, Y_10_c30, Y_10_c31, Y_10_c32, Y_10_c33, Y_10_c34, Y_10_c35, Y_10_c36, Y_10_c37, Y_10_c38, Y_10_c39, Y_10_c40, Y_10_c41, Y_10_c42, Y_10_c43, Y_10_c44 :  std_logic_vector(3 downto 0);
signal S_10_c44 :  std_logic_vector(3 downto 0);
signal R_10_c44, R_10_c45, R_10_c46, R_10_c47, R_10_c48, R_10_c49, R_10_c50, R_10_c51, R_10_c52, R_10_c53, R_10_c54, R_10_c55, R_10_c56 :  std_logic_vector(2 downto 0);
signal Cin_11_c44, Cin_11_c45 :  std_logic;
signal X_11_c33, X_11_c34, X_11_c35, X_11_c36, X_11_c37, X_11_c38, X_11_c39, X_11_c40, X_11_c41, X_11_c42, X_11_c43, X_11_c44, X_11_c45 :  std_logic_vector(3 downto 0);
signal Y_11_c0, Y_11_c1, Y_11_c2, Y_11_c3, Y_11_c4, Y_11_c5, Y_11_c6, Y_11_c7, Y_11_c8, Y_11_c9, Y_11_c10, Y_11_c11, Y_11_c12, Y_11_c13, Y_11_c14, Y_11_c15, Y_11_c16, Y_11_c17, Y_11_c18, Y_11_c19, Y_11_c20, Y_11_c21, Y_11_c22, Y_11_c23, Y_11_c24, Y_11_c25, Y_11_c26, Y_11_c27, Y_11_c28, Y_11_c29, Y_11_c30, Y_11_c31, Y_11_c32, Y_11_c33, Y_11_c34, Y_11_c35, Y_11_c36, Y_11_c37, Y_11_c38, Y_11_c39, Y_11_c40, Y_11_c41, Y_11_c42, Y_11_c43, Y_11_c44, Y_11_c45 :  std_logic_vector(3 downto 0);
signal S_11_c45 :  std_logic_vector(3 downto 0);
signal R_11_c45, R_11_c46, R_11_c47, R_11_c48, R_11_c49, R_11_c50, R_11_c51, R_11_c52, R_11_c53, R_11_c54, R_11_c55, R_11_c56 :  std_logic_vector(2 downto 0);
signal Cin_12_c45, Cin_12_c46 :  std_logic;
signal X_12_c33, X_12_c34, X_12_c35, X_12_c36, X_12_c37, X_12_c38, X_12_c39, X_12_c40, X_12_c41, X_12_c42, X_12_c43, X_12_c44, X_12_c45, X_12_c46 :  std_logic_vector(3 downto 0);
signal Y_12_c0, Y_12_c1, Y_12_c2, Y_12_c3, Y_12_c4, Y_12_c5, Y_12_c6, Y_12_c7, Y_12_c8, Y_12_c9, Y_12_c10, Y_12_c11, Y_12_c12, Y_12_c13, Y_12_c14, Y_12_c15, Y_12_c16, Y_12_c17, Y_12_c18, Y_12_c19, Y_12_c20, Y_12_c21, Y_12_c22, Y_12_c23, Y_12_c24, Y_12_c25, Y_12_c26, Y_12_c27, Y_12_c28, Y_12_c29, Y_12_c30, Y_12_c31, Y_12_c32, Y_12_c33, Y_12_c34, Y_12_c35, Y_12_c36, Y_12_c37, Y_12_c38, Y_12_c39, Y_12_c40, Y_12_c41, Y_12_c42, Y_12_c43, Y_12_c44, Y_12_c45, Y_12_c46 :  std_logic_vector(3 downto 0);
signal S_12_c46 :  std_logic_vector(3 downto 0);
signal R_12_c46, R_12_c47, R_12_c48, R_12_c49, R_12_c50, R_12_c51, R_12_c52, R_12_c53, R_12_c54, R_12_c55, R_12_c56 :  std_logic_vector(2 downto 0);
signal Cin_13_c46, Cin_13_c47 :  std_logic;
signal X_13_c33, X_13_c34, X_13_c35, X_13_c36, X_13_c37, X_13_c38, X_13_c39, X_13_c40, X_13_c41, X_13_c42, X_13_c43, X_13_c44, X_13_c45, X_13_c46, X_13_c47 :  std_logic_vector(3 downto 0);
signal Y_13_c0, Y_13_c1, Y_13_c2, Y_13_c3, Y_13_c4, Y_13_c5, Y_13_c6, Y_13_c7, Y_13_c8, Y_13_c9, Y_13_c10, Y_13_c11, Y_13_c12, Y_13_c13, Y_13_c14, Y_13_c15, Y_13_c16, Y_13_c17, Y_13_c18, Y_13_c19, Y_13_c20, Y_13_c21, Y_13_c22, Y_13_c23, Y_13_c24, Y_13_c25, Y_13_c26, Y_13_c27, Y_13_c28, Y_13_c29, Y_13_c30, Y_13_c31, Y_13_c32, Y_13_c33, Y_13_c34, Y_13_c35, Y_13_c36, Y_13_c37, Y_13_c38, Y_13_c39, Y_13_c40, Y_13_c41, Y_13_c42, Y_13_c43, Y_13_c44, Y_13_c45, Y_13_c46, Y_13_c47 :  std_logic_vector(3 downto 0);
signal S_13_c47 :  std_logic_vector(3 downto 0);
signal R_13_c47, R_13_c48, R_13_c49, R_13_c50, R_13_c51, R_13_c52, R_13_c53, R_13_c54, R_13_c55, R_13_c56 :  std_logic_vector(2 downto 0);
signal Cin_14_c47, Cin_14_c48 :  std_logic;
signal X_14_c33, X_14_c34, X_14_c35, X_14_c36, X_14_c37, X_14_c38, X_14_c39, X_14_c40, X_14_c41, X_14_c42, X_14_c43, X_14_c44, X_14_c45, X_14_c46, X_14_c47, X_14_c48 :  std_logic_vector(3 downto 0);
signal Y_14_c0, Y_14_c1, Y_14_c2, Y_14_c3, Y_14_c4, Y_14_c5, Y_14_c6, Y_14_c7, Y_14_c8, Y_14_c9, Y_14_c10, Y_14_c11, Y_14_c12, Y_14_c13, Y_14_c14, Y_14_c15, Y_14_c16, Y_14_c17, Y_14_c18, Y_14_c19, Y_14_c20, Y_14_c21, Y_14_c22, Y_14_c23, Y_14_c24, Y_14_c25, Y_14_c26, Y_14_c27, Y_14_c28, Y_14_c29, Y_14_c30, Y_14_c31, Y_14_c32, Y_14_c33, Y_14_c34, Y_14_c35, Y_14_c36, Y_14_c37, Y_14_c38, Y_14_c39, Y_14_c40, Y_14_c41, Y_14_c42, Y_14_c43, Y_14_c44, Y_14_c45, Y_14_c46, Y_14_c47, Y_14_c48 :  std_logic_vector(3 downto 0);
signal S_14_c48 :  std_logic_vector(3 downto 0);
signal R_14_c48, R_14_c49, R_14_c50, R_14_c51, R_14_c52, R_14_c53, R_14_c54, R_14_c55, R_14_c56 :  std_logic_vector(2 downto 0);
signal Cin_15_c48, Cin_15_c49 :  std_logic;
signal X_15_c33, X_15_c34, X_15_c35, X_15_c36, X_15_c37, X_15_c38, X_15_c39, X_15_c40, X_15_c41, X_15_c42, X_15_c43, X_15_c44, X_15_c45, X_15_c46, X_15_c47, X_15_c48, X_15_c49 :  std_logic_vector(3 downto 0);
signal Y_15_c0, Y_15_c1, Y_15_c2, Y_15_c3, Y_15_c4, Y_15_c5, Y_15_c6, Y_15_c7, Y_15_c8, Y_15_c9, Y_15_c10, Y_15_c11, Y_15_c12, Y_15_c13, Y_15_c14, Y_15_c15, Y_15_c16, Y_15_c17, Y_15_c18, Y_15_c19, Y_15_c20, Y_15_c21, Y_15_c22, Y_15_c23, Y_15_c24, Y_15_c25, Y_15_c26, Y_15_c27, Y_15_c28, Y_15_c29, Y_15_c30, Y_15_c31, Y_15_c32, Y_15_c33, Y_15_c34, Y_15_c35, Y_15_c36, Y_15_c37, Y_15_c38, Y_15_c39, Y_15_c40, Y_15_c41, Y_15_c42, Y_15_c43, Y_15_c44, Y_15_c45, Y_15_c46, Y_15_c47, Y_15_c48, Y_15_c49 :  std_logic_vector(3 downto 0);
signal S_15_c49 :  std_logic_vector(3 downto 0);
signal R_15_c49, R_15_c50, R_15_c51, R_15_c52, R_15_c53, R_15_c54, R_15_c55, R_15_c56 :  std_logic_vector(2 downto 0);
signal Cin_16_c49, Cin_16_c50 :  std_logic;
signal X_16_c33, X_16_c34, X_16_c35, X_16_c36, X_16_c37, X_16_c38, X_16_c39, X_16_c40, X_16_c41, X_16_c42, X_16_c43, X_16_c44, X_16_c45, X_16_c46, X_16_c47, X_16_c48, X_16_c49, X_16_c50 :  std_logic_vector(3 downto 0);
signal Y_16_c0, Y_16_c1, Y_16_c2, Y_16_c3, Y_16_c4, Y_16_c5, Y_16_c6, Y_16_c7, Y_16_c8, Y_16_c9, Y_16_c10, Y_16_c11, Y_16_c12, Y_16_c13, Y_16_c14, Y_16_c15, Y_16_c16, Y_16_c17, Y_16_c18, Y_16_c19, Y_16_c20, Y_16_c21, Y_16_c22, Y_16_c23, Y_16_c24, Y_16_c25, Y_16_c26, Y_16_c27, Y_16_c28, Y_16_c29, Y_16_c30, Y_16_c31, Y_16_c32, Y_16_c33, Y_16_c34, Y_16_c35, Y_16_c36, Y_16_c37, Y_16_c38, Y_16_c39, Y_16_c40, Y_16_c41, Y_16_c42, Y_16_c43, Y_16_c44, Y_16_c45, Y_16_c46, Y_16_c47, Y_16_c48, Y_16_c49, Y_16_c50 :  std_logic_vector(3 downto 0);
signal S_16_c50 :  std_logic_vector(3 downto 0);
signal R_16_c50, R_16_c51, R_16_c52, R_16_c53, R_16_c54, R_16_c55, R_16_c56 :  std_logic_vector(2 downto 0);
signal Cin_17_c50, Cin_17_c51 :  std_logic;
signal X_17_c33, X_17_c34, X_17_c35, X_17_c36, X_17_c37, X_17_c38, X_17_c39, X_17_c40, X_17_c41, X_17_c42, X_17_c43, X_17_c44, X_17_c45, X_17_c46, X_17_c47, X_17_c48, X_17_c49, X_17_c50, X_17_c51 :  std_logic_vector(3 downto 0);
signal Y_17_c0, Y_17_c1, Y_17_c2, Y_17_c3, Y_17_c4, Y_17_c5, Y_17_c6, Y_17_c7, Y_17_c8, Y_17_c9, Y_17_c10, Y_17_c11, Y_17_c12, Y_17_c13, Y_17_c14, Y_17_c15, Y_17_c16, Y_17_c17, Y_17_c18, Y_17_c19, Y_17_c20, Y_17_c21, Y_17_c22, Y_17_c23, Y_17_c24, Y_17_c25, Y_17_c26, Y_17_c27, Y_17_c28, Y_17_c29, Y_17_c30, Y_17_c31, Y_17_c32, Y_17_c33, Y_17_c34, Y_17_c35, Y_17_c36, Y_17_c37, Y_17_c38, Y_17_c39, Y_17_c40, Y_17_c41, Y_17_c42, Y_17_c43, Y_17_c44, Y_17_c45, Y_17_c46, Y_17_c47, Y_17_c48, Y_17_c49, Y_17_c50, Y_17_c51 :  std_logic_vector(3 downto 0);
signal S_17_c51 :  std_logic_vector(3 downto 0);
signal R_17_c51, R_17_c52, R_17_c53, R_17_c54, R_17_c55, R_17_c56 :  std_logic_vector(2 downto 0);
signal Cin_18_c51, Cin_18_c52 :  std_logic;
signal X_18_c33, X_18_c34, X_18_c35, X_18_c36, X_18_c37, X_18_c38, X_18_c39, X_18_c40, X_18_c41, X_18_c42, X_18_c43, X_18_c44, X_18_c45, X_18_c46, X_18_c47, X_18_c48, X_18_c49, X_18_c50, X_18_c51, X_18_c52 :  std_logic_vector(3 downto 0);
signal Y_18_c0, Y_18_c1, Y_18_c2, Y_18_c3, Y_18_c4, Y_18_c5, Y_18_c6, Y_18_c7, Y_18_c8, Y_18_c9, Y_18_c10, Y_18_c11, Y_18_c12, Y_18_c13, Y_18_c14, Y_18_c15, Y_18_c16, Y_18_c17, Y_18_c18, Y_18_c19, Y_18_c20, Y_18_c21, Y_18_c22, Y_18_c23, Y_18_c24, Y_18_c25, Y_18_c26, Y_18_c27, Y_18_c28, Y_18_c29, Y_18_c30, Y_18_c31, Y_18_c32, Y_18_c33, Y_18_c34, Y_18_c35, Y_18_c36, Y_18_c37, Y_18_c38, Y_18_c39, Y_18_c40, Y_18_c41, Y_18_c42, Y_18_c43, Y_18_c44, Y_18_c45, Y_18_c46, Y_18_c47, Y_18_c48, Y_18_c49, Y_18_c50, Y_18_c51, Y_18_c52 :  std_logic_vector(3 downto 0);
signal S_18_c52 :  std_logic_vector(3 downto 0);
signal R_18_c52, R_18_c53, R_18_c54, R_18_c55, R_18_c56 :  std_logic_vector(2 downto 0);
signal Cin_19_c52, Cin_19_c53 :  std_logic;
signal X_19_c33, X_19_c34, X_19_c35, X_19_c36, X_19_c37, X_19_c38, X_19_c39, X_19_c40, X_19_c41, X_19_c42, X_19_c43, X_19_c44, X_19_c45, X_19_c46, X_19_c47, X_19_c48, X_19_c49, X_19_c50, X_19_c51, X_19_c52, X_19_c53 :  std_logic_vector(3 downto 0);
signal Y_19_c0, Y_19_c1, Y_19_c2, Y_19_c3, Y_19_c4, Y_19_c5, Y_19_c6, Y_19_c7, Y_19_c8, Y_19_c9, Y_19_c10, Y_19_c11, Y_19_c12, Y_19_c13, Y_19_c14, Y_19_c15, Y_19_c16, Y_19_c17, Y_19_c18, Y_19_c19, Y_19_c20, Y_19_c21, Y_19_c22, Y_19_c23, Y_19_c24, Y_19_c25, Y_19_c26, Y_19_c27, Y_19_c28, Y_19_c29, Y_19_c30, Y_19_c31, Y_19_c32, Y_19_c33, Y_19_c34, Y_19_c35, Y_19_c36, Y_19_c37, Y_19_c38, Y_19_c39, Y_19_c40, Y_19_c41, Y_19_c42, Y_19_c43, Y_19_c44, Y_19_c45, Y_19_c46, Y_19_c47, Y_19_c48, Y_19_c49, Y_19_c50, Y_19_c51, Y_19_c52, Y_19_c53 :  std_logic_vector(3 downto 0);
signal S_19_c53 :  std_logic_vector(3 downto 0);
signal R_19_c53, R_19_c54, R_19_c55, R_19_c56 :  std_logic_vector(2 downto 0);
signal Cin_20_c53, Cin_20_c54 :  std_logic;
signal X_20_c33, X_20_c34, X_20_c35, X_20_c36, X_20_c37, X_20_c38, X_20_c39, X_20_c40, X_20_c41, X_20_c42, X_20_c43, X_20_c44, X_20_c45, X_20_c46, X_20_c47, X_20_c48, X_20_c49, X_20_c50, X_20_c51, X_20_c52, X_20_c53, X_20_c54 :  std_logic_vector(3 downto 0);
signal Y_20_c0, Y_20_c1, Y_20_c2, Y_20_c3, Y_20_c4, Y_20_c5, Y_20_c6, Y_20_c7, Y_20_c8, Y_20_c9, Y_20_c10, Y_20_c11, Y_20_c12, Y_20_c13, Y_20_c14, Y_20_c15, Y_20_c16, Y_20_c17, Y_20_c18, Y_20_c19, Y_20_c20, Y_20_c21, Y_20_c22, Y_20_c23, Y_20_c24, Y_20_c25, Y_20_c26, Y_20_c27, Y_20_c28, Y_20_c29, Y_20_c30, Y_20_c31, Y_20_c32, Y_20_c33, Y_20_c34, Y_20_c35, Y_20_c36, Y_20_c37, Y_20_c38, Y_20_c39, Y_20_c40, Y_20_c41, Y_20_c42, Y_20_c43, Y_20_c44, Y_20_c45, Y_20_c46, Y_20_c47, Y_20_c48, Y_20_c49, Y_20_c50, Y_20_c51, Y_20_c52, Y_20_c53, Y_20_c54 :  std_logic_vector(3 downto 0);
signal S_20_c54 :  std_logic_vector(3 downto 0);
signal R_20_c54, R_20_c55, R_20_c56 :  std_logic_vector(2 downto 0);
signal Cin_21_c54, Cin_21_c55, Cin_21_c56 :  std_logic;
signal X_21_c33, X_21_c34, X_21_c35, X_21_c36, X_21_c37, X_21_c38, X_21_c39, X_21_c40, X_21_c41, X_21_c42, X_21_c43, X_21_c44, X_21_c45, X_21_c46, X_21_c47, X_21_c48, X_21_c49, X_21_c50, X_21_c51, X_21_c52, X_21_c53, X_21_c54, X_21_c55, X_21_c56 :  std_logic_vector(3 downto 0);
signal Y_21_c0, Y_21_c1, Y_21_c2, Y_21_c3, Y_21_c4, Y_21_c5, Y_21_c6, Y_21_c7, Y_21_c8, Y_21_c9, Y_21_c10, Y_21_c11, Y_21_c12, Y_21_c13, Y_21_c14, Y_21_c15, Y_21_c16, Y_21_c17, Y_21_c18, Y_21_c19, Y_21_c20, Y_21_c21, Y_21_c22, Y_21_c23, Y_21_c24, Y_21_c25, Y_21_c26, Y_21_c27, Y_21_c28, Y_21_c29, Y_21_c30, Y_21_c31, Y_21_c32, Y_21_c33, Y_21_c34, Y_21_c35, Y_21_c36, Y_21_c37, Y_21_c38, Y_21_c39, Y_21_c40, Y_21_c41, Y_21_c42, Y_21_c43, Y_21_c44, Y_21_c45, Y_21_c46, Y_21_c47, Y_21_c48, Y_21_c49, Y_21_c50, Y_21_c51, Y_21_c52, Y_21_c53, Y_21_c54, Y_21_c55, Y_21_c56 :  std_logic_vector(3 downto 0);
signal S_21_c56 :  std_logic_vector(3 downto 0);
signal R_21_c56 :  std_logic_vector(2 downto 0);
signal Cin_22_c56 :  std_logic;
signal X_22_c33, X_22_c34, X_22_c35, X_22_c36, X_22_c37, X_22_c38, X_22_c39, X_22_c40, X_22_c41, X_22_c42, X_22_c43, X_22_c44, X_22_c45, X_22_c46, X_22_c47, X_22_c48, X_22_c49, X_22_c50, X_22_c51, X_22_c52, X_22_c53, X_22_c54, X_22_c55, X_22_c56 :  std_logic_vector(2 downto 0);
signal Y_22_c0, Y_22_c1, Y_22_c2, Y_22_c3, Y_22_c4, Y_22_c5, Y_22_c6, Y_22_c7, Y_22_c8, Y_22_c9, Y_22_c10, Y_22_c11, Y_22_c12, Y_22_c13, Y_22_c14, Y_22_c15, Y_22_c16, Y_22_c17, Y_22_c18, Y_22_c19, Y_22_c20, Y_22_c21, Y_22_c22, Y_22_c23, Y_22_c24, Y_22_c25, Y_22_c26, Y_22_c27, Y_22_c28, Y_22_c29, Y_22_c30, Y_22_c31, Y_22_c32, Y_22_c33, Y_22_c34, Y_22_c35, Y_22_c36, Y_22_c37, Y_22_c38, Y_22_c39, Y_22_c40, Y_22_c41, Y_22_c42, Y_22_c43, Y_22_c44, Y_22_c45, Y_22_c46, Y_22_c47, Y_22_c48, Y_22_c49, Y_22_c50, Y_22_c51, Y_22_c52, Y_22_c53, Y_22_c54, Y_22_c55, Y_22_c56 :  std_logic_vector(2 downto 0);
signal S_22_c56 :  std_logic_vector(2 downto 0);
signal R_22_c56 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_1_c1 <= Y_1_c0;
               Y_2_c1 <= Y_2_c0;
               Y_3_c1 <= Y_3_c0;
               Y_4_c1 <= Y_4_c0;
               Y_5_c1 <= Y_5_c0;
               Y_6_c1 <= Y_6_c0;
               Y_7_c1 <= Y_7_c0;
               Y_8_c1 <= Y_8_c0;
               Y_9_c1 <= Y_9_c0;
               Y_10_c1 <= Y_10_c0;
               Y_11_c1 <= Y_11_c0;
               Y_12_c1 <= Y_12_c0;
               Y_13_c1 <= Y_13_c0;
               Y_14_c1 <= Y_14_c0;
               Y_15_c1 <= Y_15_c0;
               Y_16_c1 <= Y_16_c0;
               Y_17_c1 <= Y_17_c0;
               Y_18_c1 <= Y_18_c0;
               Y_19_c1 <= Y_19_c0;
               Y_20_c1 <= Y_20_c0;
               Y_21_c1 <= Y_21_c0;
               Y_22_c1 <= Y_22_c0;
            end if;
            if ce_2 = '1' then
               Y_1_c2 <= Y_1_c1;
               Y_2_c2 <= Y_2_c1;
               Y_3_c2 <= Y_3_c1;
               Y_4_c2 <= Y_4_c1;
               Y_5_c2 <= Y_5_c1;
               Y_6_c2 <= Y_6_c1;
               Y_7_c2 <= Y_7_c1;
               Y_8_c2 <= Y_8_c1;
               Y_9_c2 <= Y_9_c1;
               Y_10_c2 <= Y_10_c1;
               Y_11_c2 <= Y_11_c1;
               Y_12_c2 <= Y_12_c1;
               Y_13_c2 <= Y_13_c1;
               Y_14_c2 <= Y_14_c1;
               Y_15_c2 <= Y_15_c1;
               Y_16_c2 <= Y_16_c1;
               Y_17_c2 <= Y_17_c1;
               Y_18_c2 <= Y_18_c1;
               Y_19_c2 <= Y_19_c1;
               Y_20_c2 <= Y_20_c1;
               Y_21_c2 <= Y_21_c1;
               Y_22_c2 <= Y_22_c1;
            end if;
            if ce_3 = '1' then
               Y_1_c3 <= Y_1_c2;
               Y_2_c3 <= Y_2_c2;
               Y_3_c3 <= Y_3_c2;
               Y_4_c3 <= Y_4_c2;
               Y_5_c3 <= Y_5_c2;
               Y_6_c3 <= Y_6_c2;
               Y_7_c3 <= Y_7_c2;
               Y_8_c3 <= Y_8_c2;
               Y_9_c3 <= Y_9_c2;
               Y_10_c3 <= Y_10_c2;
               Y_11_c3 <= Y_11_c2;
               Y_12_c3 <= Y_12_c2;
               Y_13_c3 <= Y_13_c2;
               Y_14_c3 <= Y_14_c2;
               Y_15_c3 <= Y_15_c2;
               Y_16_c3 <= Y_16_c2;
               Y_17_c3 <= Y_17_c2;
               Y_18_c3 <= Y_18_c2;
               Y_19_c3 <= Y_19_c2;
               Y_20_c3 <= Y_20_c2;
               Y_21_c3 <= Y_21_c2;
               Y_22_c3 <= Y_22_c2;
            end if;
            if ce_4 = '1' then
               Y_1_c4 <= Y_1_c3;
               Y_2_c4 <= Y_2_c3;
               Y_3_c4 <= Y_3_c3;
               Y_4_c4 <= Y_4_c3;
               Y_5_c4 <= Y_5_c3;
               Y_6_c4 <= Y_6_c3;
               Y_7_c4 <= Y_7_c3;
               Y_8_c4 <= Y_8_c3;
               Y_9_c4 <= Y_9_c3;
               Y_10_c4 <= Y_10_c3;
               Y_11_c4 <= Y_11_c3;
               Y_12_c4 <= Y_12_c3;
               Y_13_c4 <= Y_13_c3;
               Y_14_c4 <= Y_14_c3;
               Y_15_c4 <= Y_15_c3;
               Y_16_c4 <= Y_16_c3;
               Y_17_c4 <= Y_17_c3;
               Y_18_c4 <= Y_18_c3;
               Y_19_c4 <= Y_19_c3;
               Y_20_c4 <= Y_20_c3;
               Y_21_c4 <= Y_21_c3;
               Y_22_c4 <= Y_22_c3;
            end if;
            if ce_5 = '1' then
               Y_1_c5 <= Y_1_c4;
               Y_2_c5 <= Y_2_c4;
               Y_3_c5 <= Y_3_c4;
               Y_4_c5 <= Y_4_c4;
               Y_5_c5 <= Y_5_c4;
               Y_6_c5 <= Y_6_c4;
               Y_7_c5 <= Y_7_c4;
               Y_8_c5 <= Y_8_c4;
               Y_9_c5 <= Y_9_c4;
               Y_10_c5 <= Y_10_c4;
               Y_11_c5 <= Y_11_c4;
               Y_12_c5 <= Y_12_c4;
               Y_13_c5 <= Y_13_c4;
               Y_14_c5 <= Y_14_c4;
               Y_15_c5 <= Y_15_c4;
               Y_16_c5 <= Y_16_c4;
               Y_17_c5 <= Y_17_c4;
               Y_18_c5 <= Y_18_c4;
               Y_19_c5 <= Y_19_c4;
               Y_20_c5 <= Y_20_c4;
               Y_21_c5 <= Y_21_c4;
               Y_22_c5 <= Y_22_c4;
            end if;
            if ce_6 = '1' then
               Y_1_c6 <= Y_1_c5;
               Y_2_c6 <= Y_2_c5;
               Y_3_c6 <= Y_3_c5;
               Y_4_c6 <= Y_4_c5;
               Y_5_c6 <= Y_5_c5;
               Y_6_c6 <= Y_6_c5;
               Y_7_c6 <= Y_7_c5;
               Y_8_c6 <= Y_8_c5;
               Y_9_c6 <= Y_9_c5;
               Y_10_c6 <= Y_10_c5;
               Y_11_c6 <= Y_11_c5;
               Y_12_c6 <= Y_12_c5;
               Y_13_c6 <= Y_13_c5;
               Y_14_c6 <= Y_14_c5;
               Y_15_c6 <= Y_15_c5;
               Y_16_c6 <= Y_16_c5;
               Y_17_c6 <= Y_17_c5;
               Y_18_c6 <= Y_18_c5;
               Y_19_c6 <= Y_19_c5;
               Y_20_c6 <= Y_20_c5;
               Y_21_c6 <= Y_21_c5;
               Y_22_c6 <= Y_22_c5;
            end if;
            if ce_7 = '1' then
               Y_1_c7 <= Y_1_c6;
               Y_2_c7 <= Y_2_c6;
               Y_3_c7 <= Y_3_c6;
               Y_4_c7 <= Y_4_c6;
               Y_5_c7 <= Y_5_c6;
               Y_6_c7 <= Y_6_c6;
               Y_7_c7 <= Y_7_c6;
               Y_8_c7 <= Y_8_c6;
               Y_9_c7 <= Y_9_c6;
               Y_10_c7 <= Y_10_c6;
               Y_11_c7 <= Y_11_c6;
               Y_12_c7 <= Y_12_c6;
               Y_13_c7 <= Y_13_c6;
               Y_14_c7 <= Y_14_c6;
               Y_15_c7 <= Y_15_c6;
               Y_16_c7 <= Y_16_c6;
               Y_17_c7 <= Y_17_c6;
               Y_18_c7 <= Y_18_c6;
               Y_19_c7 <= Y_19_c6;
               Y_20_c7 <= Y_20_c6;
               Y_21_c7 <= Y_21_c6;
               Y_22_c7 <= Y_22_c6;
            end if;
            if ce_8 = '1' then
               Y_1_c8 <= Y_1_c7;
               Y_2_c8 <= Y_2_c7;
               Y_3_c8 <= Y_3_c7;
               Y_4_c8 <= Y_4_c7;
               Y_5_c8 <= Y_5_c7;
               Y_6_c8 <= Y_6_c7;
               Y_7_c8 <= Y_7_c7;
               Y_8_c8 <= Y_8_c7;
               Y_9_c8 <= Y_9_c7;
               Y_10_c8 <= Y_10_c7;
               Y_11_c8 <= Y_11_c7;
               Y_12_c8 <= Y_12_c7;
               Y_13_c8 <= Y_13_c7;
               Y_14_c8 <= Y_14_c7;
               Y_15_c8 <= Y_15_c7;
               Y_16_c8 <= Y_16_c7;
               Y_17_c8 <= Y_17_c7;
               Y_18_c8 <= Y_18_c7;
               Y_19_c8 <= Y_19_c7;
               Y_20_c8 <= Y_20_c7;
               Y_21_c8 <= Y_21_c7;
               Y_22_c8 <= Y_22_c7;
            end if;
            if ce_9 = '1' then
               Y_1_c9 <= Y_1_c8;
               Y_2_c9 <= Y_2_c8;
               Y_3_c9 <= Y_3_c8;
               Y_4_c9 <= Y_4_c8;
               Y_5_c9 <= Y_5_c8;
               Y_6_c9 <= Y_6_c8;
               Y_7_c9 <= Y_7_c8;
               Y_8_c9 <= Y_8_c8;
               Y_9_c9 <= Y_9_c8;
               Y_10_c9 <= Y_10_c8;
               Y_11_c9 <= Y_11_c8;
               Y_12_c9 <= Y_12_c8;
               Y_13_c9 <= Y_13_c8;
               Y_14_c9 <= Y_14_c8;
               Y_15_c9 <= Y_15_c8;
               Y_16_c9 <= Y_16_c8;
               Y_17_c9 <= Y_17_c8;
               Y_18_c9 <= Y_18_c8;
               Y_19_c9 <= Y_19_c8;
               Y_20_c9 <= Y_20_c8;
               Y_21_c9 <= Y_21_c8;
               Y_22_c9 <= Y_22_c8;
            end if;
            if ce_10 = '1' then
               Y_1_c10 <= Y_1_c9;
               Y_2_c10 <= Y_2_c9;
               Y_3_c10 <= Y_3_c9;
               Y_4_c10 <= Y_4_c9;
               Y_5_c10 <= Y_5_c9;
               Y_6_c10 <= Y_6_c9;
               Y_7_c10 <= Y_7_c9;
               Y_8_c10 <= Y_8_c9;
               Y_9_c10 <= Y_9_c9;
               Y_10_c10 <= Y_10_c9;
               Y_11_c10 <= Y_11_c9;
               Y_12_c10 <= Y_12_c9;
               Y_13_c10 <= Y_13_c9;
               Y_14_c10 <= Y_14_c9;
               Y_15_c10 <= Y_15_c9;
               Y_16_c10 <= Y_16_c9;
               Y_17_c10 <= Y_17_c9;
               Y_18_c10 <= Y_18_c9;
               Y_19_c10 <= Y_19_c9;
               Y_20_c10 <= Y_20_c9;
               Y_21_c10 <= Y_21_c9;
               Y_22_c10 <= Y_22_c9;
            end if;
            if ce_11 = '1' then
               Y_1_c11 <= Y_1_c10;
               Y_2_c11 <= Y_2_c10;
               Y_3_c11 <= Y_3_c10;
               Y_4_c11 <= Y_4_c10;
               Y_5_c11 <= Y_5_c10;
               Y_6_c11 <= Y_6_c10;
               Y_7_c11 <= Y_7_c10;
               Y_8_c11 <= Y_8_c10;
               Y_9_c11 <= Y_9_c10;
               Y_10_c11 <= Y_10_c10;
               Y_11_c11 <= Y_11_c10;
               Y_12_c11 <= Y_12_c10;
               Y_13_c11 <= Y_13_c10;
               Y_14_c11 <= Y_14_c10;
               Y_15_c11 <= Y_15_c10;
               Y_16_c11 <= Y_16_c10;
               Y_17_c11 <= Y_17_c10;
               Y_18_c11 <= Y_18_c10;
               Y_19_c11 <= Y_19_c10;
               Y_20_c11 <= Y_20_c10;
               Y_21_c11 <= Y_21_c10;
               Y_22_c11 <= Y_22_c10;
            end if;
            if ce_12 = '1' then
               Y_1_c12 <= Y_1_c11;
               Y_2_c12 <= Y_2_c11;
               Y_3_c12 <= Y_3_c11;
               Y_4_c12 <= Y_4_c11;
               Y_5_c12 <= Y_5_c11;
               Y_6_c12 <= Y_6_c11;
               Y_7_c12 <= Y_7_c11;
               Y_8_c12 <= Y_8_c11;
               Y_9_c12 <= Y_9_c11;
               Y_10_c12 <= Y_10_c11;
               Y_11_c12 <= Y_11_c11;
               Y_12_c12 <= Y_12_c11;
               Y_13_c12 <= Y_13_c11;
               Y_14_c12 <= Y_14_c11;
               Y_15_c12 <= Y_15_c11;
               Y_16_c12 <= Y_16_c11;
               Y_17_c12 <= Y_17_c11;
               Y_18_c12 <= Y_18_c11;
               Y_19_c12 <= Y_19_c11;
               Y_20_c12 <= Y_20_c11;
               Y_21_c12 <= Y_21_c11;
               Y_22_c12 <= Y_22_c11;
            end if;
            if ce_13 = '1' then
               Y_1_c13 <= Y_1_c12;
               Y_2_c13 <= Y_2_c12;
               Y_3_c13 <= Y_3_c12;
               Y_4_c13 <= Y_4_c12;
               Y_5_c13 <= Y_5_c12;
               Y_6_c13 <= Y_6_c12;
               Y_7_c13 <= Y_7_c12;
               Y_8_c13 <= Y_8_c12;
               Y_9_c13 <= Y_9_c12;
               Y_10_c13 <= Y_10_c12;
               Y_11_c13 <= Y_11_c12;
               Y_12_c13 <= Y_12_c12;
               Y_13_c13 <= Y_13_c12;
               Y_14_c13 <= Y_14_c12;
               Y_15_c13 <= Y_15_c12;
               Y_16_c13 <= Y_16_c12;
               Y_17_c13 <= Y_17_c12;
               Y_18_c13 <= Y_18_c12;
               Y_19_c13 <= Y_19_c12;
               Y_20_c13 <= Y_20_c12;
               Y_21_c13 <= Y_21_c12;
               Y_22_c13 <= Y_22_c12;
            end if;
            if ce_14 = '1' then
               Y_1_c14 <= Y_1_c13;
               Y_2_c14 <= Y_2_c13;
               Y_3_c14 <= Y_3_c13;
               Y_4_c14 <= Y_4_c13;
               Y_5_c14 <= Y_5_c13;
               Y_6_c14 <= Y_6_c13;
               Y_7_c14 <= Y_7_c13;
               Y_8_c14 <= Y_8_c13;
               Y_9_c14 <= Y_9_c13;
               Y_10_c14 <= Y_10_c13;
               Y_11_c14 <= Y_11_c13;
               Y_12_c14 <= Y_12_c13;
               Y_13_c14 <= Y_13_c13;
               Y_14_c14 <= Y_14_c13;
               Y_15_c14 <= Y_15_c13;
               Y_16_c14 <= Y_16_c13;
               Y_17_c14 <= Y_17_c13;
               Y_18_c14 <= Y_18_c13;
               Y_19_c14 <= Y_19_c13;
               Y_20_c14 <= Y_20_c13;
               Y_21_c14 <= Y_21_c13;
               Y_22_c14 <= Y_22_c13;
            end if;
            if ce_15 = '1' then
               Y_1_c15 <= Y_1_c14;
               Y_2_c15 <= Y_2_c14;
               Y_3_c15 <= Y_3_c14;
               Y_4_c15 <= Y_4_c14;
               Y_5_c15 <= Y_5_c14;
               Y_6_c15 <= Y_6_c14;
               Y_7_c15 <= Y_7_c14;
               Y_8_c15 <= Y_8_c14;
               Y_9_c15 <= Y_9_c14;
               Y_10_c15 <= Y_10_c14;
               Y_11_c15 <= Y_11_c14;
               Y_12_c15 <= Y_12_c14;
               Y_13_c15 <= Y_13_c14;
               Y_14_c15 <= Y_14_c14;
               Y_15_c15 <= Y_15_c14;
               Y_16_c15 <= Y_16_c14;
               Y_17_c15 <= Y_17_c14;
               Y_18_c15 <= Y_18_c14;
               Y_19_c15 <= Y_19_c14;
               Y_20_c15 <= Y_20_c14;
               Y_21_c15 <= Y_21_c14;
               Y_22_c15 <= Y_22_c14;
            end if;
            if ce_16 = '1' then
               Y_1_c16 <= Y_1_c15;
               Y_2_c16 <= Y_2_c15;
               Y_3_c16 <= Y_3_c15;
               Y_4_c16 <= Y_4_c15;
               Y_5_c16 <= Y_5_c15;
               Y_6_c16 <= Y_6_c15;
               Y_7_c16 <= Y_7_c15;
               Y_8_c16 <= Y_8_c15;
               Y_9_c16 <= Y_9_c15;
               Y_10_c16 <= Y_10_c15;
               Y_11_c16 <= Y_11_c15;
               Y_12_c16 <= Y_12_c15;
               Y_13_c16 <= Y_13_c15;
               Y_14_c16 <= Y_14_c15;
               Y_15_c16 <= Y_15_c15;
               Y_16_c16 <= Y_16_c15;
               Y_17_c16 <= Y_17_c15;
               Y_18_c16 <= Y_18_c15;
               Y_19_c16 <= Y_19_c15;
               Y_20_c16 <= Y_20_c15;
               Y_21_c16 <= Y_21_c15;
               Y_22_c16 <= Y_22_c15;
            end if;
            if ce_17 = '1' then
               Y_1_c17 <= Y_1_c16;
               Y_2_c17 <= Y_2_c16;
               Y_3_c17 <= Y_3_c16;
               Y_4_c17 <= Y_4_c16;
               Y_5_c17 <= Y_5_c16;
               Y_6_c17 <= Y_6_c16;
               Y_7_c17 <= Y_7_c16;
               Y_8_c17 <= Y_8_c16;
               Y_9_c17 <= Y_9_c16;
               Y_10_c17 <= Y_10_c16;
               Y_11_c17 <= Y_11_c16;
               Y_12_c17 <= Y_12_c16;
               Y_13_c17 <= Y_13_c16;
               Y_14_c17 <= Y_14_c16;
               Y_15_c17 <= Y_15_c16;
               Y_16_c17 <= Y_16_c16;
               Y_17_c17 <= Y_17_c16;
               Y_18_c17 <= Y_18_c16;
               Y_19_c17 <= Y_19_c16;
               Y_20_c17 <= Y_20_c16;
               Y_21_c17 <= Y_21_c16;
               Y_22_c17 <= Y_22_c16;
            end if;
            if ce_18 = '1' then
               Y_1_c18 <= Y_1_c17;
               Y_2_c18 <= Y_2_c17;
               Y_3_c18 <= Y_3_c17;
               Y_4_c18 <= Y_4_c17;
               Y_5_c18 <= Y_5_c17;
               Y_6_c18 <= Y_6_c17;
               Y_7_c18 <= Y_7_c17;
               Y_8_c18 <= Y_8_c17;
               Y_9_c18 <= Y_9_c17;
               Y_10_c18 <= Y_10_c17;
               Y_11_c18 <= Y_11_c17;
               Y_12_c18 <= Y_12_c17;
               Y_13_c18 <= Y_13_c17;
               Y_14_c18 <= Y_14_c17;
               Y_15_c18 <= Y_15_c17;
               Y_16_c18 <= Y_16_c17;
               Y_17_c18 <= Y_17_c17;
               Y_18_c18 <= Y_18_c17;
               Y_19_c18 <= Y_19_c17;
               Y_20_c18 <= Y_20_c17;
               Y_21_c18 <= Y_21_c17;
               Y_22_c18 <= Y_22_c17;
            end if;
            if ce_19 = '1' then
               Y_1_c19 <= Y_1_c18;
               Y_2_c19 <= Y_2_c18;
               Y_3_c19 <= Y_3_c18;
               Y_4_c19 <= Y_4_c18;
               Y_5_c19 <= Y_5_c18;
               Y_6_c19 <= Y_6_c18;
               Y_7_c19 <= Y_7_c18;
               Y_8_c19 <= Y_8_c18;
               Y_9_c19 <= Y_9_c18;
               Y_10_c19 <= Y_10_c18;
               Y_11_c19 <= Y_11_c18;
               Y_12_c19 <= Y_12_c18;
               Y_13_c19 <= Y_13_c18;
               Y_14_c19 <= Y_14_c18;
               Y_15_c19 <= Y_15_c18;
               Y_16_c19 <= Y_16_c18;
               Y_17_c19 <= Y_17_c18;
               Y_18_c19 <= Y_18_c18;
               Y_19_c19 <= Y_19_c18;
               Y_20_c19 <= Y_20_c18;
               Y_21_c19 <= Y_21_c18;
               Y_22_c19 <= Y_22_c18;
            end if;
            if ce_20 = '1' then
               Y_1_c20 <= Y_1_c19;
               Y_2_c20 <= Y_2_c19;
               Y_3_c20 <= Y_3_c19;
               Y_4_c20 <= Y_4_c19;
               Y_5_c20 <= Y_5_c19;
               Y_6_c20 <= Y_6_c19;
               Y_7_c20 <= Y_7_c19;
               Y_8_c20 <= Y_8_c19;
               Y_9_c20 <= Y_9_c19;
               Y_10_c20 <= Y_10_c19;
               Y_11_c20 <= Y_11_c19;
               Y_12_c20 <= Y_12_c19;
               Y_13_c20 <= Y_13_c19;
               Y_14_c20 <= Y_14_c19;
               Y_15_c20 <= Y_15_c19;
               Y_16_c20 <= Y_16_c19;
               Y_17_c20 <= Y_17_c19;
               Y_18_c20 <= Y_18_c19;
               Y_19_c20 <= Y_19_c19;
               Y_20_c20 <= Y_20_c19;
               Y_21_c20 <= Y_21_c19;
               Y_22_c20 <= Y_22_c19;
            end if;
            if ce_21 = '1' then
               Y_1_c21 <= Y_1_c20;
               Y_2_c21 <= Y_2_c20;
               Y_3_c21 <= Y_3_c20;
               Y_4_c21 <= Y_4_c20;
               Y_5_c21 <= Y_5_c20;
               Y_6_c21 <= Y_6_c20;
               Y_7_c21 <= Y_7_c20;
               Y_8_c21 <= Y_8_c20;
               Y_9_c21 <= Y_9_c20;
               Y_10_c21 <= Y_10_c20;
               Y_11_c21 <= Y_11_c20;
               Y_12_c21 <= Y_12_c20;
               Y_13_c21 <= Y_13_c20;
               Y_14_c21 <= Y_14_c20;
               Y_15_c21 <= Y_15_c20;
               Y_16_c21 <= Y_16_c20;
               Y_17_c21 <= Y_17_c20;
               Y_18_c21 <= Y_18_c20;
               Y_19_c21 <= Y_19_c20;
               Y_20_c21 <= Y_20_c20;
               Y_21_c21 <= Y_21_c20;
               Y_22_c21 <= Y_22_c20;
            end if;
            if ce_22 = '1' then
               Y_1_c22 <= Y_1_c21;
               Y_2_c22 <= Y_2_c21;
               Y_3_c22 <= Y_3_c21;
               Y_4_c22 <= Y_4_c21;
               Y_5_c22 <= Y_5_c21;
               Y_6_c22 <= Y_6_c21;
               Y_7_c22 <= Y_7_c21;
               Y_8_c22 <= Y_8_c21;
               Y_9_c22 <= Y_9_c21;
               Y_10_c22 <= Y_10_c21;
               Y_11_c22 <= Y_11_c21;
               Y_12_c22 <= Y_12_c21;
               Y_13_c22 <= Y_13_c21;
               Y_14_c22 <= Y_14_c21;
               Y_15_c22 <= Y_15_c21;
               Y_16_c22 <= Y_16_c21;
               Y_17_c22 <= Y_17_c21;
               Y_18_c22 <= Y_18_c21;
               Y_19_c22 <= Y_19_c21;
               Y_20_c22 <= Y_20_c21;
               Y_21_c22 <= Y_21_c21;
               Y_22_c22 <= Y_22_c21;
            end if;
            if ce_23 = '1' then
               Y_1_c23 <= Y_1_c22;
               Y_2_c23 <= Y_2_c22;
               Y_3_c23 <= Y_3_c22;
               Y_4_c23 <= Y_4_c22;
               Y_5_c23 <= Y_5_c22;
               Y_6_c23 <= Y_6_c22;
               Y_7_c23 <= Y_7_c22;
               Y_8_c23 <= Y_8_c22;
               Y_9_c23 <= Y_9_c22;
               Y_10_c23 <= Y_10_c22;
               Y_11_c23 <= Y_11_c22;
               Y_12_c23 <= Y_12_c22;
               Y_13_c23 <= Y_13_c22;
               Y_14_c23 <= Y_14_c22;
               Y_15_c23 <= Y_15_c22;
               Y_16_c23 <= Y_16_c22;
               Y_17_c23 <= Y_17_c22;
               Y_18_c23 <= Y_18_c22;
               Y_19_c23 <= Y_19_c22;
               Y_20_c23 <= Y_20_c22;
               Y_21_c23 <= Y_21_c22;
               Y_22_c23 <= Y_22_c22;
            end if;
            if ce_24 = '1' then
               Y_1_c24 <= Y_1_c23;
               Y_2_c24 <= Y_2_c23;
               Y_3_c24 <= Y_3_c23;
               Y_4_c24 <= Y_4_c23;
               Y_5_c24 <= Y_5_c23;
               Y_6_c24 <= Y_6_c23;
               Y_7_c24 <= Y_7_c23;
               Y_8_c24 <= Y_8_c23;
               Y_9_c24 <= Y_9_c23;
               Y_10_c24 <= Y_10_c23;
               Y_11_c24 <= Y_11_c23;
               Y_12_c24 <= Y_12_c23;
               Y_13_c24 <= Y_13_c23;
               Y_14_c24 <= Y_14_c23;
               Y_15_c24 <= Y_15_c23;
               Y_16_c24 <= Y_16_c23;
               Y_17_c24 <= Y_17_c23;
               Y_18_c24 <= Y_18_c23;
               Y_19_c24 <= Y_19_c23;
               Y_20_c24 <= Y_20_c23;
               Y_21_c24 <= Y_21_c23;
               Y_22_c24 <= Y_22_c23;
            end if;
            if ce_25 = '1' then
               Y_1_c25 <= Y_1_c24;
               Y_2_c25 <= Y_2_c24;
               Y_3_c25 <= Y_3_c24;
               Y_4_c25 <= Y_4_c24;
               Y_5_c25 <= Y_5_c24;
               Y_6_c25 <= Y_6_c24;
               Y_7_c25 <= Y_7_c24;
               Y_8_c25 <= Y_8_c24;
               Y_9_c25 <= Y_9_c24;
               Y_10_c25 <= Y_10_c24;
               Y_11_c25 <= Y_11_c24;
               Y_12_c25 <= Y_12_c24;
               Y_13_c25 <= Y_13_c24;
               Y_14_c25 <= Y_14_c24;
               Y_15_c25 <= Y_15_c24;
               Y_16_c25 <= Y_16_c24;
               Y_17_c25 <= Y_17_c24;
               Y_18_c25 <= Y_18_c24;
               Y_19_c25 <= Y_19_c24;
               Y_20_c25 <= Y_20_c24;
               Y_21_c25 <= Y_21_c24;
               Y_22_c25 <= Y_22_c24;
            end if;
            if ce_26 = '1' then
               Y_1_c26 <= Y_1_c25;
               Y_2_c26 <= Y_2_c25;
               Y_3_c26 <= Y_3_c25;
               Y_4_c26 <= Y_4_c25;
               Y_5_c26 <= Y_5_c25;
               Y_6_c26 <= Y_6_c25;
               Y_7_c26 <= Y_7_c25;
               Y_8_c26 <= Y_8_c25;
               Y_9_c26 <= Y_9_c25;
               Y_10_c26 <= Y_10_c25;
               Y_11_c26 <= Y_11_c25;
               Y_12_c26 <= Y_12_c25;
               Y_13_c26 <= Y_13_c25;
               Y_14_c26 <= Y_14_c25;
               Y_15_c26 <= Y_15_c25;
               Y_16_c26 <= Y_16_c25;
               Y_17_c26 <= Y_17_c25;
               Y_18_c26 <= Y_18_c25;
               Y_19_c26 <= Y_19_c25;
               Y_20_c26 <= Y_20_c25;
               Y_21_c26 <= Y_21_c25;
               Y_22_c26 <= Y_22_c25;
            end if;
            if ce_27 = '1' then
               Y_1_c27 <= Y_1_c26;
               Y_2_c27 <= Y_2_c26;
               Y_3_c27 <= Y_3_c26;
               Y_4_c27 <= Y_4_c26;
               Y_5_c27 <= Y_5_c26;
               Y_6_c27 <= Y_6_c26;
               Y_7_c27 <= Y_7_c26;
               Y_8_c27 <= Y_8_c26;
               Y_9_c27 <= Y_9_c26;
               Y_10_c27 <= Y_10_c26;
               Y_11_c27 <= Y_11_c26;
               Y_12_c27 <= Y_12_c26;
               Y_13_c27 <= Y_13_c26;
               Y_14_c27 <= Y_14_c26;
               Y_15_c27 <= Y_15_c26;
               Y_16_c27 <= Y_16_c26;
               Y_17_c27 <= Y_17_c26;
               Y_18_c27 <= Y_18_c26;
               Y_19_c27 <= Y_19_c26;
               Y_20_c27 <= Y_20_c26;
               Y_21_c27 <= Y_21_c26;
               Y_22_c27 <= Y_22_c26;
            end if;
            if ce_28 = '1' then
               Y_1_c28 <= Y_1_c27;
               Y_2_c28 <= Y_2_c27;
               Y_3_c28 <= Y_3_c27;
               Y_4_c28 <= Y_4_c27;
               Y_5_c28 <= Y_5_c27;
               Y_6_c28 <= Y_6_c27;
               Y_7_c28 <= Y_7_c27;
               Y_8_c28 <= Y_8_c27;
               Y_9_c28 <= Y_9_c27;
               Y_10_c28 <= Y_10_c27;
               Y_11_c28 <= Y_11_c27;
               Y_12_c28 <= Y_12_c27;
               Y_13_c28 <= Y_13_c27;
               Y_14_c28 <= Y_14_c27;
               Y_15_c28 <= Y_15_c27;
               Y_16_c28 <= Y_16_c27;
               Y_17_c28 <= Y_17_c27;
               Y_18_c28 <= Y_18_c27;
               Y_19_c28 <= Y_19_c27;
               Y_20_c28 <= Y_20_c27;
               Y_21_c28 <= Y_21_c27;
               Y_22_c28 <= Y_22_c27;
            end if;
            if ce_29 = '1' then
               Y_1_c29 <= Y_1_c28;
               Y_2_c29 <= Y_2_c28;
               Y_3_c29 <= Y_3_c28;
               Y_4_c29 <= Y_4_c28;
               Y_5_c29 <= Y_5_c28;
               Y_6_c29 <= Y_6_c28;
               Y_7_c29 <= Y_7_c28;
               Y_8_c29 <= Y_8_c28;
               Y_9_c29 <= Y_9_c28;
               Y_10_c29 <= Y_10_c28;
               Y_11_c29 <= Y_11_c28;
               Y_12_c29 <= Y_12_c28;
               Y_13_c29 <= Y_13_c28;
               Y_14_c29 <= Y_14_c28;
               Y_15_c29 <= Y_15_c28;
               Y_16_c29 <= Y_16_c28;
               Y_17_c29 <= Y_17_c28;
               Y_18_c29 <= Y_18_c28;
               Y_19_c29 <= Y_19_c28;
               Y_20_c29 <= Y_20_c28;
               Y_21_c29 <= Y_21_c28;
               Y_22_c29 <= Y_22_c28;
            end if;
            if ce_30 = '1' then
               Y_1_c30 <= Y_1_c29;
               Y_2_c30 <= Y_2_c29;
               Y_3_c30 <= Y_3_c29;
               Y_4_c30 <= Y_4_c29;
               Y_5_c30 <= Y_5_c29;
               Y_6_c30 <= Y_6_c29;
               Y_7_c30 <= Y_7_c29;
               Y_8_c30 <= Y_8_c29;
               Y_9_c30 <= Y_9_c29;
               Y_10_c30 <= Y_10_c29;
               Y_11_c30 <= Y_11_c29;
               Y_12_c30 <= Y_12_c29;
               Y_13_c30 <= Y_13_c29;
               Y_14_c30 <= Y_14_c29;
               Y_15_c30 <= Y_15_c29;
               Y_16_c30 <= Y_16_c29;
               Y_17_c30 <= Y_17_c29;
               Y_18_c30 <= Y_18_c29;
               Y_19_c30 <= Y_19_c29;
               Y_20_c30 <= Y_20_c29;
               Y_21_c30 <= Y_21_c29;
               Y_22_c30 <= Y_22_c29;
            end if;
            if ce_31 = '1' then
               Y_1_c31 <= Y_1_c30;
               Y_2_c31 <= Y_2_c30;
               Y_3_c31 <= Y_3_c30;
               Y_4_c31 <= Y_4_c30;
               Y_5_c31 <= Y_5_c30;
               Y_6_c31 <= Y_6_c30;
               Y_7_c31 <= Y_7_c30;
               Y_8_c31 <= Y_8_c30;
               Y_9_c31 <= Y_9_c30;
               Y_10_c31 <= Y_10_c30;
               Y_11_c31 <= Y_11_c30;
               Y_12_c31 <= Y_12_c30;
               Y_13_c31 <= Y_13_c30;
               Y_14_c31 <= Y_14_c30;
               Y_15_c31 <= Y_15_c30;
               Y_16_c31 <= Y_16_c30;
               Y_17_c31 <= Y_17_c30;
               Y_18_c31 <= Y_18_c30;
               Y_19_c31 <= Y_19_c30;
               Y_20_c31 <= Y_20_c30;
               Y_21_c31 <= Y_21_c30;
               Y_22_c31 <= Y_22_c30;
            end if;
            if ce_32 = '1' then
               Y_1_c32 <= Y_1_c31;
               Y_2_c32 <= Y_2_c31;
               Y_3_c32 <= Y_3_c31;
               Y_4_c32 <= Y_4_c31;
               Y_5_c32 <= Y_5_c31;
               Y_6_c32 <= Y_6_c31;
               Y_7_c32 <= Y_7_c31;
               Y_8_c32 <= Y_8_c31;
               Y_9_c32 <= Y_9_c31;
               Y_10_c32 <= Y_10_c31;
               Y_11_c32 <= Y_11_c31;
               Y_12_c32 <= Y_12_c31;
               Y_13_c32 <= Y_13_c31;
               Y_14_c32 <= Y_14_c31;
               Y_15_c32 <= Y_15_c31;
               Y_16_c32 <= Y_16_c31;
               Y_17_c32 <= Y_17_c31;
               Y_18_c32 <= Y_18_c31;
               Y_19_c32 <= Y_19_c31;
               Y_20_c32 <= Y_20_c31;
               Y_21_c32 <= Y_21_c31;
               Y_22_c32 <= Y_22_c31;
            end if;
            if ce_33 = '1' then
               Y_1_c33 <= Y_1_c32;
               Y_2_c33 <= Y_2_c32;
               Y_3_c33 <= Y_3_c32;
               Y_4_c33 <= Y_4_c32;
               Y_5_c33 <= Y_5_c32;
               Y_6_c33 <= Y_6_c32;
               Y_7_c33 <= Y_7_c32;
               Y_8_c33 <= Y_8_c32;
               Y_9_c33 <= Y_9_c32;
               Y_10_c33 <= Y_10_c32;
               Y_11_c33 <= Y_11_c32;
               Y_12_c33 <= Y_12_c32;
               Y_13_c33 <= Y_13_c32;
               Y_14_c33 <= Y_14_c32;
               Y_15_c33 <= Y_15_c32;
               Y_16_c33 <= Y_16_c32;
               Y_17_c33 <= Y_17_c32;
               Y_18_c33 <= Y_18_c32;
               Y_19_c33 <= Y_19_c32;
               Y_20_c33 <= Y_20_c32;
               Y_21_c33 <= Y_21_c32;
               Y_22_c33 <= Y_22_c32;
            end if;
            if ce_34 = '1' then
               X_1_c34 <= X_1_c33;
               Y_1_c34 <= Y_1_c33;
               X_2_c34 <= X_2_c33;
               Y_2_c34 <= Y_2_c33;
               X_3_c34 <= X_3_c33;
               Y_3_c34 <= Y_3_c33;
               X_4_c34 <= X_4_c33;
               Y_4_c34 <= Y_4_c33;
               X_5_c34 <= X_5_c33;
               Y_5_c34 <= Y_5_c33;
               X_6_c34 <= X_6_c33;
               Y_6_c34 <= Y_6_c33;
               X_7_c34 <= X_7_c33;
               Y_7_c34 <= Y_7_c33;
               X_8_c34 <= X_8_c33;
               Y_8_c34 <= Y_8_c33;
               X_9_c34 <= X_9_c33;
               Y_9_c34 <= Y_9_c33;
               X_10_c34 <= X_10_c33;
               Y_10_c34 <= Y_10_c33;
               X_11_c34 <= X_11_c33;
               Y_11_c34 <= Y_11_c33;
               X_12_c34 <= X_12_c33;
               Y_12_c34 <= Y_12_c33;
               X_13_c34 <= X_13_c33;
               Y_13_c34 <= Y_13_c33;
               X_14_c34 <= X_14_c33;
               Y_14_c34 <= Y_14_c33;
               X_15_c34 <= X_15_c33;
               Y_15_c34 <= Y_15_c33;
               X_16_c34 <= X_16_c33;
               Y_16_c34 <= Y_16_c33;
               X_17_c34 <= X_17_c33;
               Y_17_c34 <= Y_17_c33;
               X_18_c34 <= X_18_c33;
               Y_18_c34 <= Y_18_c33;
               X_19_c34 <= X_19_c33;
               Y_19_c34 <= Y_19_c33;
               X_20_c34 <= X_20_c33;
               Y_20_c34 <= Y_20_c33;
               X_21_c34 <= X_21_c33;
               Y_21_c34 <= Y_21_c33;
               X_22_c34 <= X_22_c33;
               Y_22_c34 <= Y_22_c33;
            end if;
            if ce_35 = '1' then
               Cin_1_c35 <= Cin_1_c34;
               X_1_c35 <= X_1_c34;
               Y_1_c35 <= Y_1_c34;
               X_2_c35 <= X_2_c34;
               Y_2_c35 <= Y_2_c34;
               X_3_c35 <= X_3_c34;
               Y_3_c35 <= Y_3_c34;
               X_4_c35 <= X_4_c34;
               Y_4_c35 <= Y_4_c34;
               X_5_c35 <= X_5_c34;
               Y_5_c35 <= Y_5_c34;
               X_6_c35 <= X_6_c34;
               Y_6_c35 <= Y_6_c34;
               X_7_c35 <= X_7_c34;
               Y_7_c35 <= Y_7_c34;
               X_8_c35 <= X_8_c34;
               Y_8_c35 <= Y_8_c34;
               X_9_c35 <= X_9_c34;
               Y_9_c35 <= Y_9_c34;
               X_10_c35 <= X_10_c34;
               Y_10_c35 <= Y_10_c34;
               X_11_c35 <= X_11_c34;
               Y_11_c35 <= Y_11_c34;
               X_12_c35 <= X_12_c34;
               Y_12_c35 <= Y_12_c34;
               X_13_c35 <= X_13_c34;
               Y_13_c35 <= Y_13_c34;
               X_14_c35 <= X_14_c34;
               Y_14_c35 <= Y_14_c34;
               X_15_c35 <= X_15_c34;
               Y_15_c35 <= Y_15_c34;
               X_16_c35 <= X_16_c34;
               Y_16_c35 <= Y_16_c34;
               X_17_c35 <= X_17_c34;
               Y_17_c35 <= Y_17_c34;
               X_18_c35 <= X_18_c34;
               Y_18_c35 <= Y_18_c34;
               X_19_c35 <= X_19_c34;
               Y_19_c35 <= Y_19_c34;
               X_20_c35 <= X_20_c34;
               Y_20_c35 <= Y_20_c34;
               X_21_c35 <= X_21_c34;
               Y_21_c35 <= Y_21_c34;
               X_22_c35 <= X_22_c34;
               Y_22_c35 <= Y_22_c34;
            end if;
            if ce_36 = '1' then
               R_1_c36 <= R_1_c35;
               Cin_2_c36 <= Cin_2_c35;
               X_2_c36 <= X_2_c35;
               Y_2_c36 <= Y_2_c35;
               X_3_c36 <= X_3_c35;
               Y_3_c36 <= Y_3_c35;
               X_4_c36 <= X_4_c35;
               Y_4_c36 <= Y_4_c35;
               X_5_c36 <= X_5_c35;
               Y_5_c36 <= Y_5_c35;
               X_6_c36 <= X_6_c35;
               Y_6_c36 <= Y_6_c35;
               X_7_c36 <= X_7_c35;
               Y_7_c36 <= Y_7_c35;
               X_8_c36 <= X_8_c35;
               Y_8_c36 <= Y_8_c35;
               X_9_c36 <= X_9_c35;
               Y_9_c36 <= Y_9_c35;
               X_10_c36 <= X_10_c35;
               Y_10_c36 <= Y_10_c35;
               X_11_c36 <= X_11_c35;
               Y_11_c36 <= Y_11_c35;
               X_12_c36 <= X_12_c35;
               Y_12_c36 <= Y_12_c35;
               X_13_c36 <= X_13_c35;
               Y_13_c36 <= Y_13_c35;
               X_14_c36 <= X_14_c35;
               Y_14_c36 <= Y_14_c35;
               X_15_c36 <= X_15_c35;
               Y_15_c36 <= Y_15_c35;
               X_16_c36 <= X_16_c35;
               Y_16_c36 <= Y_16_c35;
               X_17_c36 <= X_17_c35;
               Y_17_c36 <= Y_17_c35;
               X_18_c36 <= X_18_c35;
               Y_18_c36 <= Y_18_c35;
               X_19_c36 <= X_19_c35;
               Y_19_c36 <= Y_19_c35;
               X_20_c36 <= X_20_c35;
               Y_20_c36 <= Y_20_c35;
               X_21_c36 <= X_21_c35;
               Y_21_c36 <= Y_21_c35;
               X_22_c36 <= X_22_c35;
               Y_22_c36 <= Y_22_c35;
            end if;
            if ce_37 = '1' then
               R_1_c37 <= R_1_c36;
               R_2_c37 <= R_2_c36;
               Cin_3_c37 <= Cin_3_c36;
               X_3_c37 <= X_3_c36;
               Y_3_c37 <= Y_3_c36;
               X_4_c37 <= X_4_c36;
               Y_4_c37 <= Y_4_c36;
               X_5_c37 <= X_5_c36;
               Y_5_c37 <= Y_5_c36;
               X_6_c37 <= X_6_c36;
               Y_6_c37 <= Y_6_c36;
               X_7_c37 <= X_7_c36;
               Y_7_c37 <= Y_7_c36;
               X_8_c37 <= X_8_c36;
               Y_8_c37 <= Y_8_c36;
               X_9_c37 <= X_9_c36;
               Y_9_c37 <= Y_9_c36;
               X_10_c37 <= X_10_c36;
               Y_10_c37 <= Y_10_c36;
               X_11_c37 <= X_11_c36;
               Y_11_c37 <= Y_11_c36;
               X_12_c37 <= X_12_c36;
               Y_12_c37 <= Y_12_c36;
               X_13_c37 <= X_13_c36;
               Y_13_c37 <= Y_13_c36;
               X_14_c37 <= X_14_c36;
               Y_14_c37 <= Y_14_c36;
               X_15_c37 <= X_15_c36;
               Y_15_c37 <= Y_15_c36;
               X_16_c37 <= X_16_c36;
               Y_16_c37 <= Y_16_c36;
               X_17_c37 <= X_17_c36;
               Y_17_c37 <= Y_17_c36;
               X_18_c37 <= X_18_c36;
               Y_18_c37 <= Y_18_c36;
               X_19_c37 <= X_19_c36;
               Y_19_c37 <= Y_19_c36;
               X_20_c37 <= X_20_c36;
               Y_20_c37 <= Y_20_c36;
               X_21_c37 <= X_21_c36;
               Y_21_c37 <= Y_21_c36;
               X_22_c37 <= X_22_c36;
               Y_22_c37 <= Y_22_c36;
            end if;
            if ce_38 = '1' then
               R_1_c38 <= R_1_c37;
               R_2_c38 <= R_2_c37;
               R_3_c38 <= R_3_c37;
               Cin_4_c38 <= Cin_4_c37;
               X_4_c38 <= X_4_c37;
               Y_4_c38 <= Y_4_c37;
               X_5_c38 <= X_5_c37;
               Y_5_c38 <= Y_5_c37;
               X_6_c38 <= X_6_c37;
               Y_6_c38 <= Y_6_c37;
               X_7_c38 <= X_7_c37;
               Y_7_c38 <= Y_7_c37;
               X_8_c38 <= X_8_c37;
               Y_8_c38 <= Y_8_c37;
               X_9_c38 <= X_9_c37;
               Y_9_c38 <= Y_9_c37;
               X_10_c38 <= X_10_c37;
               Y_10_c38 <= Y_10_c37;
               X_11_c38 <= X_11_c37;
               Y_11_c38 <= Y_11_c37;
               X_12_c38 <= X_12_c37;
               Y_12_c38 <= Y_12_c37;
               X_13_c38 <= X_13_c37;
               Y_13_c38 <= Y_13_c37;
               X_14_c38 <= X_14_c37;
               Y_14_c38 <= Y_14_c37;
               X_15_c38 <= X_15_c37;
               Y_15_c38 <= Y_15_c37;
               X_16_c38 <= X_16_c37;
               Y_16_c38 <= Y_16_c37;
               X_17_c38 <= X_17_c37;
               Y_17_c38 <= Y_17_c37;
               X_18_c38 <= X_18_c37;
               Y_18_c38 <= Y_18_c37;
               X_19_c38 <= X_19_c37;
               Y_19_c38 <= Y_19_c37;
               X_20_c38 <= X_20_c37;
               Y_20_c38 <= Y_20_c37;
               X_21_c38 <= X_21_c37;
               Y_21_c38 <= Y_21_c37;
               X_22_c38 <= X_22_c37;
               Y_22_c38 <= Y_22_c37;
            end if;
            if ce_39 = '1' then
               R_1_c39 <= R_1_c38;
               R_2_c39 <= R_2_c38;
               R_3_c39 <= R_3_c38;
               R_4_c39 <= R_4_c38;
               Cin_5_c39 <= Cin_5_c38;
               X_5_c39 <= X_5_c38;
               Y_5_c39 <= Y_5_c38;
               X_6_c39 <= X_6_c38;
               Y_6_c39 <= Y_6_c38;
               X_7_c39 <= X_7_c38;
               Y_7_c39 <= Y_7_c38;
               X_8_c39 <= X_8_c38;
               Y_8_c39 <= Y_8_c38;
               X_9_c39 <= X_9_c38;
               Y_9_c39 <= Y_9_c38;
               X_10_c39 <= X_10_c38;
               Y_10_c39 <= Y_10_c38;
               X_11_c39 <= X_11_c38;
               Y_11_c39 <= Y_11_c38;
               X_12_c39 <= X_12_c38;
               Y_12_c39 <= Y_12_c38;
               X_13_c39 <= X_13_c38;
               Y_13_c39 <= Y_13_c38;
               X_14_c39 <= X_14_c38;
               Y_14_c39 <= Y_14_c38;
               X_15_c39 <= X_15_c38;
               Y_15_c39 <= Y_15_c38;
               X_16_c39 <= X_16_c38;
               Y_16_c39 <= Y_16_c38;
               X_17_c39 <= X_17_c38;
               Y_17_c39 <= Y_17_c38;
               X_18_c39 <= X_18_c38;
               Y_18_c39 <= Y_18_c38;
               X_19_c39 <= X_19_c38;
               Y_19_c39 <= Y_19_c38;
               X_20_c39 <= X_20_c38;
               Y_20_c39 <= Y_20_c38;
               X_21_c39 <= X_21_c38;
               Y_21_c39 <= Y_21_c38;
               X_22_c39 <= X_22_c38;
               Y_22_c39 <= Y_22_c38;
            end if;
            if ce_40 = '1' then
               R_1_c40 <= R_1_c39;
               R_2_c40 <= R_2_c39;
               R_3_c40 <= R_3_c39;
               R_4_c40 <= R_4_c39;
               R_5_c40 <= R_5_c39;
               Cin_6_c40 <= Cin_6_c39;
               X_6_c40 <= X_6_c39;
               Y_6_c40 <= Y_6_c39;
               X_7_c40 <= X_7_c39;
               Y_7_c40 <= Y_7_c39;
               X_8_c40 <= X_8_c39;
               Y_8_c40 <= Y_8_c39;
               X_9_c40 <= X_9_c39;
               Y_9_c40 <= Y_9_c39;
               X_10_c40 <= X_10_c39;
               Y_10_c40 <= Y_10_c39;
               X_11_c40 <= X_11_c39;
               Y_11_c40 <= Y_11_c39;
               X_12_c40 <= X_12_c39;
               Y_12_c40 <= Y_12_c39;
               X_13_c40 <= X_13_c39;
               Y_13_c40 <= Y_13_c39;
               X_14_c40 <= X_14_c39;
               Y_14_c40 <= Y_14_c39;
               X_15_c40 <= X_15_c39;
               Y_15_c40 <= Y_15_c39;
               X_16_c40 <= X_16_c39;
               Y_16_c40 <= Y_16_c39;
               X_17_c40 <= X_17_c39;
               Y_17_c40 <= Y_17_c39;
               X_18_c40 <= X_18_c39;
               Y_18_c40 <= Y_18_c39;
               X_19_c40 <= X_19_c39;
               Y_19_c40 <= Y_19_c39;
               X_20_c40 <= X_20_c39;
               Y_20_c40 <= Y_20_c39;
               X_21_c40 <= X_21_c39;
               Y_21_c40 <= Y_21_c39;
               X_22_c40 <= X_22_c39;
               Y_22_c40 <= Y_22_c39;
            end if;
            if ce_41 = '1' then
               R_1_c41 <= R_1_c40;
               R_2_c41 <= R_2_c40;
               R_3_c41 <= R_3_c40;
               R_4_c41 <= R_4_c40;
               R_5_c41 <= R_5_c40;
               R_6_c41 <= R_6_c40;
               Cin_7_c41 <= Cin_7_c40;
               X_7_c41 <= X_7_c40;
               Y_7_c41 <= Y_7_c40;
               X_8_c41 <= X_8_c40;
               Y_8_c41 <= Y_8_c40;
               X_9_c41 <= X_9_c40;
               Y_9_c41 <= Y_9_c40;
               X_10_c41 <= X_10_c40;
               Y_10_c41 <= Y_10_c40;
               X_11_c41 <= X_11_c40;
               Y_11_c41 <= Y_11_c40;
               X_12_c41 <= X_12_c40;
               Y_12_c41 <= Y_12_c40;
               X_13_c41 <= X_13_c40;
               Y_13_c41 <= Y_13_c40;
               X_14_c41 <= X_14_c40;
               Y_14_c41 <= Y_14_c40;
               X_15_c41 <= X_15_c40;
               Y_15_c41 <= Y_15_c40;
               X_16_c41 <= X_16_c40;
               Y_16_c41 <= Y_16_c40;
               X_17_c41 <= X_17_c40;
               Y_17_c41 <= Y_17_c40;
               X_18_c41 <= X_18_c40;
               Y_18_c41 <= Y_18_c40;
               X_19_c41 <= X_19_c40;
               Y_19_c41 <= Y_19_c40;
               X_20_c41 <= X_20_c40;
               Y_20_c41 <= Y_20_c40;
               X_21_c41 <= X_21_c40;
               Y_21_c41 <= Y_21_c40;
               X_22_c41 <= X_22_c40;
               Y_22_c41 <= Y_22_c40;
            end if;
            if ce_42 = '1' then
               R_1_c42 <= R_1_c41;
               R_2_c42 <= R_2_c41;
               R_3_c42 <= R_3_c41;
               R_4_c42 <= R_4_c41;
               R_5_c42 <= R_5_c41;
               R_6_c42 <= R_6_c41;
               R_7_c42 <= R_7_c41;
               Cin_8_c42 <= Cin_8_c41;
               X_8_c42 <= X_8_c41;
               Y_8_c42 <= Y_8_c41;
               X_9_c42 <= X_9_c41;
               Y_9_c42 <= Y_9_c41;
               X_10_c42 <= X_10_c41;
               Y_10_c42 <= Y_10_c41;
               X_11_c42 <= X_11_c41;
               Y_11_c42 <= Y_11_c41;
               X_12_c42 <= X_12_c41;
               Y_12_c42 <= Y_12_c41;
               X_13_c42 <= X_13_c41;
               Y_13_c42 <= Y_13_c41;
               X_14_c42 <= X_14_c41;
               Y_14_c42 <= Y_14_c41;
               X_15_c42 <= X_15_c41;
               Y_15_c42 <= Y_15_c41;
               X_16_c42 <= X_16_c41;
               Y_16_c42 <= Y_16_c41;
               X_17_c42 <= X_17_c41;
               Y_17_c42 <= Y_17_c41;
               X_18_c42 <= X_18_c41;
               Y_18_c42 <= Y_18_c41;
               X_19_c42 <= X_19_c41;
               Y_19_c42 <= Y_19_c41;
               X_20_c42 <= X_20_c41;
               Y_20_c42 <= Y_20_c41;
               X_21_c42 <= X_21_c41;
               Y_21_c42 <= Y_21_c41;
               X_22_c42 <= X_22_c41;
               Y_22_c42 <= Y_22_c41;
            end if;
            if ce_43 = '1' then
               R_1_c43 <= R_1_c42;
               R_2_c43 <= R_2_c42;
               R_3_c43 <= R_3_c42;
               R_4_c43 <= R_4_c42;
               R_5_c43 <= R_5_c42;
               R_6_c43 <= R_6_c42;
               R_7_c43 <= R_7_c42;
               R_8_c43 <= R_8_c42;
               Cin_9_c43 <= Cin_9_c42;
               X_9_c43 <= X_9_c42;
               Y_9_c43 <= Y_9_c42;
               X_10_c43 <= X_10_c42;
               Y_10_c43 <= Y_10_c42;
               X_11_c43 <= X_11_c42;
               Y_11_c43 <= Y_11_c42;
               X_12_c43 <= X_12_c42;
               Y_12_c43 <= Y_12_c42;
               X_13_c43 <= X_13_c42;
               Y_13_c43 <= Y_13_c42;
               X_14_c43 <= X_14_c42;
               Y_14_c43 <= Y_14_c42;
               X_15_c43 <= X_15_c42;
               Y_15_c43 <= Y_15_c42;
               X_16_c43 <= X_16_c42;
               Y_16_c43 <= Y_16_c42;
               X_17_c43 <= X_17_c42;
               Y_17_c43 <= Y_17_c42;
               X_18_c43 <= X_18_c42;
               Y_18_c43 <= Y_18_c42;
               X_19_c43 <= X_19_c42;
               Y_19_c43 <= Y_19_c42;
               X_20_c43 <= X_20_c42;
               Y_20_c43 <= Y_20_c42;
               X_21_c43 <= X_21_c42;
               Y_21_c43 <= Y_21_c42;
               X_22_c43 <= X_22_c42;
               Y_22_c43 <= Y_22_c42;
            end if;
            if ce_44 = '1' then
               R_1_c44 <= R_1_c43;
               R_2_c44 <= R_2_c43;
               R_3_c44 <= R_3_c43;
               R_4_c44 <= R_4_c43;
               R_5_c44 <= R_5_c43;
               R_6_c44 <= R_6_c43;
               R_7_c44 <= R_7_c43;
               R_8_c44 <= R_8_c43;
               R_9_c44 <= R_9_c43;
               Cin_10_c44 <= Cin_10_c43;
               X_10_c44 <= X_10_c43;
               Y_10_c44 <= Y_10_c43;
               X_11_c44 <= X_11_c43;
               Y_11_c44 <= Y_11_c43;
               X_12_c44 <= X_12_c43;
               Y_12_c44 <= Y_12_c43;
               X_13_c44 <= X_13_c43;
               Y_13_c44 <= Y_13_c43;
               X_14_c44 <= X_14_c43;
               Y_14_c44 <= Y_14_c43;
               X_15_c44 <= X_15_c43;
               Y_15_c44 <= Y_15_c43;
               X_16_c44 <= X_16_c43;
               Y_16_c44 <= Y_16_c43;
               X_17_c44 <= X_17_c43;
               Y_17_c44 <= Y_17_c43;
               X_18_c44 <= X_18_c43;
               Y_18_c44 <= Y_18_c43;
               X_19_c44 <= X_19_c43;
               Y_19_c44 <= Y_19_c43;
               X_20_c44 <= X_20_c43;
               Y_20_c44 <= Y_20_c43;
               X_21_c44 <= X_21_c43;
               Y_21_c44 <= Y_21_c43;
               X_22_c44 <= X_22_c43;
               Y_22_c44 <= Y_22_c43;
            end if;
            if ce_45 = '1' then
               R_1_c45 <= R_1_c44;
               R_2_c45 <= R_2_c44;
               R_3_c45 <= R_3_c44;
               R_4_c45 <= R_4_c44;
               R_5_c45 <= R_5_c44;
               R_6_c45 <= R_6_c44;
               R_7_c45 <= R_7_c44;
               R_8_c45 <= R_8_c44;
               R_9_c45 <= R_9_c44;
               R_10_c45 <= R_10_c44;
               Cin_11_c45 <= Cin_11_c44;
               X_11_c45 <= X_11_c44;
               Y_11_c45 <= Y_11_c44;
               X_12_c45 <= X_12_c44;
               Y_12_c45 <= Y_12_c44;
               X_13_c45 <= X_13_c44;
               Y_13_c45 <= Y_13_c44;
               X_14_c45 <= X_14_c44;
               Y_14_c45 <= Y_14_c44;
               X_15_c45 <= X_15_c44;
               Y_15_c45 <= Y_15_c44;
               X_16_c45 <= X_16_c44;
               Y_16_c45 <= Y_16_c44;
               X_17_c45 <= X_17_c44;
               Y_17_c45 <= Y_17_c44;
               X_18_c45 <= X_18_c44;
               Y_18_c45 <= Y_18_c44;
               X_19_c45 <= X_19_c44;
               Y_19_c45 <= Y_19_c44;
               X_20_c45 <= X_20_c44;
               Y_20_c45 <= Y_20_c44;
               X_21_c45 <= X_21_c44;
               Y_21_c45 <= Y_21_c44;
               X_22_c45 <= X_22_c44;
               Y_22_c45 <= Y_22_c44;
            end if;
            if ce_46 = '1' then
               R_1_c46 <= R_1_c45;
               R_2_c46 <= R_2_c45;
               R_3_c46 <= R_3_c45;
               R_4_c46 <= R_4_c45;
               R_5_c46 <= R_5_c45;
               R_6_c46 <= R_6_c45;
               R_7_c46 <= R_7_c45;
               R_8_c46 <= R_8_c45;
               R_9_c46 <= R_9_c45;
               R_10_c46 <= R_10_c45;
               R_11_c46 <= R_11_c45;
               Cin_12_c46 <= Cin_12_c45;
               X_12_c46 <= X_12_c45;
               Y_12_c46 <= Y_12_c45;
               X_13_c46 <= X_13_c45;
               Y_13_c46 <= Y_13_c45;
               X_14_c46 <= X_14_c45;
               Y_14_c46 <= Y_14_c45;
               X_15_c46 <= X_15_c45;
               Y_15_c46 <= Y_15_c45;
               X_16_c46 <= X_16_c45;
               Y_16_c46 <= Y_16_c45;
               X_17_c46 <= X_17_c45;
               Y_17_c46 <= Y_17_c45;
               X_18_c46 <= X_18_c45;
               Y_18_c46 <= Y_18_c45;
               X_19_c46 <= X_19_c45;
               Y_19_c46 <= Y_19_c45;
               X_20_c46 <= X_20_c45;
               Y_20_c46 <= Y_20_c45;
               X_21_c46 <= X_21_c45;
               Y_21_c46 <= Y_21_c45;
               X_22_c46 <= X_22_c45;
               Y_22_c46 <= Y_22_c45;
            end if;
            if ce_47 = '1' then
               R_1_c47 <= R_1_c46;
               R_2_c47 <= R_2_c46;
               R_3_c47 <= R_3_c46;
               R_4_c47 <= R_4_c46;
               R_5_c47 <= R_5_c46;
               R_6_c47 <= R_6_c46;
               R_7_c47 <= R_7_c46;
               R_8_c47 <= R_8_c46;
               R_9_c47 <= R_9_c46;
               R_10_c47 <= R_10_c46;
               R_11_c47 <= R_11_c46;
               R_12_c47 <= R_12_c46;
               Cin_13_c47 <= Cin_13_c46;
               X_13_c47 <= X_13_c46;
               Y_13_c47 <= Y_13_c46;
               X_14_c47 <= X_14_c46;
               Y_14_c47 <= Y_14_c46;
               X_15_c47 <= X_15_c46;
               Y_15_c47 <= Y_15_c46;
               X_16_c47 <= X_16_c46;
               Y_16_c47 <= Y_16_c46;
               X_17_c47 <= X_17_c46;
               Y_17_c47 <= Y_17_c46;
               X_18_c47 <= X_18_c46;
               Y_18_c47 <= Y_18_c46;
               X_19_c47 <= X_19_c46;
               Y_19_c47 <= Y_19_c46;
               X_20_c47 <= X_20_c46;
               Y_20_c47 <= Y_20_c46;
               X_21_c47 <= X_21_c46;
               Y_21_c47 <= Y_21_c46;
               X_22_c47 <= X_22_c46;
               Y_22_c47 <= Y_22_c46;
            end if;
            if ce_48 = '1' then
               R_1_c48 <= R_1_c47;
               R_2_c48 <= R_2_c47;
               R_3_c48 <= R_3_c47;
               R_4_c48 <= R_4_c47;
               R_5_c48 <= R_5_c47;
               R_6_c48 <= R_6_c47;
               R_7_c48 <= R_7_c47;
               R_8_c48 <= R_8_c47;
               R_9_c48 <= R_9_c47;
               R_10_c48 <= R_10_c47;
               R_11_c48 <= R_11_c47;
               R_12_c48 <= R_12_c47;
               R_13_c48 <= R_13_c47;
               Cin_14_c48 <= Cin_14_c47;
               X_14_c48 <= X_14_c47;
               Y_14_c48 <= Y_14_c47;
               X_15_c48 <= X_15_c47;
               Y_15_c48 <= Y_15_c47;
               X_16_c48 <= X_16_c47;
               Y_16_c48 <= Y_16_c47;
               X_17_c48 <= X_17_c47;
               Y_17_c48 <= Y_17_c47;
               X_18_c48 <= X_18_c47;
               Y_18_c48 <= Y_18_c47;
               X_19_c48 <= X_19_c47;
               Y_19_c48 <= Y_19_c47;
               X_20_c48 <= X_20_c47;
               Y_20_c48 <= Y_20_c47;
               X_21_c48 <= X_21_c47;
               Y_21_c48 <= Y_21_c47;
               X_22_c48 <= X_22_c47;
               Y_22_c48 <= Y_22_c47;
            end if;
            if ce_49 = '1' then
               R_1_c49 <= R_1_c48;
               R_2_c49 <= R_2_c48;
               R_3_c49 <= R_3_c48;
               R_4_c49 <= R_4_c48;
               R_5_c49 <= R_5_c48;
               R_6_c49 <= R_6_c48;
               R_7_c49 <= R_7_c48;
               R_8_c49 <= R_8_c48;
               R_9_c49 <= R_9_c48;
               R_10_c49 <= R_10_c48;
               R_11_c49 <= R_11_c48;
               R_12_c49 <= R_12_c48;
               R_13_c49 <= R_13_c48;
               R_14_c49 <= R_14_c48;
               Cin_15_c49 <= Cin_15_c48;
               X_15_c49 <= X_15_c48;
               Y_15_c49 <= Y_15_c48;
               X_16_c49 <= X_16_c48;
               Y_16_c49 <= Y_16_c48;
               X_17_c49 <= X_17_c48;
               Y_17_c49 <= Y_17_c48;
               X_18_c49 <= X_18_c48;
               Y_18_c49 <= Y_18_c48;
               X_19_c49 <= X_19_c48;
               Y_19_c49 <= Y_19_c48;
               X_20_c49 <= X_20_c48;
               Y_20_c49 <= Y_20_c48;
               X_21_c49 <= X_21_c48;
               Y_21_c49 <= Y_21_c48;
               X_22_c49 <= X_22_c48;
               Y_22_c49 <= Y_22_c48;
            end if;
            if ce_50 = '1' then
               R_1_c50 <= R_1_c49;
               R_2_c50 <= R_2_c49;
               R_3_c50 <= R_3_c49;
               R_4_c50 <= R_4_c49;
               R_5_c50 <= R_5_c49;
               R_6_c50 <= R_6_c49;
               R_7_c50 <= R_7_c49;
               R_8_c50 <= R_8_c49;
               R_9_c50 <= R_9_c49;
               R_10_c50 <= R_10_c49;
               R_11_c50 <= R_11_c49;
               R_12_c50 <= R_12_c49;
               R_13_c50 <= R_13_c49;
               R_14_c50 <= R_14_c49;
               R_15_c50 <= R_15_c49;
               Cin_16_c50 <= Cin_16_c49;
               X_16_c50 <= X_16_c49;
               Y_16_c50 <= Y_16_c49;
               X_17_c50 <= X_17_c49;
               Y_17_c50 <= Y_17_c49;
               X_18_c50 <= X_18_c49;
               Y_18_c50 <= Y_18_c49;
               X_19_c50 <= X_19_c49;
               Y_19_c50 <= Y_19_c49;
               X_20_c50 <= X_20_c49;
               Y_20_c50 <= Y_20_c49;
               X_21_c50 <= X_21_c49;
               Y_21_c50 <= Y_21_c49;
               X_22_c50 <= X_22_c49;
               Y_22_c50 <= Y_22_c49;
            end if;
            if ce_51 = '1' then
               R_1_c51 <= R_1_c50;
               R_2_c51 <= R_2_c50;
               R_3_c51 <= R_3_c50;
               R_4_c51 <= R_4_c50;
               R_5_c51 <= R_5_c50;
               R_6_c51 <= R_6_c50;
               R_7_c51 <= R_7_c50;
               R_8_c51 <= R_8_c50;
               R_9_c51 <= R_9_c50;
               R_10_c51 <= R_10_c50;
               R_11_c51 <= R_11_c50;
               R_12_c51 <= R_12_c50;
               R_13_c51 <= R_13_c50;
               R_14_c51 <= R_14_c50;
               R_15_c51 <= R_15_c50;
               R_16_c51 <= R_16_c50;
               Cin_17_c51 <= Cin_17_c50;
               X_17_c51 <= X_17_c50;
               Y_17_c51 <= Y_17_c50;
               X_18_c51 <= X_18_c50;
               Y_18_c51 <= Y_18_c50;
               X_19_c51 <= X_19_c50;
               Y_19_c51 <= Y_19_c50;
               X_20_c51 <= X_20_c50;
               Y_20_c51 <= Y_20_c50;
               X_21_c51 <= X_21_c50;
               Y_21_c51 <= Y_21_c50;
               X_22_c51 <= X_22_c50;
               Y_22_c51 <= Y_22_c50;
            end if;
            if ce_52 = '1' then
               R_1_c52 <= R_1_c51;
               R_2_c52 <= R_2_c51;
               R_3_c52 <= R_3_c51;
               R_4_c52 <= R_4_c51;
               R_5_c52 <= R_5_c51;
               R_6_c52 <= R_6_c51;
               R_7_c52 <= R_7_c51;
               R_8_c52 <= R_8_c51;
               R_9_c52 <= R_9_c51;
               R_10_c52 <= R_10_c51;
               R_11_c52 <= R_11_c51;
               R_12_c52 <= R_12_c51;
               R_13_c52 <= R_13_c51;
               R_14_c52 <= R_14_c51;
               R_15_c52 <= R_15_c51;
               R_16_c52 <= R_16_c51;
               R_17_c52 <= R_17_c51;
               Cin_18_c52 <= Cin_18_c51;
               X_18_c52 <= X_18_c51;
               Y_18_c52 <= Y_18_c51;
               X_19_c52 <= X_19_c51;
               Y_19_c52 <= Y_19_c51;
               X_20_c52 <= X_20_c51;
               Y_20_c52 <= Y_20_c51;
               X_21_c52 <= X_21_c51;
               Y_21_c52 <= Y_21_c51;
               X_22_c52 <= X_22_c51;
               Y_22_c52 <= Y_22_c51;
            end if;
            if ce_53 = '1' then
               R_1_c53 <= R_1_c52;
               R_2_c53 <= R_2_c52;
               R_3_c53 <= R_3_c52;
               R_4_c53 <= R_4_c52;
               R_5_c53 <= R_5_c52;
               R_6_c53 <= R_6_c52;
               R_7_c53 <= R_7_c52;
               R_8_c53 <= R_8_c52;
               R_9_c53 <= R_9_c52;
               R_10_c53 <= R_10_c52;
               R_11_c53 <= R_11_c52;
               R_12_c53 <= R_12_c52;
               R_13_c53 <= R_13_c52;
               R_14_c53 <= R_14_c52;
               R_15_c53 <= R_15_c52;
               R_16_c53 <= R_16_c52;
               R_17_c53 <= R_17_c52;
               R_18_c53 <= R_18_c52;
               Cin_19_c53 <= Cin_19_c52;
               X_19_c53 <= X_19_c52;
               Y_19_c53 <= Y_19_c52;
               X_20_c53 <= X_20_c52;
               Y_20_c53 <= Y_20_c52;
               X_21_c53 <= X_21_c52;
               Y_21_c53 <= Y_21_c52;
               X_22_c53 <= X_22_c52;
               Y_22_c53 <= Y_22_c52;
            end if;
            if ce_54 = '1' then
               R_1_c54 <= R_1_c53;
               R_2_c54 <= R_2_c53;
               R_3_c54 <= R_3_c53;
               R_4_c54 <= R_4_c53;
               R_5_c54 <= R_5_c53;
               R_6_c54 <= R_6_c53;
               R_7_c54 <= R_7_c53;
               R_8_c54 <= R_8_c53;
               R_9_c54 <= R_9_c53;
               R_10_c54 <= R_10_c53;
               R_11_c54 <= R_11_c53;
               R_12_c54 <= R_12_c53;
               R_13_c54 <= R_13_c53;
               R_14_c54 <= R_14_c53;
               R_15_c54 <= R_15_c53;
               R_16_c54 <= R_16_c53;
               R_17_c54 <= R_17_c53;
               R_18_c54 <= R_18_c53;
               R_19_c54 <= R_19_c53;
               Cin_20_c54 <= Cin_20_c53;
               X_20_c54 <= X_20_c53;
               Y_20_c54 <= Y_20_c53;
               X_21_c54 <= X_21_c53;
               Y_21_c54 <= Y_21_c53;
               X_22_c54 <= X_22_c53;
               Y_22_c54 <= Y_22_c53;
            end if;
            if ce_55 = '1' then
               R_1_c55 <= R_1_c54;
               R_2_c55 <= R_2_c54;
               R_3_c55 <= R_3_c54;
               R_4_c55 <= R_4_c54;
               R_5_c55 <= R_5_c54;
               R_6_c55 <= R_6_c54;
               R_7_c55 <= R_7_c54;
               R_8_c55 <= R_8_c54;
               R_9_c55 <= R_9_c54;
               R_10_c55 <= R_10_c54;
               R_11_c55 <= R_11_c54;
               R_12_c55 <= R_12_c54;
               R_13_c55 <= R_13_c54;
               R_14_c55 <= R_14_c54;
               R_15_c55 <= R_15_c54;
               R_16_c55 <= R_16_c54;
               R_17_c55 <= R_17_c54;
               R_18_c55 <= R_18_c54;
               R_19_c55 <= R_19_c54;
               R_20_c55 <= R_20_c54;
               Cin_21_c55 <= Cin_21_c54;
               X_21_c55 <= X_21_c54;
               Y_21_c55 <= Y_21_c54;
               X_22_c55 <= X_22_c54;
               Y_22_c55 <= Y_22_c54;
            end if;
            if ce_56 = '1' then
               R_1_c56 <= R_1_c55;
               R_2_c56 <= R_2_c55;
               R_3_c56 <= R_3_c55;
               R_4_c56 <= R_4_c55;
               R_5_c56 <= R_5_c55;
               R_6_c56 <= R_6_c55;
               R_7_c56 <= R_7_c55;
               R_8_c56 <= R_8_c55;
               R_9_c56 <= R_9_c55;
               R_10_c56 <= R_10_c55;
               R_11_c56 <= R_11_c55;
               R_12_c56 <= R_12_c55;
               R_13_c56 <= R_13_c55;
               R_14_c56 <= R_14_c55;
               R_15_c56 <= R_15_c55;
               R_16_c56 <= R_16_c55;
               R_17_c56 <= R_17_c55;
               R_18_c56 <= R_18_c55;
               R_19_c56 <= R_19_c55;
               R_20_c56 <= R_20_c55;
               Cin_21_c56 <= Cin_21_c55;
               X_21_c56 <= X_21_c55;
               Y_21_c56 <= Y_21_c55;
               X_22_c56 <= X_22_c55;
               Y_22_c56 <= Y_22_c55;
            end if;
         end if;
      end process;
   Cin_1_c34 <= Cin;
   X_1_c33 <= '0' & X(2 downto 0);
   Y_1_c0 <= '0' & Y(2 downto 0);
   S_1_c35 <= X_1_c35 + Y_1_c35 + Cin_1_c35;
   R_1_c35 <= S_1_c35(2 downto 0);
   Cin_2_c35 <= S_1_c35(3);
   X_2_c33 <= '0' & X(5 downto 3);
   Y_2_c0 <= '0' & Y(5 downto 3);
   S_2_c36 <= X_2_c36 + Y_2_c36 + Cin_2_c36;
   R_2_c36 <= S_2_c36(2 downto 0);
   Cin_3_c36 <= S_2_c36(3);
   X_3_c33 <= '0' & X(8 downto 6);
   Y_3_c0 <= '0' & Y(8 downto 6);
   S_3_c37 <= X_3_c37 + Y_3_c37 + Cin_3_c37;
   R_3_c37 <= S_3_c37(2 downto 0);
   Cin_4_c37 <= S_3_c37(3);
   X_4_c33 <= '0' & X(11 downto 9);
   Y_4_c0 <= '0' & Y(11 downto 9);
   S_4_c38 <= X_4_c38 + Y_4_c38 + Cin_4_c38;
   R_4_c38 <= S_4_c38(2 downto 0);
   Cin_5_c38 <= S_4_c38(3);
   X_5_c33 <= '0' & X(14 downto 12);
   Y_5_c0 <= '0' & Y(14 downto 12);
   S_5_c39 <= X_5_c39 + Y_5_c39 + Cin_5_c39;
   R_5_c39 <= S_5_c39(2 downto 0);
   Cin_6_c39 <= S_5_c39(3);
   X_6_c33 <= '0' & X(17 downto 15);
   Y_6_c0 <= '0' & Y(17 downto 15);
   S_6_c40 <= X_6_c40 + Y_6_c40 + Cin_6_c40;
   R_6_c40 <= S_6_c40(2 downto 0);
   Cin_7_c40 <= S_6_c40(3);
   X_7_c33 <= '0' & X(20 downto 18);
   Y_7_c0 <= '0' & Y(20 downto 18);
   S_7_c41 <= X_7_c41 + Y_7_c41 + Cin_7_c41;
   R_7_c41 <= S_7_c41(2 downto 0);
   Cin_8_c41 <= S_7_c41(3);
   X_8_c33 <= '0' & X(23 downto 21);
   Y_8_c0 <= '0' & Y(23 downto 21);
   S_8_c42 <= X_8_c42 + Y_8_c42 + Cin_8_c42;
   R_8_c42 <= S_8_c42(2 downto 0);
   Cin_9_c42 <= S_8_c42(3);
   X_9_c33 <= '0' & X(26 downto 24);
   Y_9_c0 <= '0' & Y(26 downto 24);
   S_9_c43 <= X_9_c43 + Y_9_c43 + Cin_9_c43;
   R_9_c43 <= S_9_c43(2 downto 0);
   Cin_10_c43 <= S_9_c43(3);
   X_10_c33 <= '0' & X(29 downto 27);
   Y_10_c0 <= '0' & Y(29 downto 27);
   S_10_c44 <= X_10_c44 + Y_10_c44 + Cin_10_c44;
   R_10_c44 <= S_10_c44(2 downto 0);
   Cin_11_c44 <= S_10_c44(3);
   X_11_c33 <= '0' & X(32 downto 30);
   Y_11_c0 <= '0' & Y(32 downto 30);
   S_11_c45 <= X_11_c45 + Y_11_c45 + Cin_11_c45;
   R_11_c45 <= S_11_c45(2 downto 0);
   Cin_12_c45 <= S_11_c45(3);
   X_12_c33 <= '0' & X(35 downto 33);
   Y_12_c0 <= '0' & Y(35 downto 33);
   S_12_c46 <= X_12_c46 + Y_12_c46 + Cin_12_c46;
   R_12_c46 <= S_12_c46(2 downto 0);
   Cin_13_c46 <= S_12_c46(3);
   X_13_c33 <= '0' & X(38 downto 36);
   Y_13_c0 <= '0' & Y(38 downto 36);
   S_13_c47 <= X_13_c47 + Y_13_c47 + Cin_13_c47;
   R_13_c47 <= S_13_c47(2 downto 0);
   Cin_14_c47 <= S_13_c47(3);
   X_14_c33 <= '0' & X(41 downto 39);
   Y_14_c0 <= '0' & Y(41 downto 39);
   S_14_c48 <= X_14_c48 + Y_14_c48 + Cin_14_c48;
   R_14_c48 <= S_14_c48(2 downto 0);
   Cin_15_c48 <= S_14_c48(3);
   X_15_c33 <= '0' & X(44 downto 42);
   Y_15_c0 <= '0' & Y(44 downto 42);
   S_15_c49 <= X_15_c49 + Y_15_c49 + Cin_15_c49;
   R_15_c49 <= S_15_c49(2 downto 0);
   Cin_16_c49 <= S_15_c49(3);
   X_16_c33 <= '0' & X(47 downto 45);
   Y_16_c0 <= '0' & Y(47 downto 45);
   S_16_c50 <= X_16_c50 + Y_16_c50 + Cin_16_c50;
   R_16_c50 <= S_16_c50(2 downto 0);
   Cin_17_c50 <= S_16_c50(3);
   X_17_c33 <= '0' & X(50 downto 48);
   Y_17_c0 <= '0' & Y(50 downto 48);
   S_17_c51 <= X_17_c51 + Y_17_c51 + Cin_17_c51;
   R_17_c51 <= S_17_c51(2 downto 0);
   Cin_18_c51 <= S_17_c51(3);
   X_18_c33 <= '0' & X(53 downto 51);
   Y_18_c0 <= '0' & Y(53 downto 51);
   S_18_c52 <= X_18_c52 + Y_18_c52 + Cin_18_c52;
   R_18_c52 <= S_18_c52(2 downto 0);
   Cin_19_c52 <= S_18_c52(3);
   X_19_c33 <= '0' & X(56 downto 54);
   Y_19_c0 <= '0' & Y(56 downto 54);
   S_19_c53 <= X_19_c53 + Y_19_c53 + Cin_19_c53;
   R_19_c53 <= S_19_c53(2 downto 0);
   Cin_20_c53 <= S_19_c53(3);
   X_20_c33 <= '0' & X(59 downto 57);
   Y_20_c0 <= '0' & Y(59 downto 57);
   S_20_c54 <= X_20_c54 + Y_20_c54 + Cin_20_c54;
   R_20_c54 <= S_20_c54(2 downto 0);
   Cin_21_c54 <= S_20_c54(3);
   X_21_c33 <= '0' & X(62 downto 60);
   Y_21_c0 <= '0' & Y(62 downto 60);
   S_21_c56 <= X_21_c56 + Y_21_c56 + Cin_21_c56;
   R_21_c56 <= S_21_c56(2 downto 0);
   Cin_22_c56 <= S_21_c56(3);
   X_22_c33 <= '0' & X(64 downto 63);
   Y_22_c0 <= '0' & Y(64 downto 63);
   S_22_c56 <= X_22_c56 + Y_22_c56 + Cin_22_c56;
   R_22_c56 <= S_22_c56(1 downto 0);
   R <= R_22_c56 & R_21_c56 & R_20_c56 & R_19_c56 & R_18_c56 & R_17_c56 & R_16_c56 & R_15_c56 & R_14_c56 & R_13_c56 & R_12_c56 & R_11_c56 & R_10_c56 & R_9_c56 & R_8_c56 & R_7_c56 & R_6_c56 & R_5_c56 & R_4_c56 & R_3_c56 & R_2_c56 & R_1_c56 ;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointMultiplier
--                      (FPMult_11_52_uid2_Freq800_uid3)
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 56 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointMultiplier_64_2_046000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointMultiplier_64_2_046000 is
   component IntMultiplier_53x53_106_Freq800_uid5 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33 : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             Y : in  std_logic_vector(52 downto 0);
             R : out  std_logic_vector(105 downto 0)   );
   end component;

   component IntAdder_65_Freq800_uid975 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56 : in std_logic;
             X : in  std_logic_vector(64 downto 0);
             Y : in  std_logic_vector(64 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(64 downto 0)   );
   end component;

signal sign_c0, sign_c1, sign_c2, sign_c3, sign_c4, sign_c5, sign_c6, sign_c7, sign_c8, sign_c9, sign_c10, sign_c11, sign_c12, sign_c13, sign_c14, sign_c15, sign_c16, sign_c17, sign_c18, sign_c19, sign_c20, sign_c21, sign_c22, sign_c23, sign_c24, sign_c25, sign_c26, sign_c27, sign_c28, sign_c29, sign_c30, sign_c31, sign_c32, sign_c33, sign_c34, sign_c35, sign_c36, sign_c37, sign_c38, sign_c39, sign_c40, sign_c41, sign_c42, sign_c43, sign_c44, sign_c45, sign_c46, sign_c47, sign_c48, sign_c49, sign_c50, sign_c51, sign_c52, sign_c53, sign_c54, sign_c55, sign_c56 :  std_logic;
signal expX_c0, expX_c1 :  std_logic_vector(10 downto 0);
signal expY_c0, expY_c1 :  std_logic_vector(10 downto 0);
signal expSumPreSub_c1, expSumPreSub_c2 :  std_logic_vector(12 downto 0);
signal bias_c0, bias_c1, bias_c2 :  std_logic_vector(12 downto 0);
signal expSum_c2, expSum_c3, expSum_c4, expSum_c5, expSum_c6, expSum_c7, expSum_c8, expSum_c9, expSum_c10, expSum_c11, expSum_c12, expSum_c13, expSum_c14, expSum_c15, expSum_c16, expSum_c17, expSum_c18, expSum_c19, expSum_c20, expSum_c21, expSum_c22, expSum_c23, expSum_c24, expSum_c25, expSum_c26, expSum_c27, expSum_c28, expSum_c29, expSum_c30, expSum_c31, expSum_c32, expSum_c33 :  std_logic_vector(12 downto 0);
signal sigX_c0 :  std_logic_vector(52 downto 0);
signal sigY_c0 :  std_logic_vector(52 downto 0);
signal sigProd_c33 :  std_logic_vector(105 downto 0);
signal excSel_c0 :  std_logic_vector(3 downto 0);
signal exc_c0, exc_c1, exc_c2, exc_c3, exc_c4, exc_c5, exc_c6, exc_c7, exc_c8, exc_c9, exc_c10, exc_c11, exc_c12, exc_c13, exc_c14, exc_c15, exc_c16, exc_c17, exc_c18, exc_c19, exc_c20, exc_c21, exc_c22, exc_c23, exc_c24, exc_c25, exc_c26, exc_c27, exc_c28, exc_c29, exc_c30, exc_c31, exc_c32, exc_c33, exc_c34, exc_c35, exc_c36, exc_c37, exc_c38, exc_c39, exc_c40, exc_c41, exc_c42, exc_c43, exc_c44, exc_c45, exc_c46, exc_c47, exc_c48, exc_c49, exc_c50, exc_c51, exc_c52, exc_c53, exc_c54, exc_c55, exc_c56 :  std_logic_vector(1 downto 0);
signal norm_c33 :  std_logic;
signal expPostNorm_c33 :  std_logic_vector(12 downto 0);
signal sigProdExt_c33, sigProdExt_c34 :  std_logic_vector(105 downto 0);
signal expSig_c33 :  std_logic_vector(64 downto 0);
signal sticky_c33, sticky_c34 :  std_logic;
signal guard_c34 :  std_logic;
signal round_c34 :  std_logic;
signal expSigPostRound_c56 :  std_logic_vector(64 downto 0);
signal excPostNorm_c56 :  std_logic_vector(1 downto 0);
signal finalExc_c56 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               sign_c1 <= sign_c0;
               expX_c1 <= expX_c0;
               expY_c1 <= expY_c0;
               bias_c1 <= bias_c0;
               exc_c1 <= exc_c0;
            end if;
            if ce_2 = '1' then
               sign_c2 <= sign_c1;
               expSumPreSub_c2 <= expSumPreSub_c1;
               bias_c2 <= bias_c1;
               exc_c2 <= exc_c1;
            end if;
            if ce_3 = '1' then
               sign_c3 <= sign_c2;
               expSum_c3 <= expSum_c2;
               exc_c3 <= exc_c2;
            end if;
            if ce_4 = '1' then
               sign_c4 <= sign_c3;
               expSum_c4 <= expSum_c3;
               exc_c4 <= exc_c3;
            end if;
            if ce_5 = '1' then
               sign_c5 <= sign_c4;
               expSum_c5 <= expSum_c4;
               exc_c5 <= exc_c4;
            end if;
            if ce_6 = '1' then
               sign_c6 <= sign_c5;
               expSum_c6 <= expSum_c5;
               exc_c6 <= exc_c5;
            end if;
            if ce_7 = '1' then
               sign_c7 <= sign_c6;
               expSum_c7 <= expSum_c6;
               exc_c7 <= exc_c6;
            end if;
            if ce_8 = '1' then
               sign_c8 <= sign_c7;
               expSum_c8 <= expSum_c7;
               exc_c8 <= exc_c7;
            end if;
            if ce_9 = '1' then
               sign_c9 <= sign_c8;
               expSum_c9 <= expSum_c8;
               exc_c9 <= exc_c8;
            end if;
            if ce_10 = '1' then
               sign_c10 <= sign_c9;
               expSum_c10 <= expSum_c9;
               exc_c10 <= exc_c9;
            end if;
            if ce_11 = '1' then
               sign_c11 <= sign_c10;
               expSum_c11 <= expSum_c10;
               exc_c11 <= exc_c10;
            end if;
            if ce_12 = '1' then
               sign_c12 <= sign_c11;
               expSum_c12 <= expSum_c11;
               exc_c12 <= exc_c11;
            end if;
            if ce_13 = '1' then
               sign_c13 <= sign_c12;
               expSum_c13 <= expSum_c12;
               exc_c13 <= exc_c12;
            end if;
            if ce_14 = '1' then
               sign_c14 <= sign_c13;
               expSum_c14 <= expSum_c13;
               exc_c14 <= exc_c13;
            end if;
            if ce_15 = '1' then
               sign_c15 <= sign_c14;
               expSum_c15 <= expSum_c14;
               exc_c15 <= exc_c14;
            end if;
            if ce_16 = '1' then
               sign_c16 <= sign_c15;
               expSum_c16 <= expSum_c15;
               exc_c16 <= exc_c15;
            end if;
            if ce_17 = '1' then
               sign_c17 <= sign_c16;
               expSum_c17 <= expSum_c16;
               exc_c17 <= exc_c16;
            end if;
            if ce_18 = '1' then
               sign_c18 <= sign_c17;
               expSum_c18 <= expSum_c17;
               exc_c18 <= exc_c17;
            end if;
            if ce_19 = '1' then
               sign_c19 <= sign_c18;
               expSum_c19 <= expSum_c18;
               exc_c19 <= exc_c18;
            end if;
            if ce_20 = '1' then
               sign_c20 <= sign_c19;
               expSum_c20 <= expSum_c19;
               exc_c20 <= exc_c19;
            end if;
            if ce_21 = '1' then
               sign_c21 <= sign_c20;
               expSum_c21 <= expSum_c20;
               exc_c21 <= exc_c20;
            end if;
            if ce_22 = '1' then
               sign_c22 <= sign_c21;
               expSum_c22 <= expSum_c21;
               exc_c22 <= exc_c21;
            end if;
            if ce_23 = '1' then
               sign_c23 <= sign_c22;
               expSum_c23 <= expSum_c22;
               exc_c23 <= exc_c22;
            end if;
            if ce_24 = '1' then
               sign_c24 <= sign_c23;
               expSum_c24 <= expSum_c23;
               exc_c24 <= exc_c23;
            end if;
            if ce_25 = '1' then
               sign_c25 <= sign_c24;
               expSum_c25 <= expSum_c24;
               exc_c25 <= exc_c24;
            end if;
            if ce_26 = '1' then
               sign_c26 <= sign_c25;
               expSum_c26 <= expSum_c25;
               exc_c26 <= exc_c25;
            end if;
            if ce_27 = '1' then
               sign_c27 <= sign_c26;
               expSum_c27 <= expSum_c26;
               exc_c27 <= exc_c26;
            end if;
            if ce_28 = '1' then
               sign_c28 <= sign_c27;
               expSum_c28 <= expSum_c27;
               exc_c28 <= exc_c27;
            end if;
            if ce_29 = '1' then
               sign_c29 <= sign_c28;
               expSum_c29 <= expSum_c28;
               exc_c29 <= exc_c28;
            end if;
            if ce_30 = '1' then
               sign_c30 <= sign_c29;
               expSum_c30 <= expSum_c29;
               exc_c30 <= exc_c29;
            end if;
            if ce_31 = '1' then
               sign_c31 <= sign_c30;
               expSum_c31 <= expSum_c30;
               exc_c31 <= exc_c30;
            end if;
            if ce_32 = '1' then
               sign_c32 <= sign_c31;
               expSum_c32 <= expSum_c31;
               exc_c32 <= exc_c31;
            end if;
            if ce_33 = '1' then
               sign_c33 <= sign_c32;
               expSum_c33 <= expSum_c32;
               exc_c33 <= exc_c32;
            end if;
            if ce_34 = '1' then
               sign_c34 <= sign_c33;
               exc_c34 <= exc_c33;
               sigProdExt_c34 <= sigProdExt_c33;
               sticky_c34 <= sticky_c33;
            end if;
            if ce_35 = '1' then
               sign_c35 <= sign_c34;
               exc_c35 <= exc_c34;
            end if;
            if ce_36 = '1' then
               sign_c36 <= sign_c35;
               exc_c36 <= exc_c35;
            end if;
            if ce_37 = '1' then
               sign_c37 <= sign_c36;
               exc_c37 <= exc_c36;
            end if;
            if ce_38 = '1' then
               sign_c38 <= sign_c37;
               exc_c38 <= exc_c37;
            end if;
            if ce_39 = '1' then
               sign_c39 <= sign_c38;
               exc_c39 <= exc_c38;
            end if;
            if ce_40 = '1' then
               sign_c40 <= sign_c39;
               exc_c40 <= exc_c39;
            end if;
            if ce_41 = '1' then
               sign_c41 <= sign_c40;
               exc_c41 <= exc_c40;
            end if;
            if ce_42 = '1' then
               sign_c42 <= sign_c41;
               exc_c42 <= exc_c41;
            end if;
            if ce_43 = '1' then
               sign_c43 <= sign_c42;
               exc_c43 <= exc_c42;
            end if;
            if ce_44 = '1' then
               sign_c44 <= sign_c43;
               exc_c44 <= exc_c43;
            end if;
            if ce_45 = '1' then
               sign_c45 <= sign_c44;
               exc_c45 <= exc_c44;
            end if;
            if ce_46 = '1' then
               sign_c46 <= sign_c45;
               exc_c46 <= exc_c45;
            end if;
            if ce_47 = '1' then
               sign_c47 <= sign_c46;
               exc_c47 <= exc_c46;
            end if;
            if ce_48 = '1' then
               sign_c48 <= sign_c47;
               exc_c48 <= exc_c47;
            end if;
            if ce_49 = '1' then
               sign_c49 <= sign_c48;
               exc_c49 <= exc_c48;
            end if;
            if ce_50 = '1' then
               sign_c50 <= sign_c49;
               exc_c50 <= exc_c49;
            end if;
            if ce_51 = '1' then
               sign_c51 <= sign_c50;
               exc_c51 <= exc_c50;
            end if;
            if ce_52 = '1' then
               sign_c52 <= sign_c51;
               exc_c52 <= exc_c51;
            end if;
            if ce_53 = '1' then
               sign_c53 <= sign_c52;
               exc_c53 <= exc_c52;
            end if;
            if ce_54 = '1' then
               sign_c54 <= sign_c53;
               exc_c54 <= exc_c53;
            end if;
            if ce_55 = '1' then
               sign_c55 <= sign_c54;
               exc_c55 <= exc_c54;
            end if;
            if ce_56 = '1' then
               sign_c56 <= sign_c55;
               exc_c56 <= exc_c55;
            end if;
         end if;
      end process;
   sign_c0 <= X(63) xor Y(63);
   expX_c0 <= X(62 downto 52);
   expY_c0 <= Y(62 downto 52);
   expSumPreSub_c1 <= ("00" & expX_c1) + ("00" & expY_c1);
   bias_c0 <= CONV_STD_LOGIC_VECTOR(1023,13);
   expSum_c2 <= expSumPreSub_c2 - bias_c2;
   sigX_c0 <= "1" & X(51 downto 0);
   sigY_c0 <= "1" & Y(51 downto 0);
   SignificandMultiplication: IntMultiplier_53x53_106_Freq800_uid5
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 X => sigX_c0,
                 Y => sigY_c0,
                 R => sigProd_c33);
   excSel_c0 <= X(65 downto 64) & Y(65 downto 64);
   with excSel_c0  select  
   exc_c0 <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm_c33 <= sigProd_c33(105);
   -- exponent update
   expPostNorm_c33 <= expSum_c33 + ("000000000000" & norm_c33);
   -- significand normalization shift
   sigProdExt_c33 <= sigProd_c33(104 downto 0) & "0" when norm_c33='1' else
                         sigProd_c33(103 downto 0) & "00";
   expSig_c33 <= expPostNorm_c33 & sigProdExt_c33(105 downto 54);
   sticky_c33 <= sigProdExt_c33(53);
   guard_c34 <= '0' when sigProdExt_c34(52 downto 0)="00000000000000000000000000000000000000000000000000000" else '1';
   round_c34 <= sticky_c34 and ( (guard_c34 and not(sigProdExt_c34(54))) or (sigProdExt_c34(54) ))  ;
   RoundingAdder: IntAdder_65_Freq800_uid975
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 ce_7=> ce_7,
                 ce_8=> ce_8,
                 ce_9=> ce_9,
                 ce_10=> ce_10,
                 ce_11=> ce_11,
                 ce_12=> ce_12,
                 ce_13=> ce_13,
                 ce_14=> ce_14,
                 ce_15=> ce_15,
                 ce_16=> ce_16,
                 ce_17=> ce_17,
                 ce_18=> ce_18,
                 ce_19=> ce_19,
                 ce_20=> ce_20,
                 ce_21=> ce_21,
                 ce_22=> ce_22,
                 ce_23=> ce_23,
                 ce_24=> ce_24,
                 ce_25=> ce_25,
                 ce_26=> ce_26,
                 ce_27=> ce_27,
                 ce_28=> ce_28,
                 ce_29=> ce_29,
                 ce_30=> ce_30,
                 ce_31=> ce_31,
                 ce_32=> ce_32,
                 ce_33=> ce_33,
                 ce_34=> ce_34,
                 ce_35=> ce_35,
                 ce_36=> ce_36,
                 ce_37=> ce_37,
                 ce_38=> ce_38,
                 ce_39=> ce_39,
                 ce_40=> ce_40,
                 ce_41=> ce_41,
                 ce_42=> ce_42,
                 ce_43=> ce_43,
                 ce_44=> ce_44,
                 ce_45=> ce_45,
                 ce_46=> ce_46,
                 ce_47=> ce_47,
                 ce_48=> ce_48,
                 ce_49=> ce_49,
                 ce_50=> ce_50,
                 ce_51=> ce_51,
                 ce_52=> ce_52,
                 ce_53=> ce_53,
                 ce_54=> ce_54,
                 ce_55=> ce_55,
                 ce_56=> ce_56,
                 Cin => round_c34,
                 X => expSig_c33,
                 Y => "00000000000000000000000000000000000000000000000000000000000000000",
                 R => expSigPostRound_c56);
   with expSigPostRound_c56(64 downto 63)  select 
   excPostNorm_c56 <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_c56  select  
   finalExc_c56 <= exc_c56 when  "11"|"10"|"00",
                       excPostNorm_c56 when others; 
   R <= finalExc_c56 & sign_c56 & expSigPostRound_c56(62 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid17
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid17 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid17 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid22
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid22 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid22 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid27
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid27 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid27 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid32
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid32 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid32 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid37
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid37 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid37 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid42
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid42 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid42 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid47
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid47 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid47 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid52
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid52 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid52 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid63
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid63 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid63 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid68
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid68 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid68 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid73
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid73 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid73 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid78
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid78 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid78 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid83
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid83 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid83 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid88
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid88 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid88 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid93
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid93 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid93 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid98
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid98 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid98 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid113
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid113 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid113 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid118
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid118 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid118 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid123
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid128
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid128 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid128 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid133
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid133 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid133 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid138
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid138 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid138 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid143
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid143 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid143 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid148
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid148 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid148 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid153
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid153 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid153 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid158
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid158 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid158 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid163
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid163 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid163 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid168
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid168 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid168 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid183
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid183 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid183 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid188
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid188 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid188 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid193
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid193 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid193 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid198
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid198 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid198 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid203
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid203 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid203 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid208
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid208 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid208 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid213
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid213 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid213 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid218
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid218 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid218 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid223
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid223 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid223 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid228
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid228 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid228 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid233
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid233 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid233 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid238
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid238 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid238 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid253
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid253 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid253 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid258
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid258 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid258 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid263
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid263 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid263 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid268
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid268 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid268 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid273
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid273 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid273 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid278
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid278 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid278 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid283
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid283 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid283 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid288
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid288 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid288 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid293
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid293 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid293 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid298
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid298 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid298 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid303
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid303 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid303 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid308
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid308 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid308 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid313
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid313 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid313 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq500_uid318
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq500_uid318 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq500_uid318 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq500_uid322
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq500_uid322 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq500_uid322 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq500_uid326
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq500_uid326 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq500_uid326 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq500_uid334
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq500_uid334 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq500_uid334 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq500_uid400
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq500_uid400 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq500_uid400 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq500_uid432
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq500_uid432 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq500_uid432 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq500_uid9
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq500_uid9 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq500_uid9 is
signal Mfull_c0, Mfull_c1 :  std_logic_vector(40 downto 0);
signal M_c1 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c1 <= Mfull_c1(40 downto 0);
   R <= M_c1;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq500_uid11
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq500_uid11 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq500_uid11 is
signal Mfull_c0, Mfull_c1 :  std_logic_vector(40 downto 0);
signal M_c1 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c1 <= Mfull_c1(40 downto 0);
   R <= M_c1;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq500_uid13
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq500_uid13 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq500_uid13 is
signal Mfull_c0, Mfull_c1 :  std_logic_vector(40 downto 0);
signal M_c1 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c1 <= Mfull_c1(40 downto 0);
   R <= M_c1;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid15
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid15 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid15 is
   component MultTable_Freq500_uid17 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy18_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid17
      port map ( X => Xtable_c0,
                 Y => Y1_copy18_c0);
   Y1_c0 <= Y1_copy18_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid20
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid20 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid20 is
   component MultTable_Freq500_uid22 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy23_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid22
      port map ( X => Xtable_c0,
                 Y => Y1_copy23_c0);
   Y1_c0 <= Y1_copy23_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid25
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid25 is
   component MultTable_Freq500_uid27 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy28_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid27
      port map ( X => Xtable_c0,
                 Y => Y1_copy28_c0);
   Y1_c0 <= Y1_copy28_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid30
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid30 is
   component MultTable_Freq500_uid32 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy33_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid32
      port map ( X => Xtable_c0,
                 Y => Y1_copy33_c0);
   Y1_c0 <= Y1_copy33_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid35
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid35 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid35 is
   component MultTable_Freq500_uid37 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy38_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid37
      port map ( X => Xtable_c0,
                 Y => Y1_copy38_c0);
   Y1_c0 <= Y1_copy38_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid40
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid40 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid40 is
   component MultTable_Freq500_uid42 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy43_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid42
      port map ( X => Xtable_c0,
                 Y => Y1_copy43_c0);
   Y1_c0 <= Y1_copy43_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid45
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid45 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid45 is
   component MultTable_Freq500_uid47 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy48_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid47
      port map ( X => Xtable_c0,
                 Y => Y1_copy48_c0);
   Y1_c0 <= Y1_copy48_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid50
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid50 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid50 is
   component MultTable_Freq500_uid52 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy53_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid52
      port map ( X => Xtable_c0,
                 Y => Y1_copy53_c0);
   Y1_c0 <= Y1_copy53_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq500_uid55
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq500_uid55 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq500_uid55 is
signal Mfull_c0, Mfull_c1 :  std_logic_vector(40 downto 0);
signal M_c1 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c1 <= Mfull_c1(40 downto 0);
   R <= M_c1;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq500_uid57
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq500_uid57 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq500_uid57 is
signal Mfull_c0, Mfull_c1 :  std_logic_vector(40 downto 0);
signal M_c1 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c1 <= Mfull_c1(40 downto 0);
   R <= M_c1;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq500_uid59
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq500_uid59 is
    port (clk, ce_1 : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq500_uid59 is
signal Mfull_c0, Mfull_c1 :  std_logic_vector(40 downto 0);
signal M_c1 :  std_logic_vector(40 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Mfull_c1 <= Mfull_c0;
            end if;
         end if;
      end process;
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c1 <= Mfull_c1(40 downto 0);
   R <= M_c1;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid61
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid61 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid61 is
   component MultTable_Freq500_uid63 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy64_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid63
      port map ( X => Xtable_c0,
                 Y => Y1_copy64_c0);
   Y1_c0 <= Y1_copy64_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid66
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid66 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid66 is
   component MultTable_Freq500_uid68 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy69_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid68
      port map ( X => Xtable_c0,
                 Y => Y1_copy69_c0);
   Y1_c0 <= Y1_copy69_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid71
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid71 is
   component MultTable_Freq500_uid73 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy74_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid73
      port map ( X => Xtable_c0,
                 Y => Y1_copy74_c0);
   Y1_c0 <= Y1_copy74_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid76
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid76 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid76 is
   component MultTable_Freq500_uid78 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy79_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid78
      port map ( X => Xtable_c0,
                 Y => Y1_copy79_c0);
   Y1_c0 <= Y1_copy79_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid81
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid81 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid81 is
   component MultTable_Freq500_uid83 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy84_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid83
      port map ( X => Xtable_c0,
                 Y => Y1_copy84_c0);
   Y1_c0 <= Y1_copy84_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid86
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid86 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid86 is
   component MultTable_Freq500_uid88 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy89_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid88
      port map ( X => Xtable_c0,
                 Y => Y1_copy89_c0);
   Y1_c0 <= Y1_copy89_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid91
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid91 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid91 is
   component MultTable_Freq500_uid93 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy94_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid93
      port map ( X => Xtable_c0,
                 Y => Y1_copy94_c0);
   Y1_c0 <= Y1_copy94_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq500_uid96
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid96 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid96 is
   component MultTable_Freq500_uid98 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy99_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid98
      port map ( X => Xtable_c0,
                 Y => Y1_copy99_c0);
   Y1_c0 <= Y1_copy99_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq500_uid101
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq500_uid101 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq500_uid101 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid103
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid103 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid103 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid105
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid105 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid105 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid107
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid107 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid107 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid109
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid109 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid109 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq500_uid111
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq500_uid111 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq500_uid111 is
   component MultTable_Freq500_uid113 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy114_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid113
      port map ( X => Xtable_c0,
                 Y => Y1_copy114_c0);
   Y1_c0 <= Y1_copy114_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid116
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid116 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid116 is
   component MultTable_Freq500_uid118 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy119_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid118
      port map ( X => Xtable_c0,
                 Y => Y1_copy119_c0);
   Y1_c0 <= Y1_copy119_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid121
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid121 is
   component MultTable_Freq500_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy124_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid123
      port map ( X => Xtable_c0,
                 Y => Y1_copy124_c0);
   Y1_c0 <= Y1_copy124_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid126
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid126 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid126 is
   component MultTable_Freq500_uid128 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy129_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid128
      port map ( X => Xtable_c0,
                 Y => Y1_copy129_c0);
   Y1_c0 <= Y1_copy129_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid131
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid131 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid131 is
   component MultTable_Freq500_uid133 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy134_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid133
      port map ( X => Xtable_c0,
                 Y => Y1_copy134_c0);
   Y1_c0 <= Y1_copy134_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid136
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid136 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid136 is
   component MultTable_Freq500_uid138 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy139_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid138
      port map ( X => Xtable_c0,
                 Y => Y1_copy139_c0);
   Y1_c0 <= Y1_copy139_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq500_uid141
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq500_uid141 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq500_uid141 is
   component MultTable_Freq500_uid143 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy144_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid143
      port map ( X => Xtable_c0,
                 Y => Y1_copy144_c0);
   Y1_c0 <= Y1_copy144_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid146
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid146 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid146 is
   component MultTable_Freq500_uid148 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy149_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid148
      port map ( X => Xtable_c0,
                 Y => Y1_copy149_c0);
   Y1_c0 <= Y1_copy149_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid151
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid151 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid151 is
   component MultTable_Freq500_uid153 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy154_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid153
      port map ( X => Xtable_c0,
                 Y => Y1_copy154_c0);
   Y1_c0 <= Y1_copy154_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid156
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid156 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid156 is
   component MultTable_Freq500_uid158 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy159_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid158
      port map ( X => Xtable_c0,
                 Y => Y1_copy159_c0);
   Y1_c0 <= Y1_copy159_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid161
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid161 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid161 is
   component MultTable_Freq500_uid163 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy164_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid163
      port map ( X => Xtable_c0,
                 Y => Y1_copy164_c0);
   Y1_c0 <= Y1_copy164_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid166
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid166 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid166 is
   component MultTable_Freq500_uid168 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy169_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid168
      port map ( X => Xtable_c0,
                 Y => Y1_copy169_c0);
   Y1_c0 <= Y1_copy169_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq500_uid171
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq500_uid171 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq500_uid171 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid173
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid173 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid173 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid175
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid175 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid175 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid177
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid177 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid177 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid179
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid179 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid179 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq500_uid181
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq500_uid181 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq500_uid181 is
   component MultTable_Freq500_uid183 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy184_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid183
      port map ( X => Xtable_c0,
                 Y => Y1_copy184_c0);
   Y1_c0 <= Y1_copy184_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid186
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid186 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid186 is
   component MultTable_Freq500_uid188 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy189_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid188
      port map ( X => Xtable_c0,
                 Y => Y1_copy189_c0);
   Y1_c0 <= Y1_copy189_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid191
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid191 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid191 is
   component MultTable_Freq500_uid193 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy194_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid193
      port map ( X => Xtable_c0,
                 Y => Y1_copy194_c0);
   Y1_c0 <= Y1_copy194_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid196
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid196 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid196 is
   component MultTable_Freq500_uid198 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy199_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid198
      port map ( X => Xtable_c0,
                 Y => Y1_copy199_c0);
   Y1_c0 <= Y1_copy199_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid201
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid201 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid201 is
   component MultTable_Freq500_uid203 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy204_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid203
      port map ( X => Xtable_c0,
                 Y => Y1_copy204_c0);
   Y1_c0 <= Y1_copy204_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid206
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid206 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid206 is
   component MultTable_Freq500_uid208 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy209_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid208
      port map ( X => Xtable_c0,
                 Y => Y1_copy209_c0);
   Y1_c0 <= Y1_copy209_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq500_uid211
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq500_uid211 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq500_uid211 is
   component MultTable_Freq500_uid213 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy214_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid213
      port map ( X => Xtable_c0,
                 Y => Y1_copy214_c0);
   Y1_c0 <= Y1_copy214_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid216
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid216 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid216 is
   component MultTable_Freq500_uid218 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy219_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid218
      port map ( X => Xtable_c0,
                 Y => Y1_copy219_c0);
   Y1_c0 <= Y1_copy219_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid221
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid221 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid221 is
   component MultTable_Freq500_uid223 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy224_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid223
      port map ( X => Xtable_c0,
                 Y => Y1_copy224_c0);
   Y1_c0 <= Y1_copy224_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid226
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid226 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid226 is
   component MultTable_Freq500_uid228 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy229_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid228
      port map ( X => Xtable_c0,
                 Y => Y1_copy229_c0);
   Y1_c0 <= Y1_copy229_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid231
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid231 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid231 is
   component MultTable_Freq500_uid233 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy234_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid233
      port map ( X => Xtable_c0,
                 Y => Y1_copy234_c0);
   Y1_c0 <= Y1_copy234_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid236
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid236 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid236 is
   component MultTable_Freq500_uid238 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy239_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid238
      port map ( X => Xtable_c0,
                 Y => Y1_copy239_c0);
   Y1_c0 <= Y1_copy239_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq500_uid241
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq500_uid241 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq500_uid241 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid243
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid243 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid243 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid245
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid245 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid245 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid247
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid247 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid247 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq500_uid249
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq500_uid249 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq500_uid249 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq500_uid251
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq500_uid251 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq500_uid251 is
   component MultTable_Freq500_uid253 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy254_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid253
      port map ( X => Xtable_c0,
                 Y => Y1_copy254_c0);
   Y1_c0 <= Y1_copy254_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid256
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid256 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid256 is
   component MultTable_Freq500_uid258 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy259_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid258
      port map ( X => Xtable_c0,
                 Y => Y1_copy259_c0);
   Y1_c0 <= Y1_copy259_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid261
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid261 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid261 is
   component MultTable_Freq500_uid263 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy264_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid263
      port map ( X => Xtable_c0,
                 Y => Y1_copy264_c0);
   Y1_c0 <= Y1_copy264_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid266
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid266 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid266 is
   component MultTable_Freq500_uid268 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy269_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid268
      port map ( X => Xtable_c0,
                 Y => Y1_copy269_c0);
   Y1_c0 <= Y1_copy269_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid271
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid271 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid271 is
   component MultTable_Freq500_uid273 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy274_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid273
      port map ( X => Xtable_c0,
                 Y => Y1_copy274_c0);
   Y1_c0 <= Y1_copy274_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid276
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid276 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid276 is
   component MultTable_Freq500_uid278 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy279_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid278
      port map ( X => Xtable_c0,
                 Y => Y1_copy279_c0);
   Y1_c0 <= Y1_copy279_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq500_uid281
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq500_uid281 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq500_uid281 is
   component MultTable_Freq500_uid283 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy284_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid283
      port map ( X => Xtable_c0,
                 Y => Y1_copy284_c0);
   Y1_c0 <= Y1_copy284_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid286
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid286 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid286 is
   component MultTable_Freq500_uid288 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy289_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid288
      port map ( X => Xtable_c0,
                 Y => Y1_copy289_c0);
   Y1_c0 <= Y1_copy289_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid291
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid291 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid291 is
   component MultTable_Freq500_uid293 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy294_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid293
      port map ( X => Xtable_c0,
                 Y => Y1_copy294_c0);
   Y1_c0 <= Y1_copy294_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid296
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid296 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid296 is
   component MultTable_Freq500_uid298 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy299_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid298
      port map ( X => Xtable_c0,
                 Y => Y1_copy299_c0);
   Y1_c0 <= Y1_copy299_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid301
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid301 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid301 is
   component MultTable_Freq500_uid303 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy304_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid303
      port map ( X => Xtable_c0,
                 Y => Y1_copy304_c0);
   Y1_c0 <= Y1_copy304_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq500_uid306
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq500_uid306 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq500_uid306 is
   component MultTable_Freq500_uid308 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy309_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid308
      port map ( X => Xtable_c0,
                 Y => Y1_copy309_c0);
   Y1_c0 <= Y1_copy309_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq500_uid311
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq500_uid311 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq500_uid311 is
   component MultTable_Freq500_uid313 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy314_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid313
      port map ( X => Xtable_c0,
                 Y => Y1_copy314_c0);
   Y1_c0 <= Y1_copy314_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x3_Freq500_uid316
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq500_uid316 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq500_uid316 is
   component MultTable_Freq500_uid318 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy319_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq500_uid318
      port map ( X => Xtable_c0,
                 Y => Y1_copy319_c0);
   Y1_c0 <= Y1_copy319_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_84_Freq500_uid930
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_84_Freq500_uid930 is
    port (clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(83 downto 0);
          Y : in  std_logic_vector(83 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(83 downto 0)   );
end entity;

architecture arch of IntAdder_84_Freq500_uid930 is
signal Cin_0_c0, Cin_0_c1, Cin_0_c2, Cin_0_c3 :  std_logic;
signal X_0_c2, X_0_c3 :  std_logic_vector(67 downto 0);
signal Y_0_c2, Y_0_c3 :  std_logic_vector(67 downto 0);
signal S_0_c3 :  std_logic_vector(67 downto 0);
signal R_0_c3, R_0_c4 :  std_logic_vector(66 downto 0);
signal Cin_1_c3, Cin_1_c4 :  std_logic;
signal X_1_c2, X_1_c3, X_1_c4 :  std_logic_vector(17 downto 0);
signal Y_1_c2, Y_1_c3, Y_1_c4 :  std_logic_vector(17 downto 0);
signal S_1_c4 :  std_logic_vector(17 downto 0);
signal R_1_c4 :  std_logic_vector(16 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_0_c1 <= Cin_0_c0;
            end if;
            if ce_2 = '1' then
               Cin_0_c2 <= Cin_0_c1;
            end if;
            if ce_3 = '1' then
               Cin_0_c3 <= Cin_0_c2;
               X_0_c3 <= X_0_c2;
               Y_0_c3 <= Y_0_c2;
               X_1_c3 <= X_1_c2;
               Y_1_c3 <= Y_1_c2;
            end if;
            if ce_4 = '1' then
               R_0_c4 <= R_0_c3;
               Cin_1_c4 <= Cin_1_c3;
               X_1_c4 <= X_1_c3;
               Y_1_c4 <= Y_1_c3;
            end if;
         end if;
      end process;
   Cin_0_c0 <= Cin;
   X_0_c2 <= '0' & X(66 downto 0);
   Y_0_c2 <= '0' & Y(66 downto 0);
   S_0_c3 <= X_0_c3 + Y_0_c3 + Cin_0_c3;
   R_0_c3 <= S_0_c3(66 downto 0);
   Cin_1_c3 <= S_0_c3(67);
   X_1_c2 <= '0' & X(83 downto 67);
   Y_1_c2 <= '0' & Y(83 downto 67);
   S_1_c4 <= X_1_c4 + Y_1_c4 + Cin_1_c4;
   R_1_c4 <= S_1_c4(16 downto 0);
   R <= R_1_c4 & R_0_c4 ;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_53x53_106_Freq500_uid5
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_53x53_106_Freq500_uid5 is
    port (clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          Y : in  std_logic_vector(52 downto 0);
          R : out  std_logic_vector(105 downto 0)   );
end entity;

architecture arch of IntMultiplier_53x53_106_Freq500_uid5 is
   component DSPBlock_17x24_Freq500_uid9 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq500_uid11 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq500_uid13 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid15 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid20 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid35 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid40 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid45 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid50 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq500_uid55 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq500_uid57 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq500_uid59 is
      port ( clk, ce_1 : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid61 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid66 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid76 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid81 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid86 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid91 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid96 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq500_uid101 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid103 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid105 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid107 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid109 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq500_uid111 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid116 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid126 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid131 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid136 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq500_uid141 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid146 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid151 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid156 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid161 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid166 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq500_uid171 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid173 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid175 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid177 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid179 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq500_uid181 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid186 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid191 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid196 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid201 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid206 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq500_uid211 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid216 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid221 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid226 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid231 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid236 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq500_uid241 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid243 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid245 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid247 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq500_uid249 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq500_uid251 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid256 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid261 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid266 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid271 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid276 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq500_uid281 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid286 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid291 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid296 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid301 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq500_uid306 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq500_uid311 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq500_uid316 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq500_uid322 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq500_uid326 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq500_uid334 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq500_uid400 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq500_uid432 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntAdder_84_Freq500_uid930 is
      port ( clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
             X : in  std_logic_vector(83 downto 0);
             Y : in  std_logic_vector(83 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(83 downto 0)   );
   end component;

signal XX_m6_c0 :  std_logic_vector(52 downto 0);
signal YY_m6_c0 :  std_logic_vector(52 downto 0);
signal tile_0_X_c0 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_0_output_c1 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c1 :  unsigned(40-0 downto 0);
signal bh7_w0_0_c1, bh7_w0_0_c2 :  std_logic;
signal bh7_w1_0_c1, bh7_w1_0_c2 :  std_logic;
signal bh7_w2_0_c1, bh7_w2_0_c2 :  std_logic;
signal bh7_w3_0_c1, bh7_w3_0_c2 :  std_logic;
signal bh7_w4_0_c1, bh7_w4_0_c2 :  std_logic;
signal bh7_w5_0_c1, bh7_w5_0_c2 :  std_logic;
signal bh7_w6_0_c1, bh7_w6_0_c2 :  std_logic;
signal bh7_w7_0_c1, bh7_w7_0_c2 :  std_logic;
signal bh7_w8_0_c1, bh7_w8_0_c2 :  std_logic;
signal bh7_w9_0_c1, bh7_w9_0_c2 :  std_logic;
signal bh7_w10_0_c1, bh7_w10_0_c2 :  std_logic;
signal bh7_w11_0_c1, bh7_w11_0_c2 :  std_logic;
signal bh7_w12_0_c1, bh7_w12_0_c2 :  std_logic;
signal bh7_w13_0_c1, bh7_w13_0_c2 :  std_logic;
signal bh7_w14_0_c1, bh7_w14_0_c2 :  std_logic;
signal bh7_w15_0_c1, bh7_w15_0_c2 :  std_logic;
signal bh7_w16_0_c1, bh7_w16_0_c2 :  std_logic;
signal bh7_w17_0_c1 :  std_logic;
signal bh7_w18_0_c1 :  std_logic;
signal bh7_w19_0_c1 :  std_logic;
signal bh7_w20_0_c1 :  std_logic;
signal bh7_w21_0_c1 :  std_logic;
signal bh7_w22_0_c1 :  std_logic;
signal bh7_w23_0_c1 :  std_logic;
signal bh7_w24_0_c1 :  std_logic;
signal bh7_w25_0_c1 :  std_logic;
signal bh7_w26_0_c1 :  std_logic;
signal bh7_w27_0_c1 :  std_logic;
signal bh7_w28_0_c1 :  std_logic;
signal bh7_w29_0_c1 :  std_logic;
signal bh7_w30_0_c1 :  std_logic;
signal bh7_w31_0_c1 :  std_logic;
signal bh7_w32_0_c1 :  std_logic;
signal bh7_w33_0_c1 :  std_logic;
signal bh7_w34_0_c1 :  std_logic;
signal bh7_w35_0_c1 :  std_logic;
signal bh7_w36_0_c1 :  std_logic;
signal bh7_w37_0_c1 :  std_logic;
signal bh7_w38_0_c1 :  std_logic;
signal bh7_w39_0_c1 :  std_logic;
signal bh7_w40_0_c1 :  std_logic;
signal tile_1_X_c0 :  std_logic_vector(16 downto 0);
signal tile_1_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_1_output_c1 :  std_logic_vector(40 downto 0);
signal tile_1_filtered_output_c1 :  unsigned(40-0 downto 0);
signal bh7_w17_1_c1 :  std_logic;
signal bh7_w18_1_c1 :  std_logic;
signal bh7_w19_1_c1 :  std_logic;
signal bh7_w20_1_c1 :  std_logic;
signal bh7_w21_1_c1 :  std_logic;
signal bh7_w22_1_c1 :  std_logic;
signal bh7_w23_1_c1 :  std_logic;
signal bh7_w24_1_c1 :  std_logic;
signal bh7_w25_1_c1 :  std_logic;
signal bh7_w26_1_c1 :  std_logic;
signal bh7_w27_1_c1 :  std_logic;
signal bh7_w28_1_c1 :  std_logic;
signal bh7_w29_1_c1 :  std_logic;
signal bh7_w30_1_c1 :  std_logic;
signal bh7_w31_1_c1 :  std_logic;
signal bh7_w32_1_c1 :  std_logic;
signal bh7_w33_1_c1 :  std_logic;
signal bh7_w34_1_c1 :  std_logic;
signal bh7_w35_1_c1 :  std_logic;
signal bh7_w36_1_c1 :  std_logic;
signal bh7_w37_1_c1 :  std_logic;
signal bh7_w38_1_c1 :  std_logic;
signal bh7_w39_1_c1 :  std_logic;
signal bh7_w40_1_c1 :  std_logic;
signal bh7_w41_0_c1 :  std_logic;
signal bh7_w42_0_c1 :  std_logic;
signal bh7_w43_0_c1 :  std_logic;
signal bh7_w44_0_c1 :  std_logic;
signal bh7_w45_0_c1 :  std_logic;
signal bh7_w46_0_c1 :  std_logic;
signal bh7_w47_0_c1 :  std_logic;
signal bh7_w48_0_c1 :  std_logic;
signal bh7_w49_0_c1 :  std_logic;
signal bh7_w50_0_c1 :  std_logic;
signal bh7_w51_0_c1 :  std_logic;
signal bh7_w52_0_c1 :  std_logic;
signal bh7_w53_0_c1 :  std_logic;
signal bh7_w54_0_c1 :  std_logic;
signal bh7_w55_0_c1 :  std_logic;
signal bh7_w56_0_c1 :  std_logic;
signal bh7_w57_0_c1 :  std_logic;
signal tile_2_X_c0 :  std_logic_vector(16 downto 0);
signal tile_2_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_2_output_c1 :  std_logic_vector(40 downto 0);
signal tile_2_filtered_output_c1 :  unsigned(40-0 downto 0);
signal bh7_w34_2_c1 :  std_logic;
signal bh7_w35_2_c1 :  std_logic;
signal bh7_w36_2_c1 :  std_logic;
signal bh7_w37_2_c1 :  std_logic;
signal bh7_w38_2_c1 :  std_logic;
signal bh7_w39_2_c1 :  std_logic;
signal bh7_w40_2_c1 :  std_logic;
signal bh7_w41_1_c1 :  std_logic;
signal bh7_w42_1_c1 :  std_logic;
signal bh7_w43_1_c1 :  std_logic;
signal bh7_w44_1_c1 :  std_logic;
signal bh7_w45_1_c1 :  std_logic;
signal bh7_w46_1_c1 :  std_logic;
signal bh7_w47_1_c1 :  std_logic;
signal bh7_w48_1_c1 :  std_logic;
signal bh7_w49_1_c1 :  std_logic;
signal bh7_w50_1_c1 :  std_logic;
signal bh7_w51_1_c1 :  std_logic;
signal bh7_w52_1_c1 :  std_logic;
signal bh7_w53_1_c1 :  std_logic;
signal bh7_w54_1_c1 :  std_logic;
signal bh7_w55_1_c1 :  std_logic;
signal bh7_w56_1_c1 :  std_logic;
signal bh7_w57_1_c1 :  std_logic;
signal bh7_w58_0_c1 :  std_logic;
signal bh7_w59_0_c1 :  std_logic;
signal bh7_w60_0_c1 :  std_logic;
signal bh7_w61_0_c1 :  std_logic;
signal bh7_w62_0_c1 :  std_logic;
signal bh7_w63_0_c1 :  std_logic;
signal bh7_w64_0_c1 :  std_logic;
signal bh7_w65_0_c1 :  std_logic;
signal bh7_w66_0_c1 :  std_logic;
signal bh7_w67_0_c1 :  std_logic;
signal bh7_w68_0_c1 :  std_logic;
signal bh7_w69_0_c1 :  std_logic;
signal bh7_w70_0_c1 :  std_logic;
signal bh7_w71_0_c1 :  std_logic;
signal bh7_w72_0_c1 :  std_logic;
signal bh7_w73_0_c1 :  std_logic;
signal bh7_w74_0_c1 :  std_logic;
signal tile_3_X_c0 :  std_logic_vector(1 downto 0);
signal tile_3_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_3_output_c0 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w72_1_c0 :  std_logic;
signal bh7_w73_1_c0 :  std_logic;
signal bh7_w74_1_c0 :  std_logic;
signal bh7_w75_0_c0 :  std_logic;
signal bh7_w76_0_c0 :  std_logic;
signal tile_4_X_c0 :  std_logic_vector(1 downto 0);
signal tile_4_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_4_output_c0 :  std_logic_vector(4 downto 0);
signal tile_4_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w69_1_c0 :  std_logic;
signal bh7_w70_1_c0 :  std_logic;
signal bh7_w71_1_c0 :  std_logic;
signal bh7_w72_2_c0 :  std_logic;
signal bh7_w73_2_c0 :  std_logic;
signal tile_5_X_c0 :  std_logic_vector(1 downto 0);
signal tile_5_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_5_output_c0 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w66_1_c0 :  std_logic;
signal bh7_w67_1_c0 :  std_logic;
signal bh7_w68_1_c0 :  std_logic;
signal bh7_w69_2_c0 :  std_logic;
signal bh7_w70_2_c0 :  std_logic;
signal tile_6_X_c0 :  std_logic_vector(1 downto 0);
signal tile_6_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_6_output_c0 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w63_1_c0 :  std_logic;
signal bh7_w64_1_c0 :  std_logic;
signal bh7_w65_1_c0 :  std_logic;
signal bh7_w66_2_c0 :  std_logic;
signal bh7_w67_2_c0 :  std_logic;
signal tile_7_X_c0 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_7_output_c0 :  std_logic_vector(4 downto 0);
signal tile_7_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_1_c0 :  std_logic;
signal bh7_w61_1_c0 :  std_logic;
signal bh7_w62_1_c0 :  std_logic;
signal bh7_w63_2_c0 :  std_logic;
signal bh7_w64_2_c0 :  std_logic;
signal tile_8_X_c0 :  std_logic_vector(1 downto 0);
signal tile_8_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_8_output_c0 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_2_c0 :  std_logic;
signal bh7_w58_1_c0 :  std_logic;
signal bh7_w59_1_c0 :  std_logic;
signal bh7_w60_2_c0 :  std_logic;
signal bh7_w61_2_c0 :  std_logic;
signal tile_9_X_c0 :  std_logic_vector(1 downto 0);
signal tile_9_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_9_output_c0 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_2_c0 :  std_logic;
signal bh7_w55_2_c0 :  std_logic;
signal bh7_w56_2_c0 :  std_logic;
signal bh7_w57_3_c0 :  std_logic;
signal bh7_w58_2_c0 :  std_logic;
signal tile_10_X_c0 :  std_logic_vector(1 downto 0);
signal tile_10_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_10_output_c0 :  std_logic_vector(4 downto 0);
signal tile_10_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_2_c0 :  std_logic;
signal bh7_w52_2_c0 :  std_logic;
signal bh7_w53_2_c0 :  std_logic;
signal bh7_w54_3_c0 :  std_logic;
signal bh7_w55_3_c0 :  std_logic;
signal tile_11_X_c0 :  std_logic_vector(16 downto 0);
signal tile_11_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_11_output_c1 :  std_logic_vector(40 downto 0);
signal tile_11_filtered_output_c1 :  unsigned(40-0 downto 0);
signal bh7_w24_2_c1 :  std_logic;
signal bh7_w25_2_c1 :  std_logic;
signal bh7_w26_2_c1 :  std_logic;
signal bh7_w27_2_c1 :  std_logic;
signal bh7_w28_2_c1 :  std_logic;
signal bh7_w29_2_c1 :  std_logic;
signal bh7_w30_2_c1 :  std_logic;
signal bh7_w31_2_c1 :  std_logic;
signal bh7_w32_2_c1 :  std_logic;
signal bh7_w33_2_c1 :  std_logic;
signal bh7_w34_3_c1 :  std_logic;
signal bh7_w35_3_c1 :  std_logic;
signal bh7_w36_3_c1 :  std_logic;
signal bh7_w37_3_c1 :  std_logic;
signal bh7_w38_3_c1 :  std_logic;
signal bh7_w39_3_c1 :  std_logic;
signal bh7_w40_3_c1 :  std_logic;
signal bh7_w41_2_c1 :  std_logic;
signal bh7_w42_2_c1 :  std_logic;
signal bh7_w43_2_c1 :  std_logic;
signal bh7_w44_2_c1 :  std_logic;
signal bh7_w45_2_c1 :  std_logic;
signal bh7_w46_2_c1 :  std_logic;
signal bh7_w47_2_c1 :  std_logic;
signal bh7_w48_2_c1 :  std_logic;
signal bh7_w49_2_c1 :  std_logic;
signal bh7_w50_2_c1 :  std_logic;
signal bh7_w51_3_c1 :  std_logic;
signal bh7_w52_3_c1 :  std_logic;
signal bh7_w53_3_c1 :  std_logic;
signal bh7_w54_4_c1 :  std_logic;
signal bh7_w55_4_c1 :  std_logic;
signal bh7_w56_3_c1 :  std_logic;
signal bh7_w57_4_c1 :  std_logic;
signal bh7_w58_3_c1 :  std_logic;
signal bh7_w59_2_c1 :  std_logic;
signal bh7_w60_3_c1 :  std_logic;
signal bh7_w61_3_c1 :  std_logic;
signal bh7_w62_2_c1 :  std_logic;
signal bh7_w63_3_c1 :  std_logic;
signal bh7_w64_3_c1 :  std_logic;
signal tile_12_X_c0 :  std_logic_vector(16 downto 0);
signal tile_12_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_12_output_c1 :  std_logic_vector(40 downto 0);
signal tile_12_filtered_output_c1 :  unsigned(40-0 downto 0);
signal bh7_w41_3_c1 :  std_logic;
signal bh7_w42_3_c1 :  std_logic;
signal bh7_w43_3_c1 :  std_logic;
signal bh7_w44_3_c1 :  std_logic;
signal bh7_w45_3_c1 :  std_logic;
signal bh7_w46_3_c1 :  std_logic;
signal bh7_w47_3_c1 :  std_logic;
signal bh7_w48_3_c1 :  std_logic;
signal bh7_w49_3_c1 :  std_logic;
signal bh7_w50_3_c1 :  std_logic;
signal bh7_w51_4_c1 :  std_logic;
signal bh7_w52_4_c1 :  std_logic;
signal bh7_w53_4_c1 :  std_logic;
signal bh7_w54_5_c1 :  std_logic;
signal bh7_w55_5_c1 :  std_logic;
signal bh7_w56_4_c1 :  std_logic;
signal bh7_w57_5_c1 :  std_logic;
signal bh7_w58_4_c1 :  std_logic;
signal bh7_w59_3_c1 :  std_logic;
signal bh7_w60_4_c1 :  std_logic;
signal bh7_w61_4_c1 :  std_logic;
signal bh7_w62_3_c1 :  std_logic;
signal bh7_w63_4_c1 :  std_logic;
signal bh7_w64_4_c1 :  std_logic;
signal bh7_w65_2_c1 :  std_logic;
signal bh7_w66_3_c1 :  std_logic;
signal bh7_w67_3_c1 :  std_logic;
signal bh7_w68_2_c1 :  std_logic;
signal bh7_w69_3_c1 :  std_logic;
signal bh7_w70_3_c1 :  std_logic;
signal bh7_w71_2_c1 :  std_logic;
signal bh7_w72_3_c1 :  std_logic;
signal bh7_w73_3_c1 :  std_logic;
signal bh7_w74_2_c1 :  std_logic;
signal bh7_w75_1_c1 :  std_logic;
signal bh7_w76_1_c1 :  std_logic;
signal bh7_w77_0_c1 :  std_logic;
signal bh7_w78_0_c1 :  std_logic;
signal bh7_w79_0_c1 :  std_logic;
signal bh7_w80_0_c1 :  std_logic;
signal bh7_w81_0_c1 :  std_logic;
signal tile_13_X_c0 :  std_logic_vector(16 downto 0);
signal tile_13_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_13_output_c1 :  std_logic_vector(40 downto 0);
signal tile_13_filtered_output_c1 :  unsigned(40-0 downto 0);
signal bh7_w58_5_c1 :  std_logic;
signal bh7_w59_4_c1 :  std_logic;
signal bh7_w60_5_c1 :  std_logic;
signal bh7_w61_5_c1 :  std_logic;
signal bh7_w62_4_c1 :  std_logic;
signal bh7_w63_5_c1 :  std_logic;
signal bh7_w64_5_c1 :  std_logic;
signal bh7_w65_3_c1 :  std_logic;
signal bh7_w66_4_c1 :  std_logic;
signal bh7_w67_4_c1 :  std_logic;
signal bh7_w68_3_c1 :  std_logic;
signal bh7_w69_4_c1 :  std_logic;
signal bh7_w70_4_c1 :  std_logic;
signal bh7_w71_3_c1 :  std_logic;
signal bh7_w72_4_c1 :  std_logic;
signal bh7_w73_4_c1 :  std_logic;
signal bh7_w74_3_c1 :  std_logic;
signal bh7_w75_2_c1 :  std_logic;
signal bh7_w76_2_c1 :  std_logic;
signal bh7_w77_1_c1 :  std_logic;
signal bh7_w78_1_c1 :  std_logic;
signal bh7_w79_1_c1 :  std_logic;
signal bh7_w80_1_c1 :  std_logic;
signal bh7_w81_1_c1 :  std_logic;
signal bh7_w82_0_c1 :  std_logic;
signal bh7_w83_0_c1 :  std_logic;
signal bh7_w84_0_c1 :  std_logic;
signal bh7_w85_0_c1 :  std_logic;
signal bh7_w86_0_c1 :  std_logic;
signal bh7_w87_0_c1 :  std_logic;
signal bh7_w88_0_c1 :  std_logic;
signal bh7_w89_0_c1 :  std_logic;
signal bh7_w90_0_c1 :  std_logic;
signal bh7_w91_0_c1 :  std_logic;
signal bh7_w92_0_c1 :  std_logic;
signal bh7_w93_0_c1 :  std_logic;
signal bh7_w94_0_c1 :  std_logic;
signal bh7_w95_0_c1 :  std_logic;
signal bh7_w96_0_c1 :  std_logic;
signal bh7_w97_0_c1 :  std_logic;
signal bh7_w98_0_c1 :  std_logic;
signal tile_14_X_c0 :  std_logic_vector(1 downto 0);
signal tile_14_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_14_output_c0 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_1_c0 :  std_logic;
signal bh7_w97_1_c0 :  std_logic;
signal bh7_w98_1_c0 :  std_logic;
signal bh7_w99_0_c0 :  std_logic;
signal bh7_w100_0_c0 :  std_logic;
signal tile_15_X_c0 :  std_logic_vector(1 downto 0);
signal tile_15_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_15_output_c0 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_1_c0 :  std_logic;
signal bh7_w94_1_c0 :  std_logic;
signal bh7_w95_1_c0 :  std_logic;
signal bh7_w96_2_c0 :  std_logic;
signal bh7_w97_2_c0 :  std_logic;
signal tile_16_X_c0 :  std_logic_vector(1 downto 0);
signal tile_16_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_16_output_c0 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_1_c0 :  std_logic;
signal bh7_w91_1_c0 :  std_logic;
signal bh7_w92_1_c0 :  std_logic;
signal bh7_w93_2_c0 :  std_logic;
signal bh7_w94_2_c0 :  std_logic;
signal tile_17_X_c0 :  std_logic_vector(1 downto 0);
signal tile_17_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_17_output_c0 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_1_c0 :  std_logic;
signal bh7_w88_1_c0 :  std_logic;
signal bh7_w89_1_c0 :  std_logic;
signal bh7_w90_2_c0 :  std_logic;
signal bh7_w91_2_c0 :  std_logic;
signal tile_18_X_c0 :  std_logic_vector(1 downto 0);
signal tile_18_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_18_output_c0 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_1_c0 :  std_logic;
signal bh7_w85_1_c0 :  std_logic;
signal bh7_w86_1_c0 :  std_logic;
signal bh7_w87_2_c0 :  std_logic;
signal bh7_w88_2_c0 :  std_logic;
signal tile_19_X_c0 :  std_logic_vector(1 downto 0);
signal tile_19_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_19_output_c0 :  std_logic_vector(4 downto 0);
signal tile_19_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w81_2_c0 :  std_logic;
signal bh7_w82_1_c0 :  std_logic;
signal bh7_w83_1_c0 :  std_logic;
signal bh7_w84_2_c0 :  std_logic;
signal bh7_w85_2_c0 :  std_logic;
signal tile_20_X_c0 :  std_logic_vector(1 downto 0);
signal tile_20_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_20_output_c0 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w78_2_c0 :  std_logic;
signal bh7_w79_2_c0 :  std_logic;
signal bh7_w80_2_c0 :  std_logic;
signal bh7_w81_3_c0 :  std_logic;
signal bh7_w82_2_c0 :  std_logic;
signal tile_21_X_c0 :  std_logic_vector(1 downto 0);
signal tile_21_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_21_output_c0 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w75_3_c0 :  std_logic;
signal bh7_w76_3_c0 :  std_logic;
signal bh7_w77_2_c0 :  std_logic;
signal bh7_w78_3_c0 :  std_logic;
signal bh7_w79_3_c0 :  std_logic;
signal tile_22_X_c0 :  std_logic_vector(0 downto 0);
signal tile_22_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_22_output_c0 :  std_logic_vector(0 downto 0);
signal tile_22_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w68_4_c0 :  std_logic;
signal tile_23_X_c0 :  std_logic_vector(3 downto 0);
signal tile_23_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_23_output_c0 :  std_logic_vector(3 downto 0);
signal tile_23_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w64_6_c0 :  std_logic;
signal bh7_w65_4_c0 :  std_logic;
signal bh7_w66_5_c0 :  std_logic;
signal bh7_w67_5_c0 :  std_logic;
signal tile_24_X_c0 :  std_logic_vector(3 downto 0);
signal tile_24_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_24_output_c0 :  std_logic_vector(3 downto 0);
signal tile_24_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w60_6_c0 :  std_logic;
signal bh7_w61_6_c0 :  std_logic;
signal bh7_w62_5_c0 :  std_logic;
signal bh7_w63_6_c0 :  std_logic;
signal tile_25_X_c0 :  std_logic_vector(3 downto 0);
signal tile_25_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_25_output_c0 :  std_logic_vector(3 downto 0);
signal tile_25_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w56_5_c0 :  std_logic;
signal bh7_w57_6_c0 :  std_logic;
signal bh7_w58_6_c0 :  std_logic;
signal bh7_w59_5_c0 :  std_logic;
signal tile_26_X_c0 :  std_logic_vector(3 downto 0);
signal tile_26_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_26_output_c0 :  std_logic_vector(3 downto 0);
signal tile_26_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w52_5_c0 :  std_logic;
signal bh7_w53_5_c0 :  std_logic;
signal bh7_w54_6_c0 :  std_logic;
signal bh7_w55_6_c0 :  std_logic;
signal tile_27_X_c0 :  std_logic_vector(1 downto 0);
signal tile_27_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_27_output_c0 :  std_logic_vector(3 downto 0);
signal tile_27_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w65_5_c0 :  std_logic;
signal bh7_w66_6_c0 :  std_logic;
signal bh7_w67_6_c0 :  std_logic;
signal bh7_w68_5_c0 :  std_logic;
signal tile_28_X_c0 :  std_logic_vector(2 downto 0);
signal tile_28_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_28_output_c0 :  std_logic_vector(4 downto 0);
signal tile_28_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w62_6_c0 :  std_logic;
signal bh7_w63_7_c0 :  std_logic;
signal bh7_w64_7_c0 :  std_logic;
signal bh7_w65_6_c0 :  std_logic;
signal bh7_w66_7_c0 :  std_logic;
signal tile_29_X_c0 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_29_output_c0 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w59_6_c0 :  std_logic;
signal bh7_w60_7_c0 :  std_logic;
signal bh7_w61_7_c0 :  std_logic;
signal bh7_w62_7_c0 :  std_logic;
signal bh7_w63_8_c0 :  std_logic;
signal tile_30_X_c0 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_30_output_c0 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w56_6_c0 :  std_logic;
signal bh7_w57_7_c0 :  std_logic;
signal bh7_w58_7_c0 :  std_logic;
signal bh7_w59_7_c0 :  std_logic;
signal bh7_w60_8_c0 :  std_logic;
signal tile_31_X_c0 :  std_logic_vector(2 downto 0);
signal tile_31_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_31_output_c0 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w53_6_c0 :  std_logic;
signal bh7_w54_7_c0 :  std_logic;
signal bh7_w55_7_c0 :  std_logic;
signal bh7_w56_7_c0 :  std_logic;
signal bh7_w57_8_c0 :  std_logic;
signal tile_32_X_c0 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_32_output_c0 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w50_4_c0 :  std_logic;
signal bh7_w51_5_c0 :  std_logic;
signal bh7_w52_6_c0 :  std_logic;
signal bh7_w53_7_c0 :  std_logic;
signal bh7_w54_8_c0 :  std_logic;
signal tile_33_X_c0 :  std_logic_vector(1 downto 0);
signal tile_33_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_33_output_c0 :  std_logic_vector(3 downto 0);
signal tile_33_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w63_9_c0 :  std_logic;
signal bh7_w64_8_c0 :  std_logic;
signal bh7_w65_7_c0 :  std_logic;
signal bh7_w66_8_c0 :  std_logic;
signal tile_34_X_c0 :  std_logic_vector(2 downto 0);
signal tile_34_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_34_output_c0 :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_9_c0 :  std_logic;
signal bh7_w61_8_c0 :  std_logic;
signal bh7_w62_8_c0 :  std_logic;
signal bh7_w63_10_c0 :  std_logic;
signal bh7_w64_9_c0 :  std_logic;
signal tile_35_X_c0 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_35_output_c0 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_9_c0 :  std_logic;
signal bh7_w58_8_c0 :  std_logic;
signal bh7_w59_8_c0 :  std_logic;
signal bh7_w60_10_c0 :  std_logic;
signal bh7_w61_9_c0 :  std_logic;
signal tile_36_X_c0 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_36_output_c0 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_9_c0 :  std_logic;
signal bh7_w55_8_c0 :  std_logic;
signal bh7_w56_8_c0 :  std_logic;
signal bh7_w57_10_c0 :  std_logic;
signal bh7_w58_9_c0 :  std_logic;
signal tile_37_X_c0 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_37_output_c0 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_6_c0 :  std_logic;
signal bh7_w52_7_c0 :  std_logic;
signal bh7_w53_8_c0 :  std_logic;
signal bh7_w54_10_c0 :  std_logic;
signal bh7_w55_9_c0 :  std_logic;
signal tile_38_X_c0 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_38_output_c0 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w48_4_c0, bh7_w48_4_c1 :  std_logic;
signal bh7_w49_4_c0 :  std_logic;
signal bh7_w50_5_c0 :  std_logic;
signal bh7_w51_7_c0 :  std_logic;
signal bh7_w52_8_c0 :  std_logic;
signal tile_39_X_c0 :  std_logic_vector(0 downto 0);
signal tile_39_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_39_output_c0 :  std_logic_vector(0 downto 0);
signal tile_39_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w85_3_c0 :  std_logic;
signal tile_40_X_c0 :  std_logic_vector(3 downto 0);
signal tile_40_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_40_output_c0 :  std_logic_vector(3 downto 0);
signal tile_40_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w81_4_c0 :  std_logic;
signal bh7_w82_3_c0 :  std_logic;
signal bh7_w83_2_c0 :  std_logic;
signal bh7_w84_3_c0 :  std_logic;
signal tile_41_X_c0 :  std_logic_vector(3 downto 0);
signal tile_41_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_41_output_c0 :  std_logic_vector(3 downto 0);
signal tile_41_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w77_3_c0 :  std_logic;
signal bh7_w78_4_c0 :  std_logic;
signal bh7_w79_4_c0 :  std_logic;
signal bh7_w80_3_c0 :  std_logic;
signal tile_42_X_c0 :  std_logic_vector(3 downto 0);
signal tile_42_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_42_output_c0 :  std_logic_vector(3 downto 0);
signal tile_42_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w73_5_c0 :  std_logic;
signal bh7_w74_4_c0 :  std_logic;
signal bh7_w75_4_c0 :  std_logic;
signal bh7_w76_4_c0 :  std_logic;
signal tile_43_X_c0 :  std_logic_vector(3 downto 0);
signal tile_43_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_43_output_c0 :  std_logic_vector(3 downto 0);
signal tile_43_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w69_5_c0 :  std_logic;
signal bh7_w70_5_c0 :  std_logic;
signal bh7_w71_4_c0 :  std_logic;
signal bh7_w72_5_c0 :  std_logic;
signal tile_44_X_c0 :  std_logic_vector(1 downto 0);
signal tile_44_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_44_output_c0 :  std_logic_vector(3 downto 0);
signal tile_44_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w82_4_c0 :  std_logic;
signal bh7_w83_3_c0 :  std_logic;
signal bh7_w84_4_c0 :  std_logic;
signal bh7_w85_4_c0 :  std_logic;
signal tile_45_X_c0 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_45_output_c0 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w79_5_c0 :  std_logic;
signal bh7_w80_4_c0 :  std_logic;
signal bh7_w81_5_c0 :  std_logic;
signal bh7_w82_5_c0 :  std_logic;
signal bh7_w83_4_c0 :  std_logic;
signal tile_46_X_c0 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_46_output_c0 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w76_5_c0 :  std_logic;
signal bh7_w77_4_c0 :  std_logic;
signal bh7_w78_5_c0 :  std_logic;
signal bh7_w79_6_c0 :  std_logic;
signal bh7_w80_5_c0 :  std_logic;
signal tile_47_X_c0 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_47_output_c0 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w73_6_c0 :  std_logic;
signal bh7_w74_5_c0 :  std_logic;
signal bh7_w75_5_c0 :  std_logic;
signal bh7_w76_6_c0 :  std_logic;
signal bh7_w77_5_c0 :  std_logic;
signal tile_48_X_c0 :  std_logic_vector(2 downto 0);
signal tile_48_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_48_output_c0 :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w70_6_c0 :  std_logic;
signal bh7_w71_5_c0 :  std_logic;
signal bh7_w72_6_c0 :  std_logic;
signal bh7_w73_7_c0 :  std_logic;
signal bh7_w74_6_c0 :  std_logic;
signal tile_49_X_c0 :  std_logic_vector(2 downto 0);
signal tile_49_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_49_output_c0 :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w67_7_c0 :  std_logic;
signal bh7_w68_6_c0 :  std_logic;
signal bh7_w69_6_c0 :  std_logic;
signal bh7_w70_7_c0 :  std_logic;
signal bh7_w71_6_c0 :  std_logic;
signal tile_50_X_c0 :  std_logic_vector(1 downto 0);
signal tile_50_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_50_output_c0 :  std_logic_vector(3 downto 0);
signal tile_50_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w80_6_c0 :  std_logic;
signal bh7_w81_6_c0 :  std_logic;
signal bh7_w82_6_c0 :  std_logic;
signal bh7_w83_5_c0 :  std_logic;
signal tile_51_X_c0 :  std_logic_vector(2 downto 0);
signal tile_51_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_51_output_c0 :  std_logic_vector(4 downto 0);
signal tile_51_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w77_6_c0 :  std_logic;
signal bh7_w78_6_c0 :  std_logic;
signal bh7_w79_7_c0 :  std_logic;
signal bh7_w80_7_c0 :  std_logic;
signal bh7_w81_7_c0 :  std_logic;
signal tile_52_X_c0 :  std_logic_vector(2 downto 0);
signal tile_52_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_52_output_c0 :  std_logic_vector(4 downto 0);
signal tile_52_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w74_7_c0 :  std_logic;
signal bh7_w75_6_c0 :  std_logic;
signal bh7_w76_7_c0 :  std_logic;
signal bh7_w77_7_c0 :  std_logic;
signal bh7_w78_7_c0 :  std_logic;
signal tile_53_X_c0 :  std_logic_vector(2 downto 0);
signal tile_53_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_53_output_c0 :  std_logic_vector(4 downto 0);
signal tile_53_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w71_7_c0 :  std_logic;
signal bh7_w72_7_c0 :  std_logic;
signal bh7_w73_8_c0 :  std_logic;
signal bh7_w74_8_c0 :  std_logic;
signal bh7_w75_7_c0 :  std_logic;
signal tile_54_X_c0 :  std_logic_vector(2 downto 0);
signal tile_54_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_54_output_c0 :  std_logic_vector(4 downto 0);
signal tile_54_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w68_7_c0 :  std_logic;
signal bh7_w69_7_c0 :  std_logic;
signal bh7_w70_8_c0 :  std_logic;
signal bh7_w71_8_c0 :  std_logic;
signal bh7_w72_8_c0 :  std_logic;
signal tile_55_X_c0 :  std_logic_vector(2 downto 0);
signal tile_55_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_55_output_c0 :  std_logic_vector(4 downto 0);
signal tile_55_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w65_8_c0 :  std_logic;
signal bh7_w66_9_c0 :  std_logic;
signal bh7_w67_8_c0 :  std_logic;
signal bh7_w68_8_c0 :  std_logic;
signal bh7_w69_8_c0 :  std_logic;
signal tile_56_X_c0 :  std_logic_vector(0 downto 0);
signal tile_56_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_56_output_c0 :  std_logic_vector(0 downto 0);
signal tile_56_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w102_0_c0 :  std_logic;
signal tile_57_X_c0 :  std_logic_vector(3 downto 0);
signal tile_57_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_57_output_c0 :  std_logic_vector(3 downto 0);
signal tile_57_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w98_2_c0 :  std_logic;
signal bh7_w99_1_c0 :  std_logic;
signal bh7_w100_1_c0 :  std_logic;
signal bh7_w101_0_c0 :  std_logic;
signal tile_58_X_c0 :  std_logic_vector(3 downto 0);
signal tile_58_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_58_output_c0 :  std_logic_vector(3 downto 0);
signal tile_58_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w94_3_c0 :  std_logic;
signal bh7_w95_2_c0 :  std_logic;
signal bh7_w96_3_c0 :  std_logic;
signal bh7_w97_3_c0 :  std_logic;
signal tile_59_X_c0 :  std_logic_vector(3 downto 0);
signal tile_59_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_59_output_c0 :  std_logic_vector(3 downto 0);
signal tile_59_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w90_3_c0 :  std_logic;
signal bh7_w91_3_c0 :  std_logic;
signal bh7_w92_2_c0 :  std_logic;
signal bh7_w93_3_c0 :  std_logic;
signal tile_60_X_c0 :  std_logic_vector(3 downto 0);
signal tile_60_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_60_output_c0 :  std_logic_vector(3 downto 0);
signal tile_60_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w86_2_c0 :  std_logic;
signal bh7_w87_3_c0 :  std_logic;
signal bh7_w88_3_c0 :  std_logic;
signal bh7_w89_2_c0 :  std_logic;
signal tile_61_X_c0 :  std_logic_vector(1 downto 0);
signal tile_61_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_61_output_c0 :  std_logic_vector(3 downto 0);
signal tile_61_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w99_2_c0 :  std_logic;
signal bh7_w100_2_c0 :  std_logic;
signal bh7_w101_1_c0 :  std_logic;
signal bh7_w102_1_c0 :  std_logic;
signal tile_62_X_c0 :  std_logic_vector(2 downto 0);
signal tile_62_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_62_output_c0 :  std_logic_vector(4 downto 0);
signal tile_62_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_4_c0 :  std_logic;
signal bh7_w97_4_c0 :  std_logic;
signal bh7_w98_3_c0 :  std_logic;
signal bh7_w99_3_c0 :  std_logic;
signal bh7_w100_3_c0 :  std_logic;
signal tile_63_X_c0 :  std_logic_vector(2 downto 0);
signal tile_63_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_63_output_c0 :  std_logic_vector(4 downto 0);
signal tile_63_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_4_c0 :  std_logic;
signal bh7_w94_4_c0 :  std_logic;
signal bh7_w95_3_c0 :  std_logic;
signal bh7_w96_5_c0 :  std_logic;
signal bh7_w97_5_c0 :  std_logic;
signal tile_64_X_c0 :  std_logic_vector(2 downto 0);
signal tile_64_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_64_output_c0 :  std_logic_vector(4 downto 0);
signal tile_64_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_4_c0 :  std_logic;
signal bh7_w91_4_c0 :  std_logic;
signal bh7_w92_3_c0 :  std_logic;
signal bh7_w93_5_c0 :  std_logic;
signal bh7_w94_5_c0 :  std_logic;
signal tile_65_X_c0 :  std_logic_vector(2 downto 0);
signal tile_65_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_65_output_c0 :  std_logic_vector(4 downto 0);
signal tile_65_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_4_c0 :  std_logic;
signal bh7_w88_4_c0 :  std_logic;
signal bh7_w89_3_c0 :  std_logic;
signal bh7_w90_5_c0 :  std_logic;
signal bh7_w91_5_c0 :  std_logic;
signal tile_66_X_c0 :  std_logic_vector(2 downto 0);
signal tile_66_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_66_output_c0 :  std_logic_vector(4 downto 0);
signal tile_66_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_5_c0 :  std_logic;
signal bh7_w85_5_c0 :  std_logic;
signal bh7_w86_3_c0 :  std_logic;
signal bh7_w87_5_c0 :  std_logic;
signal bh7_w88_5_c0 :  std_logic;
signal tile_67_X_c0 :  std_logic_vector(1 downto 0);
signal tile_67_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_67_output_c0 :  std_logic_vector(3 downto 0);
signal tile_67_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w97_6_c0 :  std_logic;
signal bh7_w98_4_c0 :  std_logic;
signal bh7_w99_4_c0 :  std_logic;
signal bh7_w100_4_c0 :  std_logic;
signal tile_68_X_c0 :  std_logic_vector(2 downto 0);
signal tile_68_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_68_output_c0 :  std_logic_vector(4 downto 0);
signal tile_68_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w94_6_c0 :  std_logic;
signal bh7_w95_4_c0 :  std_logic;
signal bh7_w96_6_c0 :  std_logic;
signal bh7_w97_7_c0 :  std_logic;
signal bh7_w98_5_c0 :  std_logic;
signal tile_69_X_c0 :  std_logic_vector(2 downto 0);
signal tile_69_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_69_output_c0 :  std_logic_vector(4 downto 0);
signal tile_69_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w91_6_c0 :  std_logic;
signal bh7_w92_4_c0 :  std_logic;
signal bh7_w93_6_c0 :  std_logic;
signal bh7_w94_7_c0 :  std_logic;
signal bh7_w95_5_c0 :  std_logic;
signal tile_70_X_c0 :  std_logic_vector(2 downto 0);
signal tile_70_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_70_output_c0 :  std_logic_vector(4 downto 0);
signal tile_70_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w88_6_c0 :  std_logic;
signal bh7_w89_4_c0 :  std_logic;
signal bh7_w90_6_c0 :  std_logic;
signal bh7_w91_7_c0 :  std_logic;
signal bh7_w92_5_c0 :  std_logic;
signal tile_71_X_c0 :  std_logic_vector(2 downto 0);
signal tile_71_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_71_output_c0 :  std_logic_vector(4 downto 0);
signal tile_71_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w85_6_c0 :  std_logic;
signal bh7_w86_4_c0 :  std_logic;
signal bh7_w87_6_c0 :  std_logic;
signal bh7_w88_7_c0 :  std_logic;
signal bh7_w89_5_c0 :  std_logic;
signal tile_72_X_c0 :  std_logic_vector(2 downto 0);
signal tile_72_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_72_output_c0 :  std_logic_vector(4 downto 0);
signal tile_72_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w82_7_c0 :  std_logic;
signal bh7_w83_6_c0 :  std_logic;
signal bh7_w84_6_c0 :  std_logic;
signal bh7_w85_7_c0 :  std_logic;
signal bh7_w86_5_c0 :  std_logic;
signal tile_73_X_c0 :  std_logic_vector(1 downto 0);
signal tile_73_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_73_output_c0 :  std_logic_vector(3 downto 0);
signal tile_73_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w102_2_c0 :  std_logic;
signal bh7_w103_0_c0 :  std_logic;
signal bh7_w104_0_c0 :  std_logic;
signal bh7_w105_0_c0 :  std_logic;
signal tile_74_X_c0 :  std_logic_vector(1 downto 0);
signal tile_74_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_74_output_c0 :  std_logic_vector(4 downto 0);
signal tile_74_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w99_5_c0 :  std_logic;
signal bh7_w100_5_c0 :  std_logic;
signal bh7_w101_2_c0 :  std_logic;
signal bh7_w102_3_c0 :  std_logic;
signal bh7_w103_1_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid323_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid323_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid323_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w49_5_c0 :  std_logic;
signal bh7_w50_6_c0 :  std_logic;
signal bh7_w51_8_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid323_Out0_copy324_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid327_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid327_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid327_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w51_9_c0 :  std_logic;
signal bh7_w52_9_c0 :  std_logic;
signal bh7_w53_9_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid327_Out0_copy328_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid329_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid329_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid329_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w52_10_c0 :  std_logic;
signal bh7_w53_10_c0 :  std_logic;
signal bh7_w54_11_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid329_Out0_copy330_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid331_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid331_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid331_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w53_11_c0 :  std_logic;
signal bh7_w54_12_c0 :  std_logic;
signal bh7_w55_10_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid331_Out0_copy332_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid335_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid335_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w54_13_c0 :  std_logic;
signal bh7_w55_11_c0 :  std_logic;
signal bh7_w56_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid335_Out0_copy336_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid337_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid337_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w55_12_c0 :  std_logic;
signal bh7_w56_10_c0 :  std_logic;
signal bh7_w57_11_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid337_Out0_copy338_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid339_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid339_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid339_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w56_11_c0 :  std_logic;
signal bh7_w57_12_c0 :  std_logic;
signal bh7_w58_10_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid339_Out0_copy340_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid341_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid341_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w57_13_c0 :  std_logic;
signal bh7_w58_11_c0 :  std_logic;
signal bh7_w59_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid341_Out0_copy342_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid343_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid343_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w58_12_c0 :  std_logic;
signal bh7_w59_10_c0 :  std_logic;
signal bh7_w60_11_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid343_Out0_copy344_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid345_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid345_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid345_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w59_11_c0 :  std_logic;
signal bh7_w60_12_c0 :  std_logic;
signal bh7_w61_10_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid345_Out0_copy346_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid347_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid347_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w60_13_c0 :  std_logic;
signal bh7_w61_11_c0 :  std_logic;
signal bh7_w62_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid347_Out0_copy348_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid349_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid349_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w61_12_c0 :  std_logic;
signal bh7_w62_10_c0 :  std_logic;
signal bh7_w63_11_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid349_Out0_copy350_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid351_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid351_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid351_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w62_11_c0 :  std_logic;
signal bh7_w63_12_c0 :  std_logic;
signal bh7_w64_10_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid351_Out0_copy352_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid353_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid353_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w63_13_c0 :  std_logic;
signal bh7_w64_11_c0 :  std_logic;
signal bh7_w65_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid353_Out0_copy354_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid355_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid355_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w64_12_c0 :  std_logic;
signal bh7_w65_10_c0 :  std_logic;
signal bh7_w66_10_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid355_Out0_copy356_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid357_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid357_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w65_11_c0 :  std_logic;
signal bh7_w66_11_c0 :  std_logic;
signal bh7_w67_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid357_Out0_copy358_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid359_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid359_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_12_c0 :  std_logic;
signal bh7_w67_10_c0 :  std_logic;
signal bh7_w68_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid359_Out0_copy360_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid361_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid361_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w67_11_c0 :  std_logic;
signal bh7_w68_10_c0 :  std_logic;
signal bh7_w69_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid361_Out0_copy362_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid363_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid363_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_11_c0 :  std_logic;
signal bh7_w69_10_c0 :  std_logic;
signal bh7_w70_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid363_Out0_copy364_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid365_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid365_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w69_11_c0 :  std_logic;
signal bh7_w70_10_c0 :  std_logic;
signal bh7_w71_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid365_Out0_copy366_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid367_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid367_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_11_c0 :  std_logic;
signal bh7_w71_10_c0 :  std_logic;
signal bh7_w72_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid367_Out0_copy368_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid369_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid369_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w71_11_c0 :  std_logic;
signal bh7_w72_10_c0 :  std_logic;
signal bh7_w73_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid369_Out0_copy370_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid371_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid371_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_11_c0 :  std_logic;
signal bh7_w73_10_c0 :  std_logic;
signal bh7_w74_9_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid371_Out0_copy372_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid373_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid373_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w73_11_c0 :  std_logic;
signal bh7_w74_10_c0 :  std_logic;
signal bh7_w75_8_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid373_Out0_copy374_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid375_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid375_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_11_c0 :  std_logic;
signal bh7_w75_9_c0 :  std_logic;
signal bh7_w76_8_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid375_Out0_copy376_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid377_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid377_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w75_10_c0 :  std_logic;
signal bh7_w76_9_c0 :  std_logic;
signal bh7_w77_8_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid377_Out0_copy378_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid379_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid379_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_10_c0 :  std_logic;
signal bh7_w77_9_c0 :  std_logic;
signal bh7_w78_8_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid379_Out0_copy380_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid381_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid381_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w77_10_c0 :  std_logic;
signal bh7_w78_9_c0 :  std_logic;
signal bh7_w79_8_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid381_Out0_copy382_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid383_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid383_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_10_c0 :  std_logic;
signal bh7_w79_9_c0 :  std_logic;
signal bh7_w80_8_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid383_Out0_copy384_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid385_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid385_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w79_10_c0 :  std_logic;
signal bh7_w80_9_c0 :  std_logic;
signal bh7_w81_8_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid385_Out0_copy386_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid387_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid387_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_10_c0 :  std_logic;
signal bh7_w81_9_c0 :  std_logic;
signal bh7_w82_8_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid387_Out0_copy388_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid389_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid389_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w81_10_c0 :  std_logic;
signal bh7_w82_9_c0 :  std_logic;
signal bh7_w83_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid389_Out0_copy390_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid391_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid391_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_10_c0 :  std_logic;
signal bh7_w83_8_c0 :  std_logic;
signal bh7_w84_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid391_Out0_copy392_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid393_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid393_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w83_9_c0 :  std_logic;
signal bh7_w84_8_c0 :  std_logic;
signal bh7_w85_8_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid393_Out0_copy394_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid395_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid395_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w84_9_c0 :  std_logic;
signal bh7_w85_9_c0 :  std_logic;
signal bh7_w86_6_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid395_Out0_copy396_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid397_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid397_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w85_10_c0 :  std_logic;
signal bh7_w86_7_c0 :  std_logic;
signal bh7_w87_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid397_Out0_copy398_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid401_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid401_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w86_8_c0 :  std_logic;
signal bh7_w87_8_c0 :  std_logic;
signal bh7_w88_8_c0 :  std_logic;
signal Compressor_5_3_Freq500_uid400_bh7_uid401_Out0_copy402_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid403_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid403_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w87_9_c0 :  std_logic;
signal bh7_w88_9_c0 :  std_logic;
signal bh7_w89_6_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid403_Out0_copy404_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid405_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid405_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w88_10_c0 :  std_logic;
signal bh7_w89_7_c0 :  std_logic;
signal bh7_w90_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid405_Out0_copy406_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid407_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid407_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w89_8_c0 :  std_logic;
signal bh7_w90_8_c0 :  std_logic;
signal bh7_w91_8_c0 :  std_logic;
signal Compressor_5_3_Freq500_uid400_bh7_uid407_Out0_copy408_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid409_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid409_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w90_9_c0 :  std_logic;
signal bh7_w91_9_c0 :  std_logic;
signal bh7_w92_6_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid409_Out0_copy410_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid411_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid411_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w91_10_c0 :  std_logic;
signal bh7_w92_7_c0 :  std_logic;
signal bh7_w93_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid411_Out0_copy412_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid413_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid413_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w92_8_c0 :  std_logic;
signal bh7_w93_8_c0 :  std_logic;
signal bh7_w94_8_c0 :  std_logic;
signal Compressor_5_3_Freq500_uid400_bh7_uid413_Out0_copy414_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid415_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid415_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w93_9_c0 :  std_logic;
signal bh7_w94_9_c0 :  std_logic;
signal bh7_w95_6_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid415_Out0_copy416_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid417_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid417_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w94_10_c0 :  std_logic;
signal bh7_w95_7_c0 :  std_logic;
signal bh7_w96_7_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid417_Out0_copy418_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid419_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid419_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w95_8_c0 :  std_logic;
signal bh7_w96_8_c0 :  std_logic;
signal bh7_w97_8_c0 :  std_logic;
signal Compressor_5_3_Freq500_uid400_bh7_uid419_Out0_copy420_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid421_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid421_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w96_9_c0 :  std_logic;
signal bh7_w97_9_c0 :  std_logic;
signal bh7_w98_6_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid421_Out0_copy422_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid423_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid423_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w97_10_c0 :  std_logic;
signal bh7_w98_7_c0 :  std_logic;
signal bh7_w99_6_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid423_Out0_copy424_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid425_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid425_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w98_8_c0 :  std_logic;
signal bh7_w99_7_c0 :  std_logic;
signal bh7_w100_6_c0 :  std_logic;
signal Compressor_5_3_Freq500_uid400_bh7_uid425_Out0_copy426_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid427_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid427_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w99_8_c0 :  std_logic;
signal bh7_w100_7_c0 :  std_logic;
signal bh7_w101_3_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid427_Out0_copy428_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid429_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid429_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w100_8_c0 :  std_logic;
signal bh7_w101_4_c0 :  std_logic;
signal bh7_w102_4_c0 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid429_Out0_copy430_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid433_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid433_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w101_5_c0 :  std_logic;
signal bh7_w102_5_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid433_Out0_copy434_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid435_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid435_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid435_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w102_6_c0 :  std_logic;
signal bh7_w103_2_c0 :  std_logic;
signal bh7_w104_1_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid435_Out0_copy436_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid437_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid437_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid437_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w51_10_c0 :  std_logic;
signal bh7_w52_11_c0 :  std_logic;
signal bh7_w53_12_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid437_Out0_copy438_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid439_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid439_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid439_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w53_13_c0 :  std_logic;
signal bh7_w54_14_c0 :  std_logic;
signal bh7_w55_13_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid439_Out0_copy440_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid441_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid441_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w55_14_c0 :  std_logic;
signal bh7_w56_12_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid441_Out0_copy442_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid443_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid443_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid443_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w56_13_c0 :  std_logic;
signal bh7_w57_14_c0 :  std_logic;
signal bh7_w58_13_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid443_Out0_copy444_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid445_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid445_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w57_15_c0 :  std_logic;
signal bh7_w58_14_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid445_Out0_copy446_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid447_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid447_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w58_15_c0 :  std_logic;
signal bh7_w59_12_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid447_Out0_copy448_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid449_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid449_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid449_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w59_13_c0 :  std_logic;
signal bh7_w60_14_c0 :  std_logic;
signal bh7_w61_13_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid449_Out0_copy450_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid451_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid451_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w60_15_c0 :  std_logic;
signal bh7_w61_14_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid451_Out0_copy452_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid453_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid453_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w61_15_c0 :  std_logic;
signal bh7_w62_12_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid453_Out0_copy454_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid455_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid455_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid455_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w62_13_c0 :  std_logic;
signal bh7_w63_14_c0 :  std_logic;
signal bh7_w64_13_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid455_Out0_copy456_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid457_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid457_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w63_15_c0 :  std_logic;
signal bh7_w64_14_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid457_Out0_copy458_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid459_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid459_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid459_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w64_15_c0 :  std_logic;
signal bh7_w65_12_c0 :  std_logic;
signal bh7_w66_13_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid459_Out0_copy460_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid461_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid461_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid461_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_14_c0 :  std_logic;
signal bh7_w67_12_c0 :  std_logic;
signal bh7_w68_12_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid461_Out0_copy462_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid463_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid463_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w67_13_c0 :  std_logic;
signal bh7_w68_13_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid463_Out0_copy464_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid465_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid465_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid465_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_14_c0 :  std_logic;
signal bh7_w69_12_c0 :  std_logic;
signal bh7_w70_12_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid465_Out0_copy466_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid467_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid467_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid467_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_13_c0 :  std_logic;
signal bh7_w71_12_c0 :  std_logic;
signal bh7_w72_12_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid467_Out0_copy468_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid469_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid469_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid469_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_13_c0 :  std_logic;
signal bh7_w73_12_c0 :  std_logic;
signal bh7_w74_12_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid469_Out0_copy470_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid471_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid471_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid471_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_13_c0 :  std_logic;
signal bh7_w75_11_c0 :  std_logic;
signal bh7_w76_11_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid471_Out0_copy472_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid473_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid473_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid473_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_12_c0 :  std_logic;
signal bh7_w77_11_c0 :  std_logic;
signal bh7_w78_11_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid473_Out0_copy474_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid475_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid475_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid475_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_12_c0 :  std_logic;
signal bh7_w79_11_c0 :  std_logic;
signal bh7_w80_11_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid475_Out0_copy476_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid477_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid477_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid477_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_12_c0 :  std_logic;
signal bh7_w81_11_c0 :  std_logic;
signal bh7_w82_11_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid477_Out0_copy478_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid479_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid479_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid479_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_12_c0 :  std_logic;
signal bh7_w83_10_c0 :  std_logic;
signal bh7_w84_10_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid479_Out0_copy480_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid481_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid481_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w83_11_c0 :  std_logic;
signal bh7_w84_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid481_Out0_copy482_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid483_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid483_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w84_12_c0 :  std_logic;
signal bh7_w85_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid483_Out0_copy484_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid485_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid485_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid485_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w85_12_c0 :  std_logic;
signal bh7_w86_9_c0 :  std_logic;
signal bh7_w87_10_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid485_Out0_copy486_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid487_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid487_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w86_10_c0 :  std_logic;
signal bh7_w87_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid487_Out0_copy488_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid489_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid489_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w87_12_c0 :  std_logic;
signal bh7_w88_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid489_Out0_copy490_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid491_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid491_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid491_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w88_12_c0 :  std_logic;
signal bh7_w89_9_c0 :  std_logic;
signal bh7_w90_10_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid491_Out0_copy492_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid493_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid493_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w89_10_c0 :  std_logic;
signal bh7_w90_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid493_Out0_copy494_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid495_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid495_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w90_12_c0 :  std_logic;
signal bh7_w91_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid495_Out0_copy496_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid497_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid497_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid497_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w91_12_c0 :  std_logic;
signal bh7_w92_9_c0 :  std_logic;
signal bh7_w93_10_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid497_Out0_copy498_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid499_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid499_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w92_10_c0 :  std_logic;
signal bh7_w93_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid499_Out0_copy500_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid501_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid501_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w93_12_c0 :  std_logic;
signal bh7_w94_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid501_Out0_copy502_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid503_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid503_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid503_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w94_12_c0 :  std_logic;
signal bh7_w95_9_c0 :  std_logic;
signal bh7_w96_10_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid503_Out0_copy504_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid505_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid505_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w95_10_c0 :  std_logic;
signal bh7_w96_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid505_Out0_copy506_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid507_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid507_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w96_12_c0 :  std_logic;
signal bh7_w97_11_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid507_Out0_copy508_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid509_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid509_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid509_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w97_12_c0 :  std_logic;
signal bh7_w98_9_c0 :  std_logic;
signal bh7_w99_9_c0 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid509_Out0_copy510_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid511_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid511_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w98_10_c0 :  std_logic;
signal bh7_w99_10_c0 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid511_Out0_copy512_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid513_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid513_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid513_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w99_11_c0 :  std_logic;
signal bh7_w100_9_c0 :  std_logic;
signal bh7_w101_6_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid513_Out0_copy514_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid515_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid515_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid515_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w101_7_c0 :  std_logic;
signal bh7_w102_7_c0 :  std_logic;
signal bh7_w103_3_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid515_Out0_copy516_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid517_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid517_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid517_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w103_4_c0 :  std_logic;
signal bh7_w104_2_c0 :  std_logic;
signal bh7_w105_1_c0 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid517_Out0_copy518_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid519_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid519_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w53_14_c1 :  std_logic;
signal bh7_w54_15_c1 :  std_logic;
signal bh7_w55_15_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_copy520_c0, Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_copy520_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid521_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid521_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w55_16_c1 :  std_logic;
signal bh7_w56_14_c1 :  std_logic;
signal bh7_w57_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_copy522_c0, Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_copy522_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid523_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w57_17_c1 :  std_logic;
signal bh7_w58_16_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_copy524_c0, Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_copy524_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid525_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid525_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w58_17_c1 :  std_logic;
signal bh7_w59_14_c1 :  std_logic;
signal bh7_w60_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_copy526_c0, Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_copy526_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid527_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w60_17_c1 :  std_logic;
signal bh7_w61_16_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_copy528_c0, Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_copy528_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid529_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid529_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w61_17_c1 :  std_logic;
signal bh7_w62_14_c1 :  std_logic;
signal bh7_w63_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_copy530_c0, Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_copy530_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid531_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w63_17_c1 :  std_logic;
signal bh7_w64_16_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_copy532_c0, Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_copy532_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid533_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid533_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_17_c1 :  std_logic;
signal bh7_w65_13_c1 :  std_logic;
signal bh7_w66_15_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_copy534_c0, Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_copy534_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid535_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid535_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w66_16_c1 :  std_logic;
signal bh7_w67_14_c1 :  std_logic;
signal bh7_w68_15_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_copy536_c0, Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_copy536_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid537_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid537_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_16_c1 :  std_logic;
signal bh7_w69_13_c1 :  std_logic;
signal bh7_w70_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_copy538_c0, Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_copy538_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid539_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid539_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_15_c1 :  std_logic;
signal bh7_w71_13_c1 :  std_logic;
signal bh7_w72_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_copy540_c0, Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_copy540_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid541_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid541_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_15_c1 :  std_logic;
signal bh7_w73_13_c1 :  std_logic;
signal bh7_w74_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_copy542_c0, Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_copy542_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid543_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid543_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_15_c1 :  std_logic;
signal bh7_w75_12_c1 :  std_logic;
signal bh7_w76_13_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_copy544_c0, Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_copy544_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid545_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid545_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_14_c1 :  std_logic;
signal bh7_w77_12_c1 :  std_logic;
signal bh7_w78_13_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_copy546_c0, Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_copy546_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid547_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid547_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_14_c1 :  std_logic;
signal bh7_w79_12_c1 :  std_logic;
signal bh7_w80_13_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_copy548_c0, Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_copy548_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid549_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid549_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_14_c1 :  std_logic;
signal bh7_w81_12_c1 :  std_logic;
signal bh7_w82_13_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_copy550_c0, Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_copy550_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid551_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid551_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_14_c1 :  std_logic;
signal bh7_w83_12_c1 :  std_logic;
signal bh7_w84_13_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_copy552_c0, Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_copy552_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid553_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid553_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_14_c1 :  std_logic;
signal bh7_w85_13_c1 :  std_logic;
signal bh7_w86_11_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_copy554_c0, Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_copy554_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid555_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w86_12_c1 :  std_logic;
signal bh7_w87_13_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_copy556_c0, Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_copy556_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid557_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid557_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w87_14_c1 :  std_logic;
signal bh7_w88_13_c1 :  std_logic;
signal bh7_w89_11_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_copy558_c0, Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_copy558_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid559_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w89_12_c1 :  std_logic;
signal bh7_w90_13_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_copy560_c0, Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_copy560_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid561_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid561_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w90_14_c1 :  std_logic;
signal bh7_w91_13_c1 :  std_logic;
signal bh7_w92_11_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_copy562_c0, Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_copy562_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid563_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w92_12_c1 :  std_logic;
signal bh7_w93_13_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_copy564_c0, Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_copy564_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid565_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid565_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w93_14_c1 :  std_logic;
signal bh7_w94_13_c1 :  std_logic;
signal bh7_w95_11_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_copy566_c0, Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_copy566_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid567_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w95_12_c1 :  std_logic;
signal bh7_w96_13_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_copy568_c0, Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_copy568_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid569_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid569_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w96_14_c1 :  std_logic;
signal bh7_w97_13_c1 :  std_logic;
signal bh7_w98_11_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_copy570_c0, Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_copy570_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid571_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w98_12_c1 :  std_logic;
signal bh7_w99_12_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_copy572_c0, Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_copy572_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid573_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid573_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w99_13_c1 :  std_logic;
signal bh7_w100_10_c1 :  std_logic;
signal bh7_w101_8_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_copy574_c0, Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_copy574_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid575_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid575_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w101_9_c1 :  std_logic;
signal bh7_w102_8_c1 :  std_logic;
signal bh7_w103_5_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_copy576_c0, Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_copy576_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid577_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid577_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w103_6_c1 :  std_logic;
signal bh7_w104_3_c1 :  std_logic;
signal bh7_w105_2_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_copy578_c0, Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_copy578_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid579_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid579_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w105_3_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid579_Out0_copy580_c0, Compressor_3_2_Freq500_uid432_bh7_uid579_Out0_copy580_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid581_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid581_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid581_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w55_17_c1 :  std_logic;
signal bh7_w56_15_c1 :  std_logic;
signal bh7_w57_18_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid581_Out0_copy582_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid583_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid583_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid583_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w57_19_c1 :  std_logic;
signal bh7_w58_18_c1 :  std_logic;
signal bh7_w59_15_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid583_Out0_copy584_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid585_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid585_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid585_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w60_18_c1 :  std_logic;
signal bh7_w61_18_c1 :  std_logic;
signal bh7_w62_15_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid585_Out0_copy586_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid587_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid587_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid587_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w63_18_c1 :  std_logic;
signal bh7_w64_18_c1 :  std_logic;
signal bh7_w65_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid587_Out0_copy588_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid589_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid589_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid589_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w66_17_c1 :  std_logic;
signal bh7_w67_15_c1 :  std_logic;
signal bh7_w68_17_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid589_Out0_copy590_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid591_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid591_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid591_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_18_c1 :  std_logic;
signal bh7_w69_14_c1 :  std_logic;
signal bh7_w70_16_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid591_Out0_copy592_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid593_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid593_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid593_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_17_c1 :  std_logic;
signal bh7_w71_14_c1 :  std_logic;
signal bh7_w72_16_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid593_Out0_copy594_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid595_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid595_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid595_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_17_c1 :  std_logic;
signal bh7_w73_14_c1 :  std_logic;
signal bh7_w74_16_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid595_Out0_copy596_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid597_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid597_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid597_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_17_c1 :  std_logic;
signal bh7_w75_13_c1 :  std_logic;
signal bh7_w76_15_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid597_Out0_copy598_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid599_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid599_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid599_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_16_c1 :  std_logic;
signal bh7_w77_13_c1 :  std_logic;
signal bh7_w78_15_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid599_Out0_copy600_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid601_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid601_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid601_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_16_c1 :  std_logic;
signal bh7_w79_13_c1 :  std_logic;
signal bh7_w80_15_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid601_Out0_copy602_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid603_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid603_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid603_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_16_c1 :  std_logic;
signal bh7_w81_13_c1 :  std_logic;
signal bh7_w82_15_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid603_Out0_copy604_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid605_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid605_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid605_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_16_c1 :  std_logic;
signal bh7_w83_13_c1 :  std_logic;
signal bh7_w84_15_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid605_Out0_copy606_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid607_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid607_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid607_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_16_c1 :  std_logic;
signal bh7_w85_14_c1 :  std_logic;
signal bh7_w86_13_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid607_Out0_copy608_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid609_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid609_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid609_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_14_c1 :  std_logic;
signal bh7_w87_15_c1 :  std_logic;
signal bh7_w88_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid609_Out0_copy610_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid611_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid611_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid611_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w89_13_c1 :  std_logic;
signal bh7_w90_15_c1 :  std_logic;
signal bh7_w91_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid611_Out0_copy612_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid613_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid613_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid613_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w92_13_c1 :  std_logic;
signal bh7_w93_15_c1 :  std_logic;
signal bh7_w94_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid613_Out0_copy614_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid615_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid615_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid615_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w95_13_c1 :  std_logic;
signal bh7_w96_15_c1 :  std_logic;
signal bh7_w97_14_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid615_Out0_copy616_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid617_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid617_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid617_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w98_13_c1 :  std_logic;
signal bh7_w99_14_c1 :  std_logic;
signal bh7_w100_11_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid617_Out0_copy618_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid619_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid619_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid619_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w101_10_c1 :  std_logic;
signal bh7_w102_9_c1 :  std_logic;
signal bh7_w103_7_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid619_Out0_copy620_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid621_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid621_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid621_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w103_8_c1 :  std_logic;
signal bh7_w104_4_c1 :  std_logic;
signal bh7_w105_4_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid621_Out0_copy622_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid623_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid623_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid623_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid623_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w105_5_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid623_Out0_copy624_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid625_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid625_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid625_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w17_2_c1, bh7_w17_2_c2 :  std_logic;
signal bh7_w18_2_c1, bh7_w18_2_c2 :  std_logic;
signal bh7_w19_2_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid625_Out0_copy626_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid627_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid627_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid627_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w19_3_c1 :  std_logic;
signal bh7_w20_2_c1 :  std_logic;
signal bh7_w21_2_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid627_Out0_copy628_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid629_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid629_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid629_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_3_c1 :  std_logic;
signal bh7_w22_2_c1 :  std_logic;
signal bh7_w23_2_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid629_Out0_copy630_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid631_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid631_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w23_3_c1 :  std_logic;
signal bh7_w24_3_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid631_Out0_copy632_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid633_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid633_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid633_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w24_4_c1 :  std_logic;
signal bh7_w25_3_c1 :  std_logic;
signal bh7_w26_3_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid633_Out0_copy634_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid635_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid635_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid635_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w26_4_c1 :  std_logic;
signal bh7_w27_3_c1 :  std_logic;
signal bh7_w28_3_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid635_Out0_copy636_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid637_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid637_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid637_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w28_4_c1 :  std_logic;
signal bh7_w29_3_c1 :  std_logic;
signal bh7_w30_3_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid637_Out0_copy638_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid639_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid639_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid639_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w30_4_c1 :  std_logic;
signal bh7_w31_3_c1 :  std_logic;
signal bh7_w32_3_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid639_Out0_copy640_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid641_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid641_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid641_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w32_4_c1 :  std_logic;
signal bh7_w33_3_c1 :  std_logic;
signal bh7_w34_4_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid641_Out0_copy642_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid643_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid643_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid643_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w34_5_c1 :  std_logic;
signal bh7_w35_4_c1 :  std_logic;
signal bh7_w36_4_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid643_Out0_copy644_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid645_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid645_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w35_5_c1 :  std_logic;
signal bh7_w36_5_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid645_Out0_copy646_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid647_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid647_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid647_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w36_6_c1 :  std_logic;
signal bh7_w37_4_c1 :  std_logic;
signal bh7_w38_4_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid647_Out0_copy648_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid649_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid649_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w37_5_c1 :  std_logic;
signal bh7_w38_5_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid649_Out0_copy650_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid651_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid651_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid651_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w38_6_c1 :  std_logic;
signal bh7_w39_4_c1 :  std_logic;
signal bh7_w40_4_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid651_Out0_copy652_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid653_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid653_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w39_5_c1 :  std_logic;
signal bh7_w40_5_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid653_Out0_copy654_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid655_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid655_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid655_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w40_6_c1 :  std_logic;
signal bh7_w41_4_c1 :  std_logic;
signal bh7_w42_4_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid655_Out0_copy656_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid657_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid657_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w41_5_c1 :  std_logic;
signal bh7_w42_5_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid657_Out0_copy658_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid659_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid659_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid659_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w42_6_c1 :  std_logic;
signal bh7_w43_4_c1 :  std_logic;
signal bh7_w44_4_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid659_Out0_copy660_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid661_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid661_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w43_5_c1 :  std_logic;
signal bh7_w44_5_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid661_Out0_copy662_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid663_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid663_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid663_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w44_6_c1 :  std_logic;
signal bh7_w45_4_c1 :  std_logic;
signal bh7_w46_4_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid663_Out0_copy664_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid665_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid665_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w45_5_c1 :  std_logic;
signal bh7_w46_5_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid665_Out0_copy666_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid667_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid667_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid667_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w46_6_c1 :  std_logic;
signal bh7_w47_4_c1 :  std_logic;
signal bh7_w48_5_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid667_Out0_copy668_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid669_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid669_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w47_5_c1 :  std_logic;
signal bh7_w48_6_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid669_Out0_copy670_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid671_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid671_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid671_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid671_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w48_7_c1 :  std_logic;
signal bh7_w49_6_c1, bh7_w49_6_c2 :  std_logic;
signal bh7_w50_7_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid671_Out0_copy672_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid673_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid673_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid673_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid673_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w49_7_c1 :  std_logic;
signal bh7_w50_8_c1 :  std_logic;
signal bh7_w51_11_c1, bh7_w51_11_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid673_Out0_copy674_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid675_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid675_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid675_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid675_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w50_9_c1 :  std_logic;
signal bh7_w51_12_c1 :  std_logic;
signal bh7_w52_12_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid675_Out0_copy676_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid677_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid677_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid677_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid677_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w51_13_c1 :  std_logic;
signal bh7_w52_13_c1 :  std_logic;
signal bh7_w53_15_c1, bh7_w53_15_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid677_Out0_copy678_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid679_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid679_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid679_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w52_14_c1 :  std_logic;
signal bh7_w53_16_c1 :  std_logic;
signal bh7_w54_16_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid679_Out0_copy680_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid681_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid681_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid681_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w53_17_c1 :  std_logic;
signal bh7_w54_17_c1 :  std_logic;
signal bh7_w55_18_c1, bh7_w55_18_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid681_Out0_copy682_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid683_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid683_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid683_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w54_18_c1 :  std_logic;
signal bh7_w55_19_c1 :  std_logic;
signal bh7_w56_16_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid683_Out0_copy684_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid685_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid685_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid685_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w55_20_c1 :  std_logic;
signal bh7_w56_17_c1 :  std_logic;
signal bh7_w57_20_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid685_Out0_copy686_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid687_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid687_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w56_18_c1 :  std_logic;
signal bh7_w57_21_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid687_Out0_copy688_c1 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid689_In0_c1 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid689_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w57_22_c1 :  std_logic;
signal bh7_w58_19_c1 :  std_logic;
signal bh7_w59_16_c1 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid689_Out0_copy690_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid691_In0_c1 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq500_uid400_bh7_uid691_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w58_20_c1 :  std_logic;
signal bh7_w59_17_c1 :  std_logic;
signal bh7_w60_19_c1 :  std_logic;
signal Compressor_5_3_Freq500_uid400_bh7_uid691_Out0_copy692_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid693_In0_c1 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid693_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_18_c1 :  std_logic;
signal bh7_w60_20_c1 :  std_logic;
signal bh7_w61_19_c1 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid693_Out0_copy694_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid695_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid695_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid695_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w60_21_c1 :  std_logic;
signal bh7_w61_20_c1 :  std_logic;
signal bh7_w62_16_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid695_Out0_copy696_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid697_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid697_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w61_21_c1 :  std_logic;
signal bh7_w62_17_c1, bh7_w62_17_c2 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid697_Out0_copy698_c1 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid699_In0_c1 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq500_uid334_bh7_uid699_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_18_c1 :  std_logic;
signal bh7_w63_19_c1 :  std_logic;
signal bh7_w64_19_c1 :  std_logic;
signal Compressor_6_3_Freq500_uid334_bh7_uid699_Out0_copy700_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid701_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid701_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid701_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w63_20_c1 :  std_logic;
signal bh7_w64_20_c1 :  std_logic;
signal bh7_w65_15_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid701_Out0_copy702_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid703_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid703_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid703_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_21_c1, bh7_w64_21_c2 :  std_logic;
signal bh7_w65_16_c1 :  std_logic;
signal bh7_w66_18_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid703_Out0_copy704_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid705_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid705_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid705_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w65_17_c1 :  std_logic;
signal bh7_w66_19_c1 :  std_logic;
signal bh7_w67_16_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid705_Out0_copy706_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid707_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid707_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w66_20_c1, bh7_w66_20_c2 :  std_logic;
signal bh7_w67_17_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid707_Out0_copy708_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid709_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid709_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid709_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w67_18_c1 :  std_logic;
signal bh7_w68_19_c1 :  std_logic;
signal bh7_w69_15_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid709_Out0_copy710_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid711_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid711_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid711_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_20_c1 :  std_logic;
signal bh7_w69_16_c1 :  std_logic;
signal bh7_w70_18_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid711_Out0_copy712_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid713_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid713_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w69_17_c1 :  std_logic;
signal bh7_w70_19_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid713_Out0_copy714_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid715_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid715_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid715_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_20_c1 :  std_logic;
signal bh7_w71_15_c1 :  std_logic;
signal bh7_w72_18_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid715_Out0_copy716_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid717_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid717_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w71_16_c1, bh7_w71_16_c2 :  std_logic;
signal bh7_w72_19_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid717_Out0_copy718_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid719_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid719_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid719_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_20_c1 :  std_logic;
signal bh7_w73_15_c1 :  std_logic;
signal bh7_w74_18_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid719_Out0_copy720_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid721_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid721_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w73_16_c1, bh7_w73_16_c2 :  std_logic;
signal bh7_w74_19_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid721_Out0_copy722_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid723_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid723_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid723_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_20_c1 :  std_logic;
signal bh7_w75_14_c1 :  std_logic;
signal bh7_w76_17_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid723_Out0_copy724_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid725_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid725_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid725_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_21_c1 :  std_logic;
signal bh7_w75_15_c1, bh7_w75_15_c2 :  std_logic;
signal bh7_w76_18_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid725_Out0_copy726_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid727_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid727_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid727_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid727_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_19_c1 :  std_logic;
signal bh7_w77_14_c1 :  std_logic;
signal bh7_w78_17_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid727_Out0_copy728_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid729_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid729_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w77_15_c1 :  std_logic;
signal bh7_w78_18_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid729_Out0_copy730_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid731_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid731_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid731_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid731_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_19_c1 :  std_logic;
signal bh7_w79_14_c1 :  std_logic;
signal bh7_w80_17_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid731_Out0_copy732_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid733_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid733_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w79_15_c1 :  std_logic;
signal bh7_w80_18_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid733_Out0_copy734_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid735_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid735_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid735_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid735_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_19_c1 :  std_logic;
signal bh7_w81_14_c1 :  std_logic;
signal bh7_w82_17_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid735_Out0_copy736_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid737_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid737_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w81_15_c1 :  std_logic;
signal bh7_w82_18_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid737_Out0_copy738_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid739_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid739_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid739_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_19_c1 :  std_logic;
signal bh7_w83_14_c1, bh7_w83_14_c2 :  std_logic;
signal bh7_w84_17_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid739_Out0_copy740_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid741_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid741_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid741_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_18_c1 :  std_logic;
signal bh7_w85_15_c1 :  std_logic;
signal bh7_w86_15_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid741_Out0_copy742_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid743_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid743_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid743_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_16_c1 :  std_logic;
signal bh7_w87_16_c1 :  std_logic;
signal bh7_w88_15_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid743_Out0_copy744_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid745_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid745_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid745_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_16_c1 :  std_logic;
signal bh7_w89_14_c1 :  std_logic;
signal bh7_w90_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid745_Out0_copy746_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid747_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid747_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w90_17_c1 :  std_logic;
signal bh7_w91_15_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid747_Out0_copy748_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid749_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid749_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid749_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w91_16_c1 :  std_logic;
signal bh7_w92_14_c1, bh7_w92_14_c2 :  std_logic;
signal bh7_w93_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid749_Out0_copy750_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid751_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid751_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w93_17_c1 :  std_logic;
signal bh7_w94_15_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid751_Out0_copy752_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid753_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid753_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid753_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w94_16_c1 :  std_logic;
signal bh7_w95_14_c1, bh7_w95_14_c2 :  std_logic;
signal bh7_w96_16_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid753_Out0_copy754_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid755_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid755_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w96_17_c1 :  std_logic;
signal bh7_w97_15_c1 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid755_Out0_copy756_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid757_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid757_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid757_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w97_16_c1 :  std_logic;
signal bh7_w98_14_c1, bh7_w98_14_c2 :  std_logic;
signal bh7_w99_15_c1 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid757_Out0_copy758_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid759_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid759_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid759_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w100_12_c1 :  std_logic;
signal bh7_w101_11_c1, bh7_w101_11_c2 :  std_logic;
signal bh7_w102_10_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid759_Out0_copy760_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid761_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid761_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid761_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w103_9_c1 :  std_logic;
signal bh7_w104_5_c1, bh7_w104_5_c2 :  std_logic;
signal bh7_w105_6_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid761_Out0_copy762_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid763_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid763_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid763_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid763_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w105_7_c1 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid763_Out0_copy764_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid765_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid765_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w19_4_c2 :  std_logic;
signal bh7_w20_3_c2 :  std_logic;
signal bh7_w21_4_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_copy766_c1, Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_copy766_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid767_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid767_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w21_5_c2 :  std_logic;
signal bh7_w22_3_c2 :  std_logic;
signal bh7_w23_4_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_copy768_c1, Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_copy768_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid769_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid769_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w23_5_c2 :  std_logic;
signal bh7_w24_5_c2 :  std_logic;
signal bh7_w25_4_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_copy770_c1, Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_copy770_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid771_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid771_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w25_5_c2 :  std_logic;
signal bh7_w26_5_c2 :  std_logic;
signal bh7_w27_4_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_copy772_c1, Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_copy772_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid773_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid773_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w27_5_c2 :  std_logic;
signal bh7_w28_5_c2 :  std_logic;
signal bh7_w29_4_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_copy774_c1, Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_copy774_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid775_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid775_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w29_5_c2 :  std_logic;
signal bh7_w30_5_c2 :  std_logic;
signal bh7_w31_4_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_copy776_c1, Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_copy776_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid777_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid777_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w31_5_c2 :  std_logic;
signal bh7_w32_5_c2 :  std_logic;
signal bh7_w33_4_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_copy778_c1, Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_copy778_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid779_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid779_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w33_5_c2 :  std_logic;
signal bh7_w34_6_c2 :  std_logic;
signal bh7_w35_6_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_copy780_c1, Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_copy780_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid781_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w35_7_c2 :  std_logic;
signal bh7_w36_7_c2 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_copy782_c1, Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_copy782_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid783_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid783_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w36_8_c2 :  std_logic;
signal bh7_w37_6_c2 :  std_logic;
signal bh7_w38_7_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_copy784_c1, Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_copy784_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid785_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid785_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w38_8_c2 :  std_logic;
signal bh7_w39_6_c2 :  std_logic;
signal bh7_w40_7_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_copy786_c1, Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_copy786_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid787_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid787_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w40_8_c2 :  std_logic;
signal bh7_w41_6_c2 :  std_logic;
signal bh7_w42_7_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_copy788_c1, Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_copy788_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid789_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid789_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w42_8_c2 :  std_logic;
signal bh7_w43_6_c2 :  std_logic;
signal bh7_w44_7_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_copy790_c1, Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_copy790_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid791_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid791_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w44_8_c2 :  std_logic;
signal bh7_w45_6_c2 :  std_logic;
signal bh7_w46_7_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_copy792_c1, Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_copy792_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid793_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid793_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w46_8_c2 :  std_logic;
signal bh7_w47_6_c2 :  std_logic;
signal bh7_w48_8_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_copy794_c1, Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_copy794_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid795_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid795_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w48_9_c2 :  std_logic;
signal bh7_w49_8_c2 :  std_logic;
signal bh7_w50_10_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_copy796_c1, Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_copy796_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid797_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid797_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w50_11_c2 :  std_logic;
signal bh7_w51_14_c2 :  std_logic;
signal bh7_w52_15_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_copy798_c1, Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_copy798_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid799_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid799_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w52_16_c2 :  std_logic;
signal bh7_w53_18_c2 :  std_logic;
signal bh7_w54_19_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_copy800_c1, Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_copy800_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid801_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid801_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w54_20_c2 :  std_logic;
signal bh7_w55_21_c2 :  std_logic;
signal bh7_w56_19_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_copy802_c1, Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_copy802_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid803_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid803_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid803_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w56_20_c2 :  std_logic;
signal bh7_w57_23_c2 :  std_logic;
signal bh7_w58_21_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_copy804_c1, Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_copy804_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid805_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid805_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w57_24_c2 :  std_logic;
signal bh7_w58_22_c2 :  std_logic;
signal bh7_w59_19_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_copy806_c1, Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_copy806_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid807_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w59_20_c2 :  std_logic;
signal bh7_w60_22_c2 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_copy808_c1, Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_copy808_c2 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid809_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid809_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w60_23_c2 :  std_logic;
signal bh7_w61_22_c2 :  std_logic;
signal bh7_w62_19_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_copy810_c1, Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_copy810_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid811_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid811_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w61_23_c2 :  std_logic;
signal bh7_w62_20_c2 :  std_logic;
signal bh7_w63_21_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_copy812_c1, Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_copy812_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid813_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid813_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w63_22_c2 :  std_logic;
signal bh7_w64_22_c2 :  std_logic;
signal bh7_w65_18_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_copy814_c1, Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_copy814_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid815_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid815_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w65_19_c2 :  std_logic;
signal bh7_w66_21_c2 :  std_logic;
signal bh7_w67_19_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_copy816_c1, Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_copy816_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid817_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid817_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w67_20_c2 :  std_logic;
signal bh7_w68_21_c2 :  std_logic;
signal bh7_w69_18_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_copy818_c1, Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_copy818_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid819_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w69_19_c2 :  std_logic;
signal bh7_w70_21_c2 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_copy820_c1, Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_copy820_c2 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid821_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid821_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w70_22_c2 :  std_logic;
signal bh7_w71_17_c2 :  std_logic;
signal bh7_w72_21_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_copy822_c1, Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_copy822_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid823_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid823_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w72_22_c2 :  std_logic;
signal bh7_w73_17_c2 :  std_logic;
signal bh7_w74_22_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_copy824_c1, Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_copy824_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid825_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid825_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w74_23_c2 :  std_logic;
signal bh7_w75_16_c2 :  std_logic;
signal bh7_w76_20_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_copy826_c1, Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_copy826_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid827_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid827_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w76_21_c2 :  std_logic;
signal bh7_w77_16_c2 :  std_logic;
signal bh7_w78_20_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_copy828_c1, Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_copy828_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid829_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid829_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w78_21_c2 :  std_logic;
signal bh7_w79_16_c2 :  std_logic;
signal bh7_w80_20_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_copy830_c1, Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_copy830_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid831_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid831_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w80_21_c2 :  std_logic;
signal bh7_w81_16_c2 :  std_logic;
signal bh7_w82_20_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_copy832_c1, Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_copy832_c2 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid833_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_c2 :  std_logic_vector(1 downto 0);
signal bh7_w82_21_c2 :  std_logic;
signal bh7_w83_15_c2 :  std_logic;
signal Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_copy834_c1, Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_copy834_c2 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid835_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid835_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w84_19_c2 :  std_logic;
signal bh7_w85_16_c2 :  std_logic;
signal bh7_w86_17_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_copy836_c1, Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_copy836_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid837_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid837_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w86_18_c2 :  std_logic;
signal bh7_w87_17_c2 :  std_logic;
signal bh7_w88_17_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_copy838_c1, Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_copy838_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid839_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid839_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w88_18_c2 :  std_logic;
signal bh7_w89_15_c2 :  std_logic;
signal bh7_w90_18_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_copy840_c1, Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_copy840_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid841_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid841_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w90_19_c2 :  std_logic;
signal bh7_w91_17_c2 :  std_logic;
signal bh7_w92_15_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_copy842_c1, Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_copy842_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid843_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid843_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w93_18_c2 :  std_logic;
signal bh7_w94_17_c2 :  std_logic;
signal bh7_w95_15_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_copy844_c1, Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_copy844_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid845_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid845_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w96_18_c2 :  std_logic;
signal bh7_w97_17_c2 :  std_logic;
signal bh7_w98_15_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_copy846_c1, Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_copy846_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid847_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid847_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w99_16_c2 :  std_logic;
signal bh7_w100_13_c2 :  std_logic;
signal bh7_w101_12_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_copy848_c1, Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_copy848_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid849_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid849_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w102_11_c2 :  std_logic;
signal bh7_w103_10_c2 :  std_logic;
signal bh7_w104_6_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_copy850_c1, Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_copy850_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid851_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid851_In1_c0, Compressor_14_3_Freq500_uid326_bh7_uid851_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid851_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w105_8_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid851_Out0_copy852_c1, Compressor_14_3_Freq500_uid326_bh7_uid851_Out0_copy852_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid853_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid853_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid853_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w21_6_c2 :  std_logic;
signal bh7_w22_4_c2 :  std_logic;
signal bh7_w23_6_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid853_Out0_copy854_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid855_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid855_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid855_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w23_7_c2 :  std_logic;
signal bh7_w24_6_c2 :  std_logic;
signal bh7_w25_6_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid855_Out0_copy856_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid857_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid857_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid857_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w25_7_c2 :  std_logic;
signal bh7_w26_6_c2 :  std_logic;
signal bh7_w27_6_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid857_Out0_copy858_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid859_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid859_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid859_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w27_7_c2 :  std_logic;
signal bh7_w28_6_c2 :  std_logic;
signal bh7_w29_6_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid859_Out0_copy860_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid861_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid861_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid861_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w29_7_c2 :  std_logic;
signal bh7_w30_6_c2 :  std_logic;
signal bh7_w31_6_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid861_Out0_copy862_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid863_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid863_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid863_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w31_7_c2 :  std_logic;
signal bh7_w32_6_c2 :  std_logic;
signal bh7_w33_6_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid863_Out0_copy864_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid865_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid865_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid865_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w33_7_c2 :  std_logic;
signal bh7_w34_7_c2 :  std_logic;
signal bh7_w35_8_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid865_Out0_copy866_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid867_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid867_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid867_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w35_9_c2 :  std_logic;
signal bh7_w36_9_c2 :  std_logic;
signal bh7_w37_7_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid867_Out0_copy868_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid869_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid869_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid869_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w38_9_c2 :  std_logic;
signal bh7_w39_7_c2 :  std_logic;
signal bh7_w40_9_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid869_Out0_copy870_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid871_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid871_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid871_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w40_10_c2 :  std_logic;
signal bh7_w41_7_c2 :  std_logic;
signal bh7_w42_9_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid871_Out0_copy872_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid873_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid873_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid873_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w42_10_c2 :  std_logic;
signal bh7_w43_7_c2 :  std_logic;
signal bh7_w44_9_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid873_Out0_copy874_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid875_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid875_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid875_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w44_10_c2 :  std_logic;
signal bh7_w45_7_c2 :  std_logic;
signal bh7_w46_9_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid875_Out0_copy876_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid877_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid877_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid877_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w46_10_c2 :  std_logic;
signal bh7_w47_7_c2 :  std_logic;
signal bh7_w48_10_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid877_Out0_copy878_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid879_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid879_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid879_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w48_11_c2 :  std_logic;
signal bh7_w49_9_c2 :  std_logic;
signal bh7_w50_12_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid879_Out0_copy880_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid881_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid881_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid881_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w50_13_c2 :  std_logic;
signal bh7_w51_15_c2 :  std_logic;
signal bh7_w52_17_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid881_Out0_copy882_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid883_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid883_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid883_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w52_18_c2 :  std_logic;
signal bh7_w53_19_c2 :  std_logic;
signal bh7_w54_21_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid883_Out0_copy884_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid885_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid885_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid885_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w54_22_c2 :  std_logic;
signal bh7_w55_22_c2 :  std_logic;
signal bh7_w56_21_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid885_Out0_copy886_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid887_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid887_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid887_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w56_22_c2 :  std_logic;
signal bh7_w57_25_c2 :  std_logic;
signal bh7_w58_23_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid887_Out0_copy888_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid889_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid889_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid889_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w58_24_c2 :  std_logic;
signal bh7_w59_21_c2 :  std_logic;
signal bh7_w60_24_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid889_Out0_copy890_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid891_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid891_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid891_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w60_25_c2 :  std_logic;
signal bh7_w61_24_c2 :  std_logic;
signal bh7_w62_21_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid891_Out0_copy892_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid893_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid893_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid893_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w62_22_c2 :  std_logic;
signal bh7_w63_23_c2 :  std_logic;
signal bh7_w64_23_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid893_Out0_copy894_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid895_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid895_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid895_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w64_24_c2 :  std_logic;
signal bh7_w65_20_c2 :  std_logic;
signal bh7_w66_22_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid895_Out0_copy896_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid897_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid897_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid897_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w66_23_c2 :  std_logic;
signal bh7_w67_21_c2 :  std_logic;
signal bh7_w68_22_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid897_Out0_copy898_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid899_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid899_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid899_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w69_20_c2 :  std_logic;
signal bh7_w70_23_c2 :  std_logic;
signal bh7_w71_18_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid899_Out0_copy900_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid901_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid901_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid901_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w71_19_c2 :  std_logic;
signal bh7_w72_23_c2 :  std_logic;
signal bh7_w73_18_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid901_Out0_copy902_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid903_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid903_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid903_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w73_19_c2 :  std_logic;
signal bh7_w74_24_c2 :  std_logic;
signal bh7_w75_17_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid903_Out0_copy904_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid905_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid905_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid905_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w75_18_c2 :  std_logic;
signal bh7_w76_22_c2 :  std_logic;
signal bh7_w77_17_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid905_Out0_copy906_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid907_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid907_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid907_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w78_22_c2 :  std_logic;
signal bh7_w79_17_c2 :  std_logic;
signal bh7_w80_22_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid907_Out0_copy908_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid909_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid909_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid909_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w80_23_c2 :  std_logic;
signal bh7_w81_17_c2 :  std_logic;
signal bh7_w82_22_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid909_Out0_copy910_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid911_In0_c2 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid911_In1_c2 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq500_uid322_bh7_uid911_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w82_23_c2 :  std_logic;
signal bh7_w83_16_c2 :  std_logic;
signal bh7_w84_20_c2 :  std_logic;
signal Compressor_23_3_Freq500_uid322_bh7_uid911_Out0_copy912_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid913_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid913_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid913_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w86_19_c2 :  std_logic;
signal bh7_w87_18_c2 :  std_logic;
signal bh7_w88_19_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid913_Out0_copy914_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid915_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid915_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid915_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w88_20_c2 :  std_logic;
signal bh7_w89_16_c2 :  std_logic;
signal bh7_w90_20_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid915_Out0_copy916_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid917_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid917_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid917_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w90_21_c2 :  std_logic;
signal bh7_w91_18_c2 :  std_logic;
signal bh7_w92_16_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid917_Out0_copy918_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid919_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid919_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid919_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w92_17_c2 :  std_logic;
signal bh7_w93_19_c2 :  std_logic;
signal bh7_w94_18_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid919_Out0_copy920_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid921_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid921_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid921_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w95_16_c2 :  std_logic;
signal bh7_w96_19_c2 :  std_logic;
signal bh7_w97_18_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid921_Out0_copy922_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid923_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid923_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid923_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w98_16_c2 :  std_logic;
signal bh7_w99_17_c2 :  std_logic;
signal bh7_w100_14_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid923_Out0_copy924_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid925_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid925_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid925_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w101_13_c2 :  std_logic;
signal bh7_w102_12_c2 :  std_logic;
signal bh7_w103_11_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid925_Out0_copy926_c2 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid927_In0_c2 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid927_In1_c2 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq500_uid326_bh7_uid927_Out0_c2 :  std_logic_vector(2 downto 0);
signal bh7_w104_7_c2 :  std_logic;
signal bh7_w105_9_c2 :  std_logic;
signal Compressor_14_3_Freq500_uid326_bh7_uid927_Out0_copy928_c2 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh7_22_c2, tmp_bitheapResult_bh7_22_c3, tmp_bitheapResult_bh7_22_c4 :  std_logic_vector(22 downto 0);
signal bitheapFinalAdd_bh7_In0_c2 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_In1_c2 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh7_Out_c4 :  std_logic_vector(83 downto 0);
signal bitheapResult_bh7_c4 :  std_logic_vector(105 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               bh7_w48_4_c1 <= bh7_w48_4_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_copy520_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_copy520_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_copy522_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_copy522_c0;
               Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_copy524_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_copy524_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_copy526_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_copy526_c0;
               Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_copy528_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_copy528_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_copy530_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_copy530_c0;
               Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_copy532_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_copy532_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_copy534_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_copy534_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_copy536_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_copy536_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_copy538_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_copy538_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_copy540_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_copy540_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_copy542_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_copy542_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_copy544_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_copy544_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_copy546_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_copy546_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_copy548_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_copy548_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_copy550_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_copy550_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_copy552_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_copy552_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_copy554_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_copy554_c0;
               Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_copy556_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_copy556_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_copy558_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_copy558_c0;
               Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_copy560_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_copy560_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_copy562_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_copy562_c0;
               Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_copy564_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_copy564_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_copy566_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_copy566_c0;
               Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_copy568_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_copy568_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_copy570_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_copy570_c0;
               Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_copy572_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_copy572_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_copy574_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_copy574_c0;
               Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_copy576_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_copy576_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_copy578_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_copy578_c0;
               Compressor_3_2_Freq500_uid432_bh7_uid579_Out0_copy580_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid579_Out0_copy580_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid623_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid623_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid671_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid671_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid673_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid673_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid675_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid675_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid677_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid677_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid727_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid727_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid731_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid731_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid735_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid735_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid763_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid763_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid803_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid803_In1_c0;
               Compressor_14_3_Freq500_uid326_bh7_uid851_In1_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid851_In1_c0;
            end if;
            if ce_2 = '1' then
               bh7_w0_0_c2 <= bh7_w0_0_c1;
               bh7_w1_0_c2 <= bh7_w1_0_c1;
               bh7_w2_0_c2 <= bh7_w2_0_c1;
               bh7_w3_0_c2 <= bh7_w3_0_c1;
               bh7_w4_0_c2 <= bh7_w4_0_c1;
               bh7_w5_0_c2 <= bh7_w5_0_c1;
               bh7_w6_0_c2 <= bh7_w6_0_c1;
               bh7_w7_0_c2 <= bh7_w7_0_c1;
               bh7_w8_0_c2 <= bh7_w8_0_c1;
               bh7_w9_0_c2 <= bh7_w9_0_c1;
               bh7_w10_0_c2 <= bh7_w10_0_c1;
               bh7_w11_0_c2 <= bh7_w11_0_c1;
               bh7_w12_0_c2 <= bh7_w12_0_c1;
               bh7_w13_0_c2 <= bh7_w13_0_c1;
               bh7_w14_0_c2 <= bh7_w14_0_c1;
               bh7_w15_0_c2 <= bh7_w15_0_c1;
               bh7_w16_0_c2 <= bh7_w16_0_c1;
               bh7_w17_2_c2 <= bh7_w17_2_c1;
               bh7_w18_2_c2 <= bh7_w18_2_c1;
               bh7_w49_6_c2 <= bh7_w49_6_c1;
               bh7_w51_11_c2 <= bh7_w51_11_c1;
               bh7_w53_15_c2 <= bh7_w53_15_c1;
               bh7_w55_18_c2 <= bh7_w55_18_c1;
               bh7_w62_17_c2 <= bh7_w62_17_c1;
               bh7_w64_21_c2 <= bh7_w64_21_c1;
               bh7_w66_20_c2 <= bh7_w66_20_c1;
               bh7_w71_16_c2 <= bh7_w71_16_c1;
               bh7_w73_16_c2 <= bh7_w73_16_c1;
               bh7_w75_15_c2 <= bh7_w75_15_c1;
               bh7_w83_14_c2 <= bh7_w83_14_c1;
               bh7_w92_14_c2 <= bh7_w92_14_c1;
               bh7_w95_14_c2 <= bh7_w95_14_c1;
               bh7_w98_14_c2 <= bh7_w98_14_c1;
               bh7_w101_11_c2 <= bh7_w101_11_c1;
               bh7_w104_5_c2 <= bh7_w104_5_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_copy766_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_copy766_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_copy768_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_copy768_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_copy770_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_copy770_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_copy772_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_copy772_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_copy774_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_copy774_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_copy776_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_copy776_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_copy778_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_copy778_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_copy780_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_copy780_c1;
               Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_copy782_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_copy782_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_copy784_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_copy784_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_copy786_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_copy786_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_copy788_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_copy788_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_copy790_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_copy790_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_copy792_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_copy792_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_copy794_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_copy794_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_copy796_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_copy796_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_copy798_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_copy798_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_copy800_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_copy800_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_copy802_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_copy802_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_copy804_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_copy804_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_copy806_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_copy806_c1;
               Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_copy808_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_copy808_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_copy810_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_copy810_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_copy812_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_copy812_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_copy814_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_copy814_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_copy816_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_copy816_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_copy818_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_copy818_c1;
               Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_copy820_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_copy820_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_copy822_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_copy822_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_copy824_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_copy824_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_copy826_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_copy826_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_copy828_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_copy828_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_copy830_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_copy830_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_copy832_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_copy832_c1;
               Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_copy834_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_copy834_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_copy836_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_copy836_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_copy838_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_copy838_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_copy840_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_copy840_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_copy842_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_copy842_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_copy844_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_copy844_c1;
               Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_copy846_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_copy846_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_copy848_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_copy848_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_copy850_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_copy850_c1;
               Compressor_14_3_Freq500_uid326_bh7_uid851_Out0_copy852_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid851_Out0_copy852_c1;
            end if;
            if ce_3 = '1' then
               tmp_bitheapResult_bh7_22_c3 <= tmp_bitheapResult_bh7_22_c2;
            end if;
            if ce_4 = '1' then
               tmp_bitheapResult_bh7_22_c4 <= tmp_bitheapResult_bh7_22_c3;
            end if;
         end if;
      end process;
   XX_m6_c0 <= X ;
   YY_m6_c0 <= Y ;
   tile_0_X_c0 <= X(16 downto 0);
   tile_0_Y_c0 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq500_uid9
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 X => tile_0_X_c0,
                 Y => tile_0_Y_c0,
                 R => tile_0_output_c1);

   tile_0_filtered_output_c1 <= unsigned(tile_0_output_c1(40 downto 0));
   bh7_w0_0_c1 <= tile_0_filtered_output_c1(0);
   bh7_w1_0_c1 <= tile_0_filtered_output_c1(1);
   bh7_w2_0_c1 <= tile_0_filtered_output_c1(2);
   bh7_w3_0_c1 <= tile_0_filtered_output_c1(3);
   bh7_w4_0_c1 <= tile_0_filtered_output_c1(4);
   bh7_w5_0_c1 <= tile_0_filtered_output_c1(5);
   bh7_w6_0_c1 <= tile_0_filtered_output_c1(6);
   bh7_w7_0_c1 <= tile_0_filtered_output_c1(7);
   bh7_w8_0_c1 <= tile_0_filtered_output_c1(8);
   bh7_w9_0_c1 <= tile_0_filtered_output_c1(9);
   bh7_w10_0_c1 <= tile_0_filtered_output_c1(10);
   bh7_w11_0_c1 <= tile_0_filtered_output_c1(11);
   bh7_w12_0_c1 <= tile_0_filtered_output_c1(12);
   bh7_w13_0_c1 <= tile_0_filtered_output_c1(13);
   bh7_w14_0_c1 <= tile_0_filtered_output_c1(14);
   bh7_w15_0_c1 <= tile_0_filtered_output_c1(15);
   bh7_w16_0_c1 <= tile_0_filtered_output_c1(16);
   bh7_w17_0_c1 <= tile_0_filtered_output_c1(17);
   bh7_w18_0_c1 <= tile_0_filtered_output_c1(18);
   bh7_w19_0_c1 <= tile_0_filtered_output_c1(19);
   bh7_w20_0_c1 <= tile_0_filtered_output_c1(20);
   bh7_w21_0_c1 <= tile_0_filtered_output_c1(21);
   bh7_w22_0_c1 <= tile_0_filtered_output_c1(22);
   bh7_w23_0_c1 <= tile_0_filtered_output_c1(23);
   bh7_w24_0_c1 <= tile_0_filtered_output_c1(24);
   bh7_w25_0_c1 <= tile_0_filtered_output_c1(25);
   bh7_w26_0_c1 <= tile_0_filtered_output_c1(26);
   bh7_w27_0_c1 <= tile_0_filtered_output_c1(27);
   bh7_w28_0_c1 <= tile_0_filtered_output_c1(28);
   bh7_w29_0_c1 <= tile_0_filtered_output_c1(29);
   bh7_w30_0_c1 <= tile_0_filtered_output_c1(30);
   bh7_w31_0_c1 <= tile_0_filtered_output_c1(31);
   bh7_w32_0_c1 <= tile_0_filtered_output_c1(32);
   bh7_w33_0_c1 <= tile_0_filtered_output_c1(33);
   bh7_w34_0_c1 <= tile_0_filtered_output_c1(34);
   bh7_w35_0_c1 <= tile_0_filtered_output_c1(35);
   bh7_w36_0_c1 <= tile_0_filtered_output_c1(36);
   bh7_w37_0_c1 <= tile_0_filtered_output_c1(37);
   bh7_w38_0_c1 <= tile_0_filtered_output_c1(38);
   bh7_w39_0_c1 <= tile_0_filtered_output_c1(39);
   bh7_w40_0_c1 <= tile_0_filtered_output_c1(40);
   tile_1_X_c0 <= X(33 downto 17);
   tile_1_Y_c0 <= Y(23 downto 0);
   tile_1_mult: DSPBlock_17x24_Freq500_uid11
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 X => tile_1_X_c0,
                 Y => tile_1_Y_c0,
                 R => tile_1_output_c1);

   tile_1_filtered_output_c1 <= unsigned(tile_1_output_c1(40 downto 0));
   bh7_w17_1_c1 <= tile_1_filtered_output_c1(0);
   bh7_w18_1_c1 <= tile_1_filtered_output_c1(1);
   bh7_w19_1_c1 <= tile_1_filtered_output_c1(2);
   bh7_w20_1_c1 <= tile_1_filtered_output_c1(3);
   bh7_w21_1_c1 <= tile_1_filtered_output_c1(4);
   bh7_w22_1_c1 <= tile_1_filtered_output_c1(5);
   bh7_w23_1_c1 <= tile_1_filtered_output_c1(6);
   bh7_w24_1_c1 <= tile_1_filtered_output_c1(7);
   bh7_w25_1_c1 <= tile_1_filtered_output_c1(8);
   bh7_w26_1_c1 <= tile_1_filtered_output_c1(9);
   bh7_w27_1_c1 <= tile_1_filtered_output_c1(10);
   bh7_w28_1_c1 <= tile_1_filtered_output_c1(11);
   bh7_w29_1_c1 <= tile_1_filtered_output_c1(12);
   bh7_w30_1_c1 <= tile_1_filtered_output_c1(13);
   bh7_w31_1_c1 <= tile_1_filtered_output_c1(14);
   bh7_w32_1_c1 <= tile_1_filtered_output_c1(15);
   bh7_w33_1_c1 <= tile_1_filtered_output_c1(16);
   bh7_w34_1_c1 <= tile_1_filtered_output_c1(17);
   bh7_w35_1_c1 <= tile_1_filtered_output_c1(18);
   bh7_w36_1_c1 <= tile_1_filtered_output_c1(19);
   bh7_w37_1_c1 <= tile_1_filtered_output_c1(20);
   bh7_w38_1_c1 <= tile_1_filtered_output_c1(21);
   bh7_w39_1_c1 <= tile_1_filtered_output_c1(22);
   bh7_w40_1_c1 <= tile_1_filtered_output_c1(23);
   bh7_w41_0_c1 <= tile_1_filtered_output_c1(24);
   bh7_w42_0_c1 <= tile_1_filtered_output_c1(25);
   bh7_w43_0_c1 <= tile_1_filtered_output_c1(26);
   bh7_w44_0_c1 <= tile_1_filtered_output_c1(27);
   bh7_w45_0_c1 <= tile_1_filtered_output_c1(28);
   bh7_w46_0_c1 <= tile_1_filtered_output_c1(29);
   bh7_w47_0_c1 <= tile_1_filtered_output_c1(30);
   bh7_w48_0_c1 <= tile_1_filtered_output_c1(31);
   bh7_w49_0_c1 <= tile_1_filtered_output_c1(32);
   bh7_w50_0_c1 <= tile_1_filtered_output_c1(33);
   bh7_w51_0_c1 <= tile_1_filtered_output_c1(34);
   bh7_w52_0_c1 <= tile_1_filtered_output_c1(35);
   bh7_w53_0_c1 <= tile_1_filtered_output_c1(36);
   bh7_w54_0_c1 <= tile_1_filtered_output_c1(37);
   bh7_w55_0_c1 <= tile_1_filtered_output_c1(38);
   bh7_w56_0_c1 <= tile_1_filtered_output_c1(39);
   bh7_w57_0_c1 <= tile_1_filtered_output_c1(40);
   tile_2_X_c0 <= X(50 downto 34);
   tile_2_Y_c0 <= Y(23 downto 0);
   tile_2_mult: DSPBlock_17x24_Freq500_uid13
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 X => tile_2_X_c0,
                 Y => tile_2_Y_c0,
                 R => tile_2_output_c1);

   tile_2_filtered_output_c1 <= unsigned(tile_2_output_c1(40 downto 0));
   bh7_w34_2_c1 <= tile_2_filtered_output_c1(0);
   bh7_w35_2_c1 <= tile_2_filtered_output_c1(1);
   bh7_w36_2_c1 <= tile_2_filtered_output_c1(2);
   bh7_w37_2_c1 <= tile_2_filtered_output_c1(3);
   bh7_w38_2_c1 <= tile_2_filtered_output_c1(4);
   bh7_w39_2_c1 <= tile_2_filtered_output_c1(5);
   bh7_w40_2_c1 <= tile_2_filtered_output_c1(6);
   bh7_w41_1_c1 <= tile_2_filtered_output_c1(7);
   bh7_w42_1_c1 <= tile_2_filtered_output_c1(8);
   bh7_w43_1_c1 <= tile_2_filtered_output_c1(9);
   bh7_w44_1_c1 <= tile_2_filtered_output_c1(10);
   bh7_w45_1_c1 <= tile_2_filtered_output_c1(11);
   bh7_w46_1_c1 <= tile_2_filtered_output_c1(12);
   bh7_w47_1_c1 <= tile_2_filtered_output_c1(13);
   bh7_w48_1_c1 <= tile_2_filtered_output_c1(14);
   bh7_w49_1_c1 <= tile_2_filtered_output_c1(15);
   bh7_w50_1_c1 <= tile_2_filtered_output_c1(16);
   bh7_w51_1_c1 <= tile_2_filtered_output_c1(17);
   bh7_w52_1_c1 <= tile_2_filtered_output_c1(18);
   bh7_w53_1_c1 <= tile_2_filtered_output_c1(19);
   bh7_w54_1_c1 <= tile_2_filtered_output_c1(20);
   bh7_w55_1_c1 <= tile_2_filtered_output_c1(21);
   bh7_w56_1_c1 <= tile_2_filtered_output_c1(22);
   bh7_w57_1_c1 <= tile_2_filtered_output_c1(23);
   bh7_w58_0_c1 <= tile_2_filtered_output_c1(24);
   bh7_w59_0_c1 <= tile_2_filtered_output_c1(25);
   bh7_w60_0_c1 <= tile_2_filtered_output_c1(26);
   bh7_w61_0_c1 <= tile_2_filtered_output_c1(27);
   bh7_w62_0_c1 <= tile_2_filtered_output_c1(28);
   bh7_w63_0_c1 <= tile_2_filtered_output_c1(29);
   bh7_w64_0_c1 <= tile_2_filtered_output_c1(30);
   bh7_w65_0_c1 <= tile_2_filtered_output_c1(31);
   bh7_w66_0_c1 <= tile_2_filtered_output_c1(32);
   bh7_w67_0_c1 <= tile_2_filtered_output_c1(33);
   bh7_w68_0_c1 <= tile_2_filtered_output_c1(34);
   bh7_w69_0_c1 <= tile_2_filtered_output_c1(35);
   bh7_w70_0_c1 <= tile_2_filtered_output_c1(36);
   bh7_w71_0_c1 <= tile_2_filtered_output_c1(37);
   bh7_w72_0_c1 <= tile_2_filtered_output_c1(38);
   bh7_w73_0_c1 <= tile_2_filtered_output_c1(39);
   bh7_w74_0_c1 <= tile_2_filtered_output_c1(40);
   tile_3_X_c0 <= X(52 downto 51);
   tile_3_Y_c0 <= Y(23 downto 21);
   tile_3_mult: IntMultiplierLUT_2x3_Freq500_uid15
      port map ( clk  => clk,
                 X => tile_3_X_c0,
                 Y => tile_3_Y_c0,
                 R => tile_3_output_c0);

   tile_3_filtered_output_c0 <= unsigned(tile_3_output_c0(4 downto 0));
   bh7_w72_1_c0 <= tile_3_filtered_output_c0(0);
   bh7_w73_1_c0 <= tile_3_filtered_output_c0(1);
   bh7_w74_1_c0 <= tile_3_filtered_output_c0(2);
   bh7_w75_0_c0 <= tile_3_filtered_output_c0(3);
   bh7_w76_0_c0 <= tile_3_filtered_output_c0(4);
   tile_4_X_c0 <= X(52 downto 51);
   tile_4_Y_c0 <= Y(20 downto 18);
   tile_4_mult: IntMultiplierLUT_2x3_Freq500_uid20
      port map ( clk  => clk,
                 X => tile_4_X_c0,
                 Y => tile_4_Y_c0,
                 R => tile_4_output_c0);

   tile_4_filtered_output_c0 <= unsigned(tile_4_output_c0(4 downto 0));
   bh7_w69_1_c0 <= tile_4_filtered_output_c0(0);
   bh7_w70_1_c0 <= tile_4_filtered_output_c0(1);
   bh7_w71_1_c0 <= tile_4_filtered_output_c0(2);
   bh7_w72_2_c0 <= tile_4_filtered_output_c0(3);
   bh7_w73_2_c0 <= tile_4_filtered_output_c0(4);
   tile_5_X_c0 <= X(52 downto 51);
   tile_5_Y_c0 <= Y(17 downto 15);
   tile_5_mult: IntMultiplierLUT_2x3_Freq500_uid25
      port map ( clk  => clk,
                 X => tile_5_X_c0,
                 Y => tile_5_Y_c0,
                 R => tile_5_output_c0);

   tile_5_filtered_output_c0 <= unsigned(tile_5_output_c0(4 downto 0));
   bh7_w66_1_c0 <= tile_5_filtered_output_c0(0);
   bh7_w67_1_c0 <= tile_5_filtered_output_c0(1);
   bh7_w68_1_c0 <= tile_5_filtered_output_c0(2);
   bh7_w69_2_c0 <= tile_5_filtered_output_c0(3);
   bh7_w70_2_c0 <= tile_5_filtered_output_c0(4);
   tile_6_X_c0 <= X(52 downto 51);
   tile_6_Y_c0 <= Y(14 downto 12);
   tile_6_mult: IntMultiplierLUT_2x3_Freq500_uid30
      port map ( clk  => clk,
                 X => tile_6_X_c0,
                 Y => tile_6_Y_c0,
                 R => tile_6_output_c0);

   tile_6_filtered_output_c0 <= unsigned(tile_6_output_c0(4 downto 0));
   bh7_w63_1_c0 <= tile_6_filtered_output_c0(0);
   bh7_w64_1_c0 <= tile_6_filtered_output_c0(1);
   bh7_w65_1_c0 <= tile_6_filtered_output_c0(2);
   bh7_w66_2_c0 <= tile_6_filtered_output_c0(3);
   bh7_w67_2_c0 <= tile_6_filtered_output_c0(4);
   tile_7_X_c0 <= X(52 downto 51);
   tile_7_Y_c0 <= Y(11 downto 9);
   tile_7_mult: IntMultiplierLUT_2x3_Freq500_uid35
      port map ( clk  => clk,
                 X => tile_7_X_c0,
                 Y => tile_7_Y_c0,
                 R => tile_7_output_c0);

   tile_7_filtered_output_c0 <= unsigned(tile_7_output_c0(4 downto 0));
   bh7_w60_1_c0 <= tile_7_filtered_output_c0(0);
   bh7_w61_1_c0 <= tile_7_filtered_output_c0(1);
   bh7_w62_1_c0 <= tile_7_filtered_output_c0(2);
   bh7_w63_2_c0 <= tile_7_filtered_output_c0(3);
   bh7_w64_2_c0 <= tile_7_filtered_output_c0(4);
   tile_8_X_c0 <= X(52 downto 51);
   tile_8_Y_c0 <= Y(8 downto 6);
   tile_8_mult: IntMultiplierLUT_2x3_Freq500_uid40
      port map ( clk  => clk,
                 X => tile_8_X_c0,
                 Y => tile_8_Y_c0,
                 R => tile_8_output_c0);

   tile_8_filtered_output_c0 <= unsigned(tile_8_output_c0(4 downto 0));
   bh7_w57_2_c0 <= tile_8_filtered_output_c0(0);
   bh7_w58_1_c0 <= tile_8_filtered_output_c0(1);
   bh7_w59_1_c0 <= tile_8_filtered_output_c0(2);
   bh7_w60_2_c0 <= tile_8_filtered_output_c0(3);
   bh7_w61_2_c0 <= tile_8_filtered_output_c0(4);
   tile_9_X_c0 <= X(52 downto 51);
   tile_9_Y_c0 <= Y(5 downto 3);
   tile_9_mult: IntMultiplierLUT_2x3_Freq500_uid45
      port map ( clk  => clk,
                 X => tile_9_X_c0,
                 Y => tile_9_Y_c0,
                 R => tile_9_output_c0);

   tile_9_filtered_output_c0 <= unsigned(tile_9_output_c0(4 downto 0));
   bh7_w54_2_c0 <= tile_9_filtered_output_c0(0);
   bh7_w55_2_c0 <= tile_9_filtered_output_c0(1);
   bh7_w56_2_c0 <= tile_9_filtered_output_c0(2);
   bh7_w57_3_c0 <= tile_9_filtered_output_c0(3);
   bh7_w58_2_c0 <= tile_9_filtered_output_c0(4);
   tile_10_X_c0 <= X(52 downto 51);
   tile_10_Y_c0 <= Y(2 downto 0);
   tile_10_mult: IntMultiplierLUT_2x3_Freq500_uid50
      port map ( clk  => clk,
                 X => tile_10_X_c0,
                 Y => tile_10_Y_c0,
                 R => tile_10_output_c0);

   tile_10_filtered_output_c0 <= unsigned(tile_10_output_c0(4 downto 0));
   bh7_w51_2_c0 <= tile_10_filtered_output_c0(0);
   bh7_w52_2_c0 <= tile_10_filtered_output_c0(1);
   bh7_w53_2_c0 <= tile_10_filtered_output_c0(2);
   bh7_w54_3_c0 <= tile_10_filtered_output_c0(3);
   bh7_w55_3_c0 <= tile_10_filtered_output_c0(4);
   tile_11_X_c0 <= X(16 downto 0);
   tile_11_Y_c0 <= Y(47 downto 24);
   tile_11_mult: DSPBlock_17x24_Freq500_uid55
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 X => tile_11_X_c0,
                 Y => tile_11_Y_c0,
                 R => tile_11_output_c1);

   tile_11_filtered_output_c1 <= unsigned(tile_11_output_c1(40 downto 0));
   bh7_w24_2_c1 <= tile_11_filtered_output_c1(0);
   bh7_w25_2_c1 <= tile_11_filtered_output_c1(1);
   bh7_w26_2_c1 <= tile_11_filtered_output_c1(2);
   bh7_w27_2_c1 <= tile_11_filtered_output_c1(3);
   bh7_w28_2_c1 <= tile_11_filtered_output_c1(4);
   bh7_w29_2_c1 <= tile_11_filtered_output_c1(5);
   bh7_w30_2_c1 <= tile_11_filtered_output_c1(6);
   bh7_w31_2_c1 <= tile_11_filtered_output_c1(7);
   bh7_w32_2_c1 <= tile_11_filtered_output_c1(8);
   bh7_w33_2_c1 <= tile_11_filtered_output_c1(9);
   bh7_w34_3_c1 <= tile_11_filtered_output_c1(10);
   bh7_w35_3_c1 <= tile_11_filtered_output_c1(11);
   bh7_w36_3_c1 <= tile_11_filtered_output_c1(12);
   bh7_w37_3_c1 <= tile_11_filtered_output_c1(13);
   bh7_w38_3_c1 <= tile_11_filtered_output_c1(14);
   bh7_w39_3_c1 <= tile_11_filtered_output_c1(15);
   bh7_w40_3_c1 <= tile_11_filtered_output_c1(16);
   bh7_w41_2_c1 <= tile_11_filtered_output_c1(17);
   bh7_w42_2_c1 <= tile_11_filtered_output_c1(18);
   bh7_w43_2_c1 <= tile_11_filtered_output_c1(19);
   bh7_w44_2_c1 <= tile_11_filtered_output_c1(20);
   bh7_w45_2_c1 <= tile_11_filtered_output_c1(21);
   bh7_w46_2_c1 <= tile_11_filtered_output_c1(22);
   bh7_w47_2_c1 <= tile_11_filtered_output_c1(23);
   bh7_w48_2_c1 <= tile_11_filtered_output_c1(24);
   bh7_w49_2_c1 <= tile_11_filtered_output_c1(25);
   bh7_w50_2_c1 <= tile_11_filtered_output_c1(26);
   bh7_w51_3_c1 <= tile_11_filtered_output_c1(27);
   bh7_w52_3_c1 <= tile_11_filtered_output_c1(28);
   bh7_w53_3_c1 <= tile_11_filtered_output_c1(29);
   bh7_w54_4_c1 <= tile_11_filtered_output_c1(30);
   bh7_w55_4_c1 <= tile_11_filtered_output_c1(31);
   bh7_w56_3_c1 <= tile_11_filtered_output_c1(32);
   bh7_w57_4_c1 <= tile_11_filtered_output_c1(33);
   bh7_w58_3_c1 <= tile_11_filtered_output_c1(34);
   bh7_w59_2_c1 <= tile_11_filtered_output_c1(35);
   bh7_w60_3_c1 <= tile_11_filtered_output_c1(36);
   bh7_w61_3_c1 <= tile_11_filtered_output_c1(37);
   bh7_w62_2_c1 <= tile_11_filtered_output_c1(38);
   bh7_w63_3_c1 <= tile_11_filtered_output_c1(39);
   bh7_w64_3_c1 <= tile_11_filtered_output_c1(40);
   tile_12_X_c0 <= X(33 downto 17);
   tile_12_Y_c0 <= Y(47 downto 24);
   tile_12_mult: DSPBlock_17x24_Freq500_uid57
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 X => tile_12_X_c0,
                 Y => tile_12_Y_c0,
                 R => tile_12_output_c1);

   tile_12_filtered_output_c1 <= unsigned(tile_12_output_c1(40 downto 0));
   bh7_w41_3_c1 <= tile_12_filtered_output_c1(0);
   bh7_w42_3_c1 <= tile_12_filtered_output_c1(1);
   bh7_w43_3_c1 <= tile_12_filtered_output_c1(2);
   bh7_w44_3_c1 <= tile_12_filtered_output_c1(3);
   bh7_w45_3_c1 <= tile_12_filtered_output_c1(4);
   bh7_w46_3_c1 <= tile_12_filtered_output_c1(5);
   bh7_w47_3_c1 <= tile_12_filtered_output_c1(6);
   bh7_w48_3_c1 <= tile_12_filtered_output_c1(7);
   bh7_w49_3_c1 <= tile_12_filtered_output_c1(8);
   bh7_w50_3_c1 <= tile_12_filtered_output_c1(9);
   bh7_w51_4_c1 <= tile_12_filtered_output_c1(10);
   bh7_w52_4_c1 <= tile_12_filtered_output_c1(11);
   bh7_w53_4_c1 <= tile_12_filtered_output_c1(12);
   bh7_w54_5_c1 <= tile_12_filtered_output_c1(13);
   bh7_w55_5_c1 <= tile_12_filtered_output_c1(14);
   bh7_w56_4_c1 <= tile_12_filtered_output_c1(15);
   bh7_w57_5_c1 <= tile_12_filtered_output_c1(16);
   bh7_w58_4_c1 <= tile_12_filtered_output_c1(17);
   bh7_w59_3_c1 <= tile_12_filtered_output_c1(18);
   bh7_w60_4_c1 <= tile_12_filtered_output_c1(19);
   bh7_w61_4_c1 <= tile_12_filtered_output_c1(20);
   bh7_w62_3_c1 <= tile_12_filtered_output_c1(21);
   bh7_w63_4_c1 <= tile_12_filtered_output_c1(22);
   bh7_w64_4_c1 <= tile_12_filtered_output_c1(23);
   bh7_w65_2_c1 <= tile_12_filtered_output_c1(24);
   bh7_w66_3_c1 <= tile_12_filtered_output_c1(25);
   bh7_w67_3_c1 <= tile_12_filtered_output_c1(26);
   bh7_w68_2_c1 <= tile_12_filtered_output_c1(27);
   bh7_w69_3_c1 <= tile_12_filtered_output_c1(28);
   bh7_w70_3_c1 <= tile_12_filtered_output_c1(29);
   bh7_w71_2_c1 <= tile_12_filtered_output_c1(30);
   bh7_w72_3_c1 <= tile_12_filtered_output_c1(31);
   bh7_w73_3_c1 <= tile_12_filtered_output_c1(32);
   bh7_w74_2_c1 <= tile_12_filtered_output_c1(33);
   bh7_w75_1_c1 <= tile_12_filtered_output_c1(34);
   bh7_w76_1_c1 <= tile_12_filtered_output_c1(35);
   bh7_w77_0_c1 <= tile_12_filtered_output_c1(36);
   bh7_w78_0_c1 <= tile_12_filtered_output_c1(37);
   bh7_w79_0_c1 <= tile_12_filtered_output_c1(38);
   bh7_w80_0_c1 <= tile_12_filtered_output_c1(39);
   bh7_w81_0_c1 <= tile_12_filtered_output_c1(40);
   tile_13_X_c0 <= X(50 downto 34);
   tile_13_Y_c0 <= Y(47 downto 24);
   tile_13_mult: DSPBlock_17x24_Freq500_uid59
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 X => tile_13_X_c0,
                 Y => tile_13_Y_c0,
                 R => tile_13_output_c1);

   tile_13_filtered_output_c1 <= unsigned(tile_13_output_c1(40 downto 0));
   bh7_w58_5_c1 <= tile_13_filtered_output_c1(0);
   bh7_w59_4_c1 <= tile_13_filtered_output_c1(1);
   bh7_w60_5_c1 <= tile_13_filtered_output_c1(2);
   bh7_w61_5_c1 <= tile_13_filtered_output_c1(3);
   bh7_w62_4_c1 <= tile_13_filtered_output_c1(4);
   bh7_w63_5_c1 <= tile_13_filtered_output_c1(5);
   bh7_w64_5_c1 <= tile_13_filtered_output_c1(6);
   bh7_w65_3_c1 <= tile_13_filtered_output_c1(7);
   bh7_w66_4_c1 <= tile_13_filtered_output_c1(8);
   bh7_w67_4_c1 <= tile_13_filtered_output_c1(9);
   bh7_w68_3_c1 <= tile_13_filtered_output_c1(10);
   bh7_w69_4_c1 <= tile_13_filtered_output_c1(11);
   bh7_w70_4_c1 <= tile_13_filtered_output_c1(12);
   bh7_w71_3_c1 <= tile_13_filtered_output_c1(13);
   bh7_w72_4_c1 <= tile_13_filtered_output_c1(14);
   bh7_w73_4_c1 <= tile_13_filtered_output_c1(15);
   bh7_w74_3_c1 <= tile_13_filtered_output_c1(16);
   bh7_w75_2_c1 <= tile_13_filtered_output_c1(17);
   bh7_w76_2_c1 <= tile_13_filtered_output_c1(18);
   bh7_w77_1_c1 <= tile_13_filtered_output_c1(19);
   bh7_w78_1_c1 <= tile_13_filtered_output_c1(20);
   bh7_w79_1_c1 <= tile_13_filtered_output_c1(21);
   bh7_w80_1_c1 <= tile_13_filtered_output_c1(22);
   bh7_w81_1_c1 <= tile_13_filtered_output_c1(23);
   bh7_w82_0_c1 <= tile_13_filtered_output_c1(24);
   bh7_w83_0_c1 <= tile_13_filtered_output_c1(25);
   bh7_w84_0_c1 <= tile_13_filtered_output_c1(26);
   bh7_w85_0_c1 <= tile_13_filtered_output_c1(27);
   bh7_w86_0_c1 <= tile_13_filtered_output_c1(28);
   bh7_w87_0_c1 <= tile_13_filtered_output_c1(29);
   bh7_w88_0_c1 <= tile_13_filtered_output_c1(30);
   bh7_w89_0_c1 <= tile_13_filtered_output_c1(31);
   bh7_w90_0_c1 <= tile_13_filtered_output_c1(32);
   bh7_w91_0_c1 <= tile_13_filtered_output_c1(33);
   bh7_w92_0_c1 <= tile_13_filtered_output_c1(34);
   bh7_w93_0_c1 <= tile_13_filtered_output_c1(35);
   bh7_w94_0_c1 <= tile_13_filtered_output_c1(36);
   bh7_w95_0_c1 <= tile_13_filtered_output_c1(37);
   bh7_w96_0_c1 <= tile_13_filtered_output_c1(38);
   bh7_w97_0_c1 <= tile_13_filtered_output_c1(39);
   bh7_w98_0_c1 <= tile_13_filtered_output_c1(40);
   tile_14_X_c0 <= X(52 downto 51);
   tile_14_Y_c0 <= Y(47 downto 45);
   tile_14_mult: IntMultiplierLUT_2x3_Freq500_uid61
      port map ( clk  => clk,
                 X => tile_14_X_c0,
                 Y => tile_14_Y_c0,
                 R => tile_14_output_c0);

   tile_14_filtered_output_c0 <= unsigned(tile_14_output_c0(4 downto 0));
   bh7_w96_1_c0 <= tile_14_filtered_output_c0(0);
   bh7_w97_1_c0 <= tile_14_filtered_output_c0(1);
   bh7_w98_1_c0 <= tile_14_filtered_output_c0(2);
   bh7_w99_0_c0 <= tile_14_filtered_output_c0(3);
   bh7_w100_0_c0 <= tile_14_filtered_output_c0(4);
   tile_15_X_c0 <= X(52 downto 51);
   tile_15_Y_c0 <= Y(44 downto 42);
   tile_15_mult: IntMultiplierLUT_2x3_Freq500_uid66
      port map ( clk  => clk,
                 X => tile_15_X_c0,
                 Y => tile_15_Y_c0,
                 R => tile_15_output_c0);

   tile_15_filtered_output_c0 <= unsigned(tile_15_output_c0(4 downto 0));
   bh7_w93_1_c0 <= tile_15_filtered_output_c0(0);
   bh7_w94_1_c0 <= tile_15_filtered_output_c0(1);
   bh7_w95_1_c0 <= tile_15_filtered_output_c0(2);
   bh7_w96_2_c0 <= tile_15_filtered_output_c0(3);
   bh7_w97_2_c0 <= tile_15_filtered_output_c0(4);
   tile_16_X_c0 <= X(52 downto 51);
   tile_16_Y_c0 <= Y(41 downto 39);
   tile_16_mult: IntMultiplierLUT_2x3_Freq500_uid71
      port map ( clk  => clk,
                 X => tile_16_X_c0,
                 Y => tile_16_Y_c0,
                 R => tile_16_output_c0);

   tile_16_filtered_output_c0 <= unsigned(tile_16_output_c0(4 downto 0));
   bh7_w90_1_c0 <= tile_16_filtered_output_c0(0);
   bh7_w91_1_c0 <= tile_16_filtered_output_c0(1);
   bh7_w92_1_c0 <= tile_16_filtered_output_c0(2);
   bh7_w93_2_c0 <= tile_16_filtered_output_c0(3);
   bh7_w94_2_c0 <= tile_16_filtered_output_c0(4);
   tile_17_X_c0 <= X(52 downto 51);
   tile_17_Y_c0 <= Y(38 downto 36);
   tile_17_mult: IntMultiplierLUT_2x3_Freq500_uid76
      port map ( clk  => clk,
                 X => tile_17_X_c0,
                 Y => tile_17_Y_c0,
                 R => tile_17_output_c0);

   tile_17_filtered_output_c0 <= unsigned(tile_17_output_c0(4 downto 0));
   bh7_w87_1_c0 <= tile_17_filtered_output_c0(0);
   bh7_w88_1_c0 <= tile_17_filtered_output_c0(1);
   bh7_w89_1_c0 <= tile_17_filtered_output_c0(2);
   bh7_w90_2_c0 <= tile_17_filtered_output_c0(3);
   bh7_w91_2_c0 <= tile_17_filtered_output_c0(4);
   tile_18_X_c0 <= X(52 downto 51);
   tile_18_Y_c0 <= Y(35 downto 33);
   tile_18_mult: IntMultiplierLUT_2x3_Freq500_uid81
      port map ( clk  => clk,
                 X => tile_18_X_c0,
                 Y => tile_18_Y_c0,
                 R => tile_18_output_c0);

   tile_18_filtered_output_c0 <= unsigned(tile_18_output_c0(4 downto 0));
   bh7_w84_1_c0 <= tile_18_filtered_output_c0(0);
   bh7_w85_1_c0 <= tile_18_filtered_output_c0(1);
   bh7_w86_1_c0 <= tile_18_filtered_output_c0(2);
   bh7_w87_2_c0 <= tile_18_filtered_output_c0(3);
   bh7_w88_2_c0 <= tile_18_filtered_output_c0(4);
   tile_19_X_c0 <= X(52 downto 51);
   tile_19_Y_c0 <= Y(32 downto 30);
   tile_19_mult: IntMultiplierLUT_2x3_Freq500_uid86
      port map ( clk  => clk,
                 X => tile_19_X_c0,
                 Y => tile_19_Y_c0,
                 R => tile_19_output_c0);

   tile_19_filtered_output_c0 <= unsigned(tile_19_output_c0(4 downto 0));
   bh7_w81_2_c0 <= tile_19_filtered_output_c0(0);
   bh7_w82_1_c0 <= tile_19_filtered_output_c0(1);
   bh7_w83_1_c0 <= tile_19_filtered_output_c0(2);
   bh7_w84_2_c0 <= tile_19_filtered_output_c0(3);
   bh7_w85_2_c0 <= tile_19_filtered_output_c0(4);
   tile_20_X_c0 <= X(52 downto 51);
   tile_20_Y_c0 <= Y(29 downto 27);
   tile_20_mult: IntMultiplierLUT_2x3_Freq500_uid91
      port map ( clk  => clk,
                 X => tile_20_X_c0,
                 Y => tile_20_Y_c0,
                 R => tile_20_output_c0);

   tile_20_filtered_output_c0 <= unsigned(tile_20_output_c0(4 downto 0));
   bh7_w78_2_c0 <= tile_20_filtered_output_c0(0);
   bh7_w79_2_c0 <= tile_20_filtered_output_c0(1);
   bh7_w80_2_c0 <= tile_20_filtered_output_c0(2);
   bh7_w81_3_c0 <= tile_20_filtered_output_c0(3);
   bh7_w82_2_c0 <= tile_20_filtered_output_c0(4);
   tile_21_X_c0 <= X(52 downto 51);
   tile_21_Y_c0 <= Y(26 downto 24);
   tile_21_mult: IntMultiplierLUT_2x3_Freq500_uid96
      port map ( clk  => clk,
                 X => tile_21_X_c0,
                 Y => tile_21_Y_c0,
                 R => tile_21_output_c0);

   tile_21_filtered_output_c0 <= unsigned(tile_21_output_c0(4 downto 0));
   bh7_w75_3_c0 <= tile_21_filtered_output_c0(0);
   bh7_w76_3_c0 <= tile_21_filtered_output_c0(1);
   bh7_w77_2_c0 <= tile_21_filtered_output_c0(2);
   bh7_w78_3_c0 <= tile_21_filtered_output_c0(3);
   bh7_w79_3_c0 <= tile_21_filtered_output_c0(4);
   tile_22_X_c0 <= X(16 downto 16);
   tile_22_Y_c0 <= Y(52 downto 52);
   tile_22_mult: IntMultiplierLUT_1x1_Freq500_uid101
      port map ( clk  => clk,
                 X => tile_22_X_c0,
                 Y => tile_22_Y_c0,
                 R => tile_22_output_c0);

   tile_22_filtered_output_c0 <= unsigned(tile_22_output_c0(0 downto 0));
   bh7_w68_4_c0 <= tile_22_filtered_output_c0(0);
   tile_23_X_c0 <= X(15 downto 12);
   tile_23_Y_c0 <= Y(52 downto 52);
   tile_23_mult: IntMultiplierLUT_4x1_Freq500_uid103
      port map ( clk  => clk,
                 X => tile_23_X_c0,
                 Y => tile_23_Y_c0,
                 R => tile_23_output_c0);

   tile_23_filtered_output_c0 <= unsigned(tile_23_output_c0(3 downto 0));
   bh7_w64_6_c0 <= tile_23_filtered_output_c0(0);
   bh7_w65_4_c0 <= tile_23_filtered_output_c0(1);
   bh7_w66_5_c0 <= tile_23_filtered_output_c0(2);
   bh7_w67_5_c0 <= tile_23_filtered_output_c0(3);
   tile_24_X_c0 <= X(11 downto 8);
   tile_24_Y_c0 <= Y(52 downto 52);
   tile_24_mult: IntMultiplierLUT_4x1_Freq500_uid105
      port map ( clk  => clk,
                 X => tile_24_X_c0,
                 Y => tile_24_Y_c0,
                 R => tile_24_output_c0);

   tile_24_filtered_output_c0 <= unsigned(tile_24_output_c0(3 downto 0));
   bh7_w60_6_c0 <= tile_24_filtered_output_c0(0);
   bh7_w61_6_c0 <= tile_24_filtered_output_c0(1);
   bh7_w62_5_c0 <= tile_24_filtered_output_c0(2);
   bh7_w63_6_c0 <= tile_24_filtered_output_c0(3);
   tile_25_X_c0 <= X(7 downto 4);
   tile_25_Y_c0 <= Y(52 downto 52);
   tile_25_mult: IntMultiplierLUT_4x1_Freq500_uid107
      port map ( clk  => clk,
                 X => tile_25_X_c0,
                 Y => tile_25_Y_c0,
                 R => tile_25_output_c0);

   tile_25_filtered_output_c0 <= unsigned(tile_25_output_c0(3 downto 0));
   bh7_w56_5_c0 <= tile_25_filtered_output_c0(0);
   bh7_w57_6_c0 <= tile_25_filtered_output_c0(1);
   bh7_w58_6_c0 <= tile_25_filtered_output_c0(2);
   bh7_w59_5_c0 <= tile_25_filtered_output_c0(3);
   tile_26_X_c0 <= X(3 downto 0);
   tile_26_Y_c0 <= Y(52 downto 52);
   tile_26_mult: IntMultiplierLUT_4x1_Freq500_uid109
      port map ( clk  => clk,
                 X => tile_26_X_c0,
                 Y => tile_26_Y_c0,
                 R => tile_26_output_c0);

   tile_26_filtered_output_c0 <= unsigned(tile_26_output_c0(3 downto 0));
   bh7_w52_5_c0 <= tile_26_filtered_output_c0(0);
   bh7_w53_5_c0 <= tile_26_filtered_output_c0(1);
   bh7_w54_6_c0 <= tile_26_filtered_output_c0(2);
   bh7_w55_6_c0 <= tile_26_filtered_output_c0(3);
   tile_27_X_c0 <= X(16 downto 15);
   tile_27_Y_c0 <= Y(51 downto 50);
   tile_27_mult: IntMultiplierLUT_2x2_Freq500_uid111
      port map ( clk  => clk,
                 X => tile_27_X_c0,
                 Y => tile_27_Y_c0,
                 R => tile_27_output_c0);

   tile_27_filtered_output_c0 <= unsigned(tile_27_output_c0(3 downto 0));
   bh7_w65_5_c0 <= tile_27_filtered_output_c0(0);
   bh7_w66_6_c0 <= tile_27_filtered_output_c0(1);
   bh7_w67_6_c0 <= tile_27_filtered_output_c0(2);
   bh7_w68_5_c0 <= tile_27_filtered_output_c0(3);
   tile_28_X_c0 <= X(14 downto 12);
   tile_28_Y_c0 <= Y(51 downto 50);
   tile_28_mult: IntMultiplierLUT_3x2_Freq500_uid116
      port map ( clk  => clk,
                 X => tile_28_X_c0,
                 Y => tile_28_Y_c0,
                 R => tile_28_output_c0);

   tile_28_filtered_output_c0 <= unsigned(tile_28_output_c0(4 downto 0));
   bh7_w62_6_c0 <= tile_28_filtered_output_c0(0);
   bh7_w63_7_c0 <= tile_28_filtered_output_c0(1);
   bh7_w64_7_c0 <= tile_28_filtered_output_c0(2);
   bh7_w65_6_c0 <= tile_28_filtered_output_c0(3);
   bh7_w66_7_c0 <= tile_28_filtered_output_c0(4);
   tile_29_X_c0 <= X(11 downto 9);
   tile_29_Y_c0 <= Y(51 downto 50);
   tile_29_mult: IntMultiplierLUT_3x2_Freq500_uid121
      port map ( clk  => clk,
                 X => tile_29_X_c0,
                 Y => tile_29_Y_c0,
                 R => tile_29_output_c0);

   tile_29_filtered_output_c0 <= unsigned(tile_29_output_c0(4 downto 0));
   bh7_w59_6_c0 <= tile_29_filtered_output_c0(0);
   bh7_w60_7_c0 <= tile_29_filtered_output_c0(1);
   bh7_w61_7_c0 <= tile_29_filtered_output_c0(2);
   bh7_w62_7_c0 <= tile_29_filtered_output_c0(3);
   bh7_w63_8_c0 <= tile_29_filtered_output_c0(4);
   tile_30_X_c0 <= X(8 downto 6);
   tile_30_Y_c0 <= Y(51 downto 50);
   tile_30_mult: IntMultiplierLUT_3x2_Freq500_uid126
      port map ( clk  => clk,
                 X => tile_30_X_c0,
                 Y => tile_30_Y_c0,
                 R => tile_30_output_c0);

   tile_30_filtered_output_c0 <= unsigned(tile_30_output_c0(4 downto 0));
   bh7_w56_6_c0 <= tile_30_filtered_output_c0(0);
   bh7_w57_7_c0 <= tile_30_filtered_output_c0(1);
   bh7_w58_7_c0 <= tile_30_filtered_output_c0(2);
   bh7_w59_7_c0 <= tile_30_filtered_output_c0(3);
   bh7_w60_8_c0 <= tile_30_filtered_output_c0(4);
   tile_31_X_c0 <= X(5 downto 3);
   tile_31_Y_c0 <= Y(51 downto 50);
   tile_31_mult: IntMultiplierLUT_3x2_Freq500_uid131
      port map ( clk  => clk,
                 X => tile_31_X_c0,
                 Y => tile_31_Y_c0,
                 R => tile_31_output_c0);

   tile_31_filtered_output_c0 <= unsigned(tile_31_output_c0(4 downto 0));
   bh7_w53_6_c0 <= tile_31_filtered_output_c0(0);
   bh7_w54_7_c0 <= tile_31_filtered_output_c0(1);
   bh7_w55_7_c0 <= tile_31_filtered_output_c0(2);
   bh7_w56_7_c0 <= tile_31_filtered_output_c0(3);
   bh7_w57_8_c0 <= tile_31_filtered_output_c0(4);
   tile_32_X_c0 <= X(2 downto 0);
   tile_32_Y_c0 <= Y(51 downto 50);
   tile_32_mult: IntMultiplierLUT_3x2_Freq500_uid136
      port map ( clk  => clk,
                 X => tile_32_X_c0,
                 Y => tile_32_Y_c0,
                 R => tile_32_output_c0);

   tile_32_filtered_output_c0 <= unsigned(tile_32_output_c0(4 downto 0));
   bh7_w50_4_c0 <= tile_32_filtered_output_c0(0);
   bh7_w51_5_c0 <= tile_32_filtered_output_c0(1);
   bh7_w52_6_c0 <= tile_32_filtered_output_c0(2);
   bh7_w53_7_c0 <= tile_32_filtered_output_c0(3);
   bh7_w54_8_c0 <= tile_32_filtered_output_c0(4);
   tile_33_X_c0 <= X(16 downto 15);
   tile_33_Y_c0 <= Y(49 downto 48);
   tile_33_mult: IntMultiplierLUT_2x2_Freq500_uid141
      port map ( clk  => clk,
                 X => tile_33_X_c0,
                 Y => tile_33_Y_c0,
                 R => tile_33_output_c0);

   tile_33_filtered_output_c0 <= unsigned(tile_33_output_c0(3 downto 0));
   bh7_w63_9_c0 <= tile_33_filtered_output_c0(0);
   bh7_w64_8_c0 <= tile_33_filtered_output_c0(1);
   bh7_w65_7_c0 <= tile_33_filtered_output_c0(2);
   bh7_w66_8_c0 <= tile_33_filtered_output_c0(3);
   tile_34_X_c0 <= X(14 downto 12);
   tile_34_Y_c0 <= Y(49 downto 48);
   tile_34_mult: IntMultiplierLUT_3x2_Freq500_uid146
      port map ( clk  => clk,
                 X => tile_34_X_c0,
                 Y => tile_34_Y_c0,
                 R => tile_34_output_c0);

   tile_34_filtered_output_c0 <= unsigned(tile_34_output_c0(4 downto 0));
   bh7_w60_9_c0 <= tile_34_filtered_output_c0(0);
   bh7_w61_8_c0 <= tile_34_filtered_output_c0(1);
   bh7_w62_8_c0 <= tile_34_filtered_output_c0(2);
   bh7_w63_10_c0 <= tile_34_filtered_output_c0(3);
   bh7_w64_9_c0 <= tile_34_filtered_output_c0(4);
   tile_35_X_c0 <= X(11 downto 9);
   tile_35_Y_c0 <= Y(49 downto 48);
   tile_35_mult: IntMultiplierLUT_3x2_Freq500_uid151
      port map ( clk  => clk,
                 X => tile_35_X_c0,
                 Y => tile_35_Y_c0,
                 R => tile_35_output_c0);

   tile_35_filtered_output_c0 <= unsigned(tile_35_output_c0(4 downto 0));
   bh7_w57_9_c0 <= tile_35_filtered_output_c0(0);
   bh7_w58_8_c0 <= tile_35_filtered_output_c0(1);
   bh7_w59_8_c0 <= tile_35_filtered_output_c0(2);
   bh7_w60_10_c0 <= tile_35_filtered_output_c0(3);
   bh7_w61_9_c0 <= tile_35_filtered_output_c0(4);
   tile_36_X_c0 <= X(8 downto 6);
   tile_36_Y_c0 <= Y(49 downto 48);
   tile_36_mult: IntMultiplierLUT_3x2_Freq500_uid156
      port map ( clk  => clk,
                 X => tile_36_X_c0,
                 Y => tile_36_Y_c0,
                 R => tile_36_output_c0);

   tile_36_filtered_output_c0 <= unsigned(tile_36_output_c0(4 downto 0));
   bh7_w54_9_c0 <= tile_36_filtered_output_c0(0);
   bh7_w55_8_c0 <= tile_36_filtered_output_c0(1);
   bh7_w56_8_c0 <= tile_36_filtered_output_c0(2);
   bh7_w57_10_c0 <= tile_36_filtered_output_c0(3);
   bh7_w58_9_c0 <= tile_36_filtered_output_c0(4);
   tile_37_X_c0 <= X(5 downto 3);
   tile_37_Y_c0 <= Y(49 downto 48);
   tile_37_mult: IntMultiplierLUT_3x2_Freq500_uid161
      port map ( clk  => clk,
                 X => tile_37_X_c0,
                 Y => tile_37_Y_c0,
                 R => tile_37_output_c0);

   tile_37_filtered_output_c0 <= unsigned(tile_37_output_c0(4 downto 0));
   bh7_w51_6_c0 <= tile_37_filtered_output_c0(0);
   bh7_w52_7_c0 <= tile_37_filtered_output_c0(1);
   bh7_w53_8_c0 <= tile_37_filtered_output_c0(2);
   bh7_w54_10_c0 <= tile_37_filtered_output_c0(3);
   bh7_w55_9_c0 <= tile_37_filtered_output_c0(4);
   tile_38_X_c0 <= X(2 downto 0);
   tile_38_Y_c0 <= Y(49 downto 48);
   tile_38_mult: IntMultiplierLUT_3x2_Freq500_uid166
      port map ( clk  => clk,
                 X => tile_38_X_c0,
                 Y => tile_38_Y_c0,
                 R => tile_38_output_c0);

   tile_38_filtered_output_c0 <= unsigned(tile_38_output_c0(4 downto 0));
   bh7_w48_4_c0 <= tile_38_filtered_output_c0(0);
   bh7_w49_4_c0 <= tile_38_filtered_output_c0(1);
   bh7_w50_5_c0 <= tile_38_filtered_output_c0(2);
   bh7_w51_7_c0 <= tile_38_filtered_output_c0(3);
   bh7_w52_8_c0 <= tile_38_filtered_output_c0(4);
   tile_39_X_c0 <= X(33 downto 33);
   tile_39_Y_c0 <= Y(52 downto 52);
   tile_39_mult: IntMultiplierLUT_1x1_Freq500_uid171
      port map ( clk  => clk,
                 X => tile_39_X_c0,
                 Y => tile_39_Y_c0,
                 R => tile_39_output_c0);

   tile_39_filtered_output_c0 <= unsigned(tile_39_output_c0(0 downto 0));
   bh7_w85_3_c0 <= tile_39_filtered_output_c0(0);
   tile_40_X_c0 <= X(32 downto 29);
   tile_40_Y_c0 <= Y(52 downto 52);
   tile_40_mult: IntMultiplierLUT_4x1_Freq500_uid173
      port map ( clk  => clk,
                 X => tile_40_X_c0,
                 Y => tile_40_Y_c0,
                 R => tile_40_output_c0);

   tile_40_filtered_output_c0 <= unsigned(tile_40_output_c0(3 downto 0));
   bh7_w81_4_c0 <= tile_40_filtered_output_c0(0);
   bh7_w82_3_c0 <= tile_40_filtered_output_c0(1);
   bh7_w83_2_c0 <= tile_40_filtered_output_c0(2);
   bh7_w84_3_c0 <= tile_40_filtered_output_c0(3);
   tile_41_X_c0 <= X(28 downto 25);
   tile_41_Y_c0 <= Y(52 downto 52);
   tile_41_mult: IntMultiplierLUT_4x1_Freq500_uid175
      port map ( clk  => clk,
                 X => tile_41_X_c0,
                 Y => tile_41_Y_c0,
                 R => tile_41_output_c0);

   tile_41_filtered_output_c0 <= unsigned(tile_41_output_c0(3 downto 0));
   bh7_w77_3_c0 <= tile_41_filtered_output_c0(0);
   bh7_w78_4_c0 <= tile_41_filtered_output_c0(1);
   bh7_w79_4_c0 <= tile_41_filtered_output_c0(2);
   bh7_w80_3_c0 <= tile_41_filtered_output_c0(3);
   tile_42_X_c0 <= X(24 downto 21);
   tile_42_Y_c0 <= Y(52 downto 52);
   tile_42_mult: IntMultiplierLUT_4x1_Freq500_uid177
      port map ( clk  => clk,
                 X => tile_42_X_c0,
                 Y => tile_42_Y_c0,
                 R => tile_42_output_c0);

   tile_42_filtered_output_c0 <= unsigned(tile_42_output_c0(3 downto 0));
   bh7_w73_5_c0 <= tile_42_filtered_output_c0(0);
   bh7_w74_4_c0 <= tile_42_filtered_output_c0(1);
   bh7_w75_4_c0 <= tile_42_filtered_output_c0(2);
   bh7_w76_4_c0 <= tile_42_filtered_output_c0(3);
   tile_43_X_c0 <= X(20 downto 17);
   tile_43_Y_c0 <= Y(52 downto 52);
   tile_43_mult: IntMultiplierLUT_4x1_Freq500_uid179
      port map ( clk  => clk,
                 X => tile_43_X_c0,
                 Y => tile_43_Y_c0,
                 R => tile_43_output_c0);

   tile_43_filtered_output_c0 <= unsigned(tile_43_output_c0(3 downto 0));
   bh7_w69_5_c0 <= tile_43_filtered_output_c0(0);
   bh7_w70_5_c0 <= tile_43_filtered_output_c0(1);
   bh7_w71_4_c0 <= tile_43_filtered_output_c0(2);
   bh7_w72_5_c0 <= tile_43_filtered_output_c0(3);
   tile_44_X_c0 <= X(33 downto 32);
   tile_44_Y_c0 <= Y(51 downto 50);
   tile_44_mult: IntMultiplierLUT_2x2_Freq500_uid181
      port map ( clk  => clk,
                 X => tile_44_X_c0,
                 Y => tile_44_Y_c0,
                 R => tile_44_output_c0);

   tile_44_filtered_output_c0 <= unsigned(tile_44_output_c0(3 downto 0));
   bh7_w82_4_c0 <= tile_44_filtered_output_c0(0);
   bh7_w83_3_c0 <= tile_44_filtered_output_c0(1);
   bh7_w84_4_c0 <= tile_44_filtered_output_c0(2);
   bh7_w85_4_c0 <= tile_44_filtered_output_c0(3);
   tile_45_X_c0 <= X(31 downto 29);
   tile_45_Y_c0 <= Y(51 downto 50);
   tile_45_mult: IntMultiplierLUT_3x2_Freq500_uid186
      port map ( clk  => clk,
                 X => tile_45_X_c0,
                 Y => tile_45_Y_c0,
                 R => tile_45_output_c0);

   tile_45_filtered_output_c0 <= unsigned(tile_45_output_c0(4 downto 0));
   bh7_w79_5_c0 <= tile_45_filtered_output_c0(0);
   bh7_w80_4_c0 <= tile_45_filtered_output_c0(1);
   bh7_w81_5_c0 <= tile_45_filtered_output_c0(2);
   bh7_w82_5_c0 <= tile_45_filtered_output_c0(3);
   bh7_w83_4_c0 <= tile_45_filtered_output_c0(4);
   tile_46_X_c0 <= X(28 downto 26);
   tile_46_Y_c0 <= Y(51 downto 50);
   tile_46_mult: IntMultiplierLUT_3x2_Freq500_uid191
      port map ( clk  => clk,
                 X => tile_46_X_c0,
                 Y => tile_46_Y_c0,
                 R => tile_46_output_c0);

   tile_46_filtered_output_c0 <= unsigned(tile_46_output_c0(4 downto 0));
   bh7_w76_5_c0 <= tile_46_filtered_output_c0(0);
   bh7_w77_4_c0 <= tile_46_filtered_output_c0(1);
   bh7_w78_5_c0 <= tile_46_filtered_output_c0(2);
   bh7_w79_6_c0 <= tile_46_filtered_output_c0(3);
   bh7_w80_5_c0 <= tile_46_filtered_output_c0(4);
   tile_47_X_c0 <= X(25 downto 23);
   tile_47_Y_c0 <= Y(51 downto 50);
   tile_47_mult: IntMultiplierLUT_3x2_Freq500_uid196
      port map ( clk  => clk,
                 X => tile_47_X_c0,
                 Y => tile_47_Y_c0,
                 R => tile_47_output_c0);

   tile_47_filtered_output_c0 <= unsigned(tile_47_output_c0(4 downto 0));
   bh7_w73_6_c0 <= tile_47_filtered_output_c0(0);
   bh7_w74_5_c0 <= tile_47_filtered_output_c0(1);
   bh7_w75_5_c0 <= tile_47_filtered_output_c0(2);
   bh7_w76_6_c0 <= tile_47_filtered_output_c0(3);
   bh7_w77_5_c0 <= tile_47_filtered_output_c0(4);
   tile_48_X_c0 <= X(22 downto 20);
   tile_48_Y_c0 <= Y(51 downto 50);
   tile_48_mult: IntMultiplierLUT_3x2_Freq500_uid201
      port map ( clk  => clk,
                 X => tile_48_X_c0,
                 Y => tile_48_Y_c0,
                 R => tile_48_output_c0);

   tile_48_filtered_output_c0 <= unsigned(tile_48_output_c0(4 downto 0));
   bh7_w70_6_c0 <= tile_48_filtered_output_c0(0);
   bh7_w71_5_c0 <= tile_48_filtered_output_c0(1);
   bh7_w72_6_c0 <= tile_48_filtered_output_c0(2);
   bh7_w73_7_c0 <= tile_48_filtered_output_c0(3);
   bh7_w74_6_c0 <= tile_48_filtered_output_c0(4);
   tile_49_X_c0 <= X(19 downto 17);
   tile_49_Y_c0 <= Y(51 downto 50);
   tile_49_mult: IntMultiplierLUT_3x2_Freq500_uid206
      port map ( clk  => clk,
                 X => tile_49_X_c0,
                 Y => tile_49_Y_c0,
                 R => tile_49_output_c0);

   tile_49_filtered_output_c0 <= unsigned(tile_49_output_c0(4 downto 0));
   bh7_w67_7_c0 <= tile_49_filtered_output_c0(0);
   bh7_w68_6_c0 <= tile_49_filtered_output_c0(1);
   bh7_w69_6_c0 <= tile_49_filtered_output_c0(2);
   bh7_w70_7_c0 <= tile_49_filtered_output_c0(3);
   bh7_w71_6_c0 <= tile_49_filtered_output_c0(4);
   tile_50_X_c0 <= X(33 downto 32);
   tile_50_Y_c0 <= Y(49 downto 48);
   tile_50_mult: IntMultiplierLUT_2x2_Freq500_uid211
      port map ( clk  => clk,
                 X => tile_50_X_c0,
                 Y => tile_50_Y_c0,
                 R => tile_50_output_c0);

   tile_50_filtered_output_c0 <= unsigned(tile_50_output_c0(3 downto 0));
   bh7_w80_6_c0 <= tile_50_filtered_output_c0(0);
   bh7_w81_6_c0 <= tile_50_filtered_output_c0(1);
   bh7_w82_6_c0 <= tile_50_filtered_output_c0(2);
   bh7_w83_5_c0 <= tile_50_filtered_output_c0(3);
   tile_51_X_c0 <= X(31 downto 29);
   tile_51_Y_c0 <= Y(49 downto 48);
   tile_51_mult: IntMultiplierLUT_3x2_Freq500_uid216
      port map ( clk  => clk,
                 X => tile_51_X_c0,
                 Y => tile_51_Y_c0,
                 R => tile_51_output_c0);

   tile_51_filtered_output_c0 <= unsigned(tile_51_output_c0(4 downto 0));
   bh7_w77_6_c0 <= tile_51_filtered_output_c0(0);
   bh7_w78_6_c0 <= tile_51_filtered_output_c0(1);
   bh7_w79_7_c0 <= tile_51_filtered_output_c0(2);
   bh7_w80_7_c0 <= tile_51_filtered_output_c0(3);
   bh7_w81_7_c0 <= tile_51_filtered_output_c0(4);
   tile_52_X_c0 <= X(28 downto 26);
   tile_52_Y_c0 <= Y(49 downto 48);
   tile_52_mult: IntMultiplierLUT_3x2_Freq500_uid221
      port map ( clk  => clk,
                 X => tile_52_X_c0,
                 Y => tile_52_Y_c0,
                 R => tile_52_output_c0);

   tile_52_filtered_output_c0 <= unsigned(tile_52_output_c0(4 downto 0));
   bh7_w74_7_c0 <= tile_52_filtered_output_c0(0);
   bh7_w75_6_c0 <= tile_52_filtered_output_c0(1);
   bh7_w76_7_c0 <= tile_52_filtered_output_c0(2);
   bh7_w77_7_c0 <= tile_52_filtered_output_c0(3);
   bh7_w78_7_c0 <= tile_52_filtered_output_c0(4);
   tile_53_X_c0 <= X(25 downto 23);
   tile_53_Y_c0 <= Y(49 downto 48);
   tile_53_mult: IntMultiplierLUT_3x2_Freq500_uid226
      port map ( clk  => clk,
                 X => tile_53_X_c0,
                 Y => tile_53_Y_c0,
                 R => tile_53_output_c0);

   tile_53_filtered_output_c0 <= unsigned(tile_53_output_c0(4 downto 0));
   bh7_w71_7_c0 <= tile_53_filtered_output_c0(0);
   bh7_w72_7_c0 <= tile_53_filtered_output_c0(1);
   bh7_w73_8_c0 <= tile_53_filtered_output_c0(2);
   bh7_w74_8_c0 <= tile_53_filtered_output_c0(3);
   bh7_w75_7_c0 <= tile_53_filtered_output_c0(4);
   tile_54_X_c0 <= X(22 downto 20);
   tile_54_Y_c0 <= Y(49 downto 48);
   tile_54_mult: IntMultiplierLUT_3x2_Freq500_uid231
      port map ( clk  => clk,
                 X => tile_54_X_c0,
                 Y => tile_54_Y_c0,
                 R => tile_54_output_c0);

   tile_54_filtered_output_c0 <= unsigned(tile_54_output_c0(4 downto 0));
   bh7_w68_7_c0 <= tile_54_filtered_output_c0(0);
   bh7_w69_7_c0 <= tile_54_filtered_output_c0(1);
   bh7_w70_8_c0 <= tile_54_filtered_output_c0(2);
   bh7_w71_8_c0 <= tile_54_filtered_output_c0(3);
   bh7_w72_8_c0 <= tile_54_filtered_output_c0(4);
   tile_55_X_c0 <= X(19 downto 17);
   tile_55_Y_c0 <= Y(49 downto 48);
   tile_55_mult: IntMultiplierLUT_3x2_Freq500_uid236
      port map ( clk  => clk,
                 X => tile_55_X_c0,
                 Y => tile_55_Y_c0,
                 R => tile_55_output_c0);

   tile_55_filtered_output_c0 <= unsigned(tile_55_output_c0(4 downto 0));
   bh7_w65_8_c0 <= tile_55_filtered_output_c0(0);
   bh7_w66_9_c0 <= tile_55_filtered_output_c0(1);
   bh7_w67_8_c0 <= tile_55_filtered_output_c0(2);
   bh7_w68_8_c0 <= tile_55_filtered_output_c0(3);
   bh7_w69_8_c0 <= tile_55_filtered_output_c0(4);
   tile_56_X_c0 <= X(50 downto 50);
   tile_56_Y_c0 <= Y(52 downto 52);
   tile_56_mult: IntMultiplierLUT_1x1_Freq500_uid241
      port map ( clk  => clk,
                 X => tile_56_X_c0,
                 Y => tile_56_Y_c0,
                 R => tile_56_output_c0);

   tile_56_filtered_output_c0 <= unsigned(tile_56_output_c0(0 downto 0));
   bh7_w102_0_c0 <= tile_56_filtered_output_c0(0);
   tile_57_X_c0 <= X(49 downto 46);
   tile_57_Y_c0 <= Y(52 downto 52);
   tile_57_mult: IntMultiplierLUT_4x1_Freq500_uid243
      port map ( clk  => clk,
                 X => tile_57_X_c0,
                 Y => tile_57_Y_c0,
                 R => tile_57_output_c0);

   tile_57_filtered_output_c0 <= unsigned(tile_57_output_c0(3 downto 0));
   bh7_w98_2_c0 <= tile_57_filtered_output_c0(0);
   bh7_w99_1_c0 <= tile_57_filtered_output_c0(1);
   bh7_w100_1_c0 <= tile_57_filtered_output_c0(2);
   bh7_w101_0_c0 <= tile_57_filtered_output_c0(3);
   tile_58_X_c0 <= X(45 downto 42);
   tile_58_Y_c0 <= Y(52 downto 52);
   tile_58_mult: IntMultiplierLUT_4x1_Freq500_uid245
      port map ( clk  => clk,
                 X => tile_58_X_c0,
                 Y => tile_58_Y_c0,
                 R => tile_58_output_c0);

   tile_58_filtered_output_c0 <= unsigned(tile_58_output_c0(3 downto 0));
   bh7_w94_3_c0 <= tile_58_filtered_output_c0(0);
   bh7_w95_2_c0 <= tile_58_filtered_output_c0(1);
   bh7_w96_3_c0 <= tile_58_filtered_output_c0(2);
   bh7_w97_3_c0 <= tile_58_filtered_output_c0(3);
   tile_59_X_c0 <= X(41 downto 38);
   tile_59_Y_c0 <= Y(52 downto 52);
   tile_59_mult: IntMultiplierLUT_4x1_Freq500_uid247
      port map ( clk  => clk,
                 X => tile_59_X_c0,
                 Y => tile_59_Y_c0,
                 R => tile_59_output_c0);

   tile_59_filtered_output_c0 <= unsigned(tile_59_output_c0(3 downto 0));
   bh7_w90_3_c0 <= tile_59_filtered_output_c0(0);
   bh7_w91_3_c0 <= tile_59_filtered_output_c0(1);
   bh7_w92_2_c0 <= tile_59_filtered_output_c0(2);
   bh7_w93_3_c0 <= tile_59_filtered_output_c0(3);
   tile_60_X_c0 <= X(37 downto 34);
   tile_60_Y_c0 <= Y(52 downto 52);
   tile_60_mult: IntMultiplierLUT_4x1_Freq500_uid249
      port map ( clk  => clk,
                 X => tile_60_X_c0,
                 Y => tile_60_Y_c0,
                 R => tile_60_output_c0);

   tile_60_filtered_output_c0 <= unsigned(tile_60_output_c0(3 downto 0));
   bh7_w86_2_c0 <= tile_60_filtered_output_c0(0);
   bh7_w87_3_c0 <= tile_60_filtered_output_c0(1);
   bh7_w88_3_c0 <= tile_60_filtered_output_c0(2);
   bh7_w89_2_c0 <= tile_60_filtered_output_c0(3);
   tile_61_X_c0 <= X(50 downto 49);
   tile_61_Y_c0 <= Y(51 downto 50);
   tile_61_mult: IntMultiplierLUT_2x2_Freq500_uid251
      port map ( clk  => clk,
                 X => tile_61_X_c0,
                 Y => tile_61_Y_c0,
                 R => tile_61_output_c0);

   tile_61_filtered_output_c0 <= unsigned(tile_61_output_c0(3 downto 0));
   bh7_w99_2_c0 <= tile_61_filtered_output_c0(0);
   bh7_w100_2_c0 <= tile_61_filtered_output_c0(1);
   bh7_w101_1_c0 <= tile_61_filtered_output_c0(2);
   bh7_w102_1_c0 <= tile_61_filtered_output_c0(3);
   tile_62_X_c0 <= X(48 downto 46);
   tile_62_Y_c0 <= Y(51 downto 50);
   tile_62_mult: IntMultiplierLUT_3x2_Freq500_uid256
      port map ( clk  => clk,
                 X => tile_62_X_c0,
                 Y => tile_62_Y_c0,
                 R => tile_62_output_c0);

   tile_62_filtered_output_c0 <= unsigned(tile_62_output_c0(4 downto 0));
   bh7_w96_4_c0 <= tile_62_filtered_output_c0(0);
   bh7_w97_4_c0 <= tile_62_filtered_output_c0(1);
   bh7_w98_3_c0 <= tile_62_filtered_output_c0(2);
   bh7_w99_3_c0 <= tile_62_filtered_output_c0(3);
   bh7_w100_3_c0 <= tile_62_filtered_output_c0(4);
   tile_63_X_c0 <= X(45 downto 43);
   tile_63_Y_c0 <= Y(51 downto 50);
   tile_63_mult: IntMultiplierLUT_3x2_Freq500_uid261
      port map ( clk  => clk,
                 X => tile_63_X_c0,
                 Y => tile_63_Y_c0,
                 R => tile_63_output_c0);

   tile_63_filtered_output_c0 <= unsigned(tile_63_output_c0(4 downto 0));
   bh7_w93_4_c0 <= tile_63_filtered_output_c0(0);
   bh7_w94_4_c0 <= tile_63_filtered_output_c0(1);
   bh7_w95_3_c0 <= tile_63_filtered_output_c0(2);
   bh7_w96_5_c0 <= tile_63_filtered_output_c0(3);
   bh7_w97_5_c0 <= tile_63_filtered_output_c0(4);
   tile_64_X_c0 <= X(42 downto 40);
   tile_64_Y_c0 <= Y(51 downto 50);
   tile_64_mult: IntMultiplierLUT_3x2_Freq500_uid266
      port map ( clk  => clk,
                 X => tile_64_X_c0,
                 Y => tile_64_Y_c0,
                 R => tile_64_output_c0);

   tile_64_filtered_output_c0 <= unsigned(tile_64_output_c0(4 downto 0));
   bh7_w90_4_c0 <= tile_64_filtered_output_c0(0);
   bh7_w91_4_c0 <= tile_64_filtered_output_c0(1);
   bh7_w92_3_c0 <= tile_64_filtered_output_c0(2);
   bh7_w93_5_c0 <= tile_64_filtered_output_c0(3);
   bh7_w94_5_c0 <= tile_64_filtered_output_c0(4);
   tile_65_X_c0 <= X(39 downto 37);
   tile_65_Y_c0 <= Y(51 downto 50);
   tile_65_mult: IntMultiplierLUT_3x2_Freq500_uid271
      port map ( clk  => clk,
                 X => tile_65_X_c0,
                 Y => tile_65_Y_c0,
                 R => tile_65_output_c0);

   tile_65_filtered_output_c0 <= unsigned(tile_65_output_c0(4 downto 0));
   bh7_w87_4_c0 <= tile_65_filtered_output_c0(0);
   bh7_w88_4_c0 <= tile_65_filtered_output_c0(1);
   bh7_w89_3_c0 <= tile_65_filtered_output_c0(2);
   bh7_w90_5_c0 <= tile_65_filtered_output_c0(3);
   bh7_w91_5_c0 <= tile_65_filtered_output_c0(4);
   tile_66_X_c0 <= X(36 downto 34);
   tile_66_Y_c0 <= Y(51 downto 50);
   tile_66_mult: IntMultiplierLUT_3x2_Freq500_uid276
      port map ( clk  => clk,
                 X => tile_66_X_c0,
                 Y => tile_66_Y_c0,
                 R => tile_66_output_c0);

   tile_66_filtered_output_c0 <= unsigned(tile_66_output_c0(4 downto 0));
   bh7_w84_5_c0 <= tile_66_filtered_output_c0(0);
   bh7_w85_5_c0 <= tile_66_filtered_output_c0(1);
   bh7_w86_3_c0 <= tile_66_filtered_output_c0(2);
   bh7_w87_5_c0 <= tile_66_filtered_output_c0(3);
   bh7_w88_5_c0 <= tile_66_filtered_output_c0(4);
   tile_67_X_c0 <= X(50 downto 49);
   tile_67_Y_c0 <= Y(49 downto 48);
   tile_67_mult: IntMultiplierLUT_2x2_Freq500_uid281
      port map ( clk  => clk,
                 X => tile_67_X_c0,
                 Y => tile_67_Y_c0,
                 R => tile_67_output_c0);

   tile_67_filtered_output_c0 <= unsigned(tile_67_output_c0(3 downto 0));
   bh7_w97_6_c0 <= tile_67_filtered_output_c0(0);
   bh7_w98_4_c0 <= tile_67_filtered_output_c0(1);
   bh7_w99_4_c0 <= tile_67_filtered_output_c0(2);
   bh7_w100_4_c0 <= tile_67_filtered_output_c0(3);
   tile_68_X_c0 <= X(48 downto 46);
   tile_68_Y_c0 <= Y(49 downto 48);
   tile_68_mult: IntMultiplierLUT_3x2_Freq500_uid286
      port map ( clk  => clk,
                 X => tile_68_X_c0,
                 Y => tile_68_Y_c0,
                 R => tile_68_output_c0);

   tile_68_filtered_output_c0 <= unsigned(tile_68_output_c0(4 downto 0));
   bh7_w94_6_c0 <= tile_68_filtered_output_c0(0);
   bh7_w95_4_c0 <= tile_68_filtered_output_c0(1);
   bh7_w96_6_c0 <= tile_68_filtered_output_c0(2);
   bh7_w97_7_c0 <= tile_68_filtered_output_c0(3);
   bh7_w98_5_c0 <= tile_68_filtered_output_c0(4);
   tile_69_X_c0 <= X(45 downto 43);
   tile_69_Y_c0 <= Y(49 downto 48);
   tile_69_mult: IntMultiplierLUT_3x2_Freq500_uid291
      port map ( clk  => clk,
                 X => tile_69_X_c0,
                 Y => tile_69_Y_c0,
                 R => tile_69_output_c0);

   tile_69_filtered_output_c0 <= unsigned(tile_69_output_c0(4 downto 0));
   bh7_w91_6_c0 <= tile_69_filtered_output_c0(0);
   bh7_w92_4_c0 <= tile_69_filtered_output_c0(1);
   bh7_w93_6_c0 <= tile_69_filtered_output_c0(2);
   bh7_w94_7_c0 <= tile_69_filtered_output_c0(3);
   bh7_w95_5_c0 <= tile_69_filtered_output_c0(4);
   tile_70_X_c0 <= X(42 downto 40);
   tile_70_Y_c0 <= Y(49 downto 48);
   tile_70_mult: IntMultiplierLUT_3x2_Freq500_uid296
      port map ( clk  => clk,
                 X => tile_70_X_c0,
                 Y => tile_70_Y_c0,
                 R => tile_70_output_c0);

   tile_70_filtered_output_c0 <= unsigned(tile_70_output_c0(4 downto 0));
   bh7_w88_6_c0 <= tile_70_filtered_output_c0(0);
   bh7_w89_4_c0 <= tile_70_filtered_output_c0(1);
   bh7_w90_6_c0 <= tile_70_filtered_output_c0(2);
   bh7_w91_7_c0 <= tile_70_filtered_output_c0(3);
   bh7_w92_5_c0 <= tile_70_filtered_output_c0(4);
   tile_71_X_c0 <= X(39 downto 37);
   tile_71_Y_c0 <= Y(49 downto 48);
   tile_71_mult: IntMultiplierLUT_3x2_Freq500_uid301
      port map ( clk  => clk,
                 X => tile_71_X_c0,
                 Y => tile_71_Y_c0,
                 R => tile_71_output_c0);

   tile_71_filtered_output_c0 <= unsigned(tile_71_output_c0(4 downto 0));
   bh7_w85_6_c0 <= tile_71_filtered_output_c0(0);
   bh7_w86_4_c0 <= tile_71_filtered_output_c0(1);
   bh7_w87_6_c0 <= tile_71_filtered_output_c0(2);
   bh7_w88_7_c0 <= tile_71_filtered_output_c0(3);
   bh7_w89_5_c0 <= tile_71_filtered_output_c0(4);
   tile_72_X_c0 <= X(36 downto 34);
   tile_72_Y_c0 <= Y(49 downto 48);
   tile_72_mult: IntMultiplierLUT_3x2_Freq500_uid306
      port map ( clk  => clk,
                 X => tile_72_X_c0,
                 Y => tile_72_Y_c0,
                 R => tile_72_output_c0);

   tile_72_filtered_output_c0 <= unsigned(tile_72_output_c0(4 downto 0));
   bh7_w82_7_c0 <= tile_72_filtered_output_c0(0);
   bh7_w83_6_c0 <= tile_72_filtered_output_c0(1);
   bh7_w84_6_c0 <= tile_72_filtered_output_c0(2);
   bh7_w85_7_c0 <= tile_72_filtered_output_c0(3);
   bh7_w86_5_c0 <= tile_72_filtered_output_c0(4);
   tile_73_X_c0 <= X(52 downto 51);
   tile_73_Y_c0 <= Y(52 downto 51);
   tile_73_mult: IntMultiplierLUT_2x2_Freq500_uid311
      port map ( clk  => clk,
                 X => tile_73_X_c0,
                 Y => tile_73_Y_c0,
                 R => tile_73_output_c0);

   tile_73_filtered_output_c0 <= unsigned(tile_73_output_c0(3 downto 0));
   bh7_w102_2_c0 <= tile_73_filtered_output_c0(0);
   bh7_w103_0_c0 <= tile_73_filtered_output_c0(1);
   bh7_w104_0_c0 <= tile_73_filtered_output_c0(2);
   bh7_w105_0_c0 <= tile_73_filtered_output_c0(3);
   tile_74_X_c0 <= X(52 downto 51);
   tile_74_Y_c0 <= Y(50 downto 48);
   tile_74_mult: IntMultiplierLUT_2x3_Freq500_uid316
      port map ( clk  => clk,
                 X => tile_74_X_c0,
                 Y => tile_74_Y_c0,
                 R => tile_74_output_c0);

   tile_74_filtered_output_c0 <= unsigned(tile_74_output_c0(4 downto 0));
   bh7_w99_5_c0 <= tile_74_filtered_output_c0(0);
   bh7_w100_5_c0 <= tile_74_filtered_output_c0(1);
   bh7_w101_2_c0 <= tile_74_filtered_output_c0(2);
   bh7_w102_3_c0 <= tile_74_filtered_output_c0(3);
   bh7_w103_1_c0 <= tile_74_filtered_output_c0(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq500_uid322_bh7_uid323_In0_c0 <= "" & bh7_w49_4_c0 & "0" & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid323_In1_c0 <= "" & bh7_w50_4_c0 & bh7_w50_5_c0;
   bh7_w49_5_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid323_Out0_c0(0);
   bh7_w50_6_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid323_Out0_c0(1);
   bh7_w51_8_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid323_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid323: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid323_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid323_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid323_Out0_copy324_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid323_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid323_Out0_copy324_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid327_In0_c0 <= "" & bh7_w51_2_c0 & bh7_w51_5_c0 & bh7_w51_6_c0 & bh7_w51_7_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid327_In1_c0 <= "" & bh7_w52_2_c0;
   bh7_w51_9_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid327_Out0_c0(0);
   bh7_w52_9_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid327_Out0_c0(1);
   bh7_w53_9_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid327_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid327: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid327_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid327_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid327_Out0_copy328_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid327_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid327_Out0_copy328_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid329_In0_c0 <= "" & bh7_w52_5_c0 & bh7_w52_6_c0 & bh7_w52_7_c0 & bh7_w52_8_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid329_In1_c0 <= "" & bh7_w53_2_c0;
   bh7_w52_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid329_Out0_c0(0);
   bh7_w53_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid329_Out0_c0(1);
   bh7_w54_11_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid329_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid329: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid329_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid329_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid329_Out0_copy330_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid329_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid329_Out0_copy330_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid331_In0_c0 <= "" & bh7_w53_5_c0 & bh7_w53_6_c0 & bh7_w53_7_c0 & bh7_w53_8_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid331_In1_c0 <= "" & bh7_w54_2_c0;
   bh7_w53_11_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid331_Out0_c0(0);
   bh7_w54_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid331_Out0_c0(1);
   bh7_w55_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid331_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid331: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid331_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid331_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid331_Out0_copy332_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid331_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid331_Out0_copy332_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid335_In0_c0 <= "" & bh7_w54_3_c0 & bh7_w54_6_c0 & bh7_w54_7_c0 & bh7_w54_8_c0 & bh7_w54_9_c0 & bh7_w54_10_c0;
   bh7_w54_13_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid335_Out0_c0(0);
   bh7_w55_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid335_Out0_c0(1);
   bh7_w56_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid335_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid335: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid335_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid335_Out0_copy336_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid335_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid335_Out0_copy336_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid337_In0_c0 <= "" & bh7_w55_2_c0 & bh7_w55_3_c0 & bh7_w55_6_c0 & bh7_w55_7_c0 & bh7_w55_8_c0 & bh7_w55_9_c0;
   bh7_w55_12_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid337_Out0_c0(0);
   bh7_w56_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid337_Out0_c0(1);
   bh7_w57_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid337_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid337: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid337_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid337_Out0_copy338_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid337_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid337_Out0_copy338_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid339_In0_c0 <= "" & bh7_w56_2_c0 & bh7_w56_5_c0 & bh7_w56_6_c0 & bh7_w56_7_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid339_In1_c0 <= "" & bh7_w57_2_c0;
   bh7_w56_11_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid339_Out0_c0(0);
   bh7_w57_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid339_Out0_c0(1);
   bh7_w58_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid339_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid339: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid339_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid339_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid339_Out0_copy340_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid339_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid339_Out0_copy340_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid341_In0_c0 <= "" & bh7_w57_3_c0 & bh7_w57_6_c0 & bh7_w57_7_c0 & bh7_w57_8_c0 & bh7_w57_9_c0 & bh7_w57_10_c0;
   bh7_w57_13_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid341_Out0_c0(0);
   bh7_w58_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid341_Out0_c0(1);
   bh7_w59_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid341_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid341: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid341_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid341_Out0_copy342_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid341_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid341_Out0_copy342_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid343_In0_c0 <= "" & bh7_w58_1_c0 & bh7_w58_2_c0 & bh7_w58_6_c0 & bh7_w58_7_c0 & bh7_w58_8_c0 & bh7_w58_9_c0;
   bh7_w58_12_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid343_Out0_c0(0);
   bh7_w59_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid343_Out0_c0(1);
   bh7_w60_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid343_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid343: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid343_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid343_Out0_copy344_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid343_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid343_Out0_copy344_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid345_In0_c0 <= "" & bh7_w59_1_c0 & bh7_w59_5_c0 & bh7_w59_6_c0 & bh7_w59_7_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid345_In1_c0 <= "" & bh7_w60_1_c0;
   bh7_w59_11_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid345_Out0_c0(0);
   bh7_w60_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid345_Out0_c0(1);
   bh7_w61_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid345_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid345: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid345_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid345_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid345_Out0_copy346_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid345_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid345_Out0_copy346_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid347_In0_c0 <= "" & bh7_w60_2_c0 & bh7_w60_6_c0 & bh7_w60_7_c0 & bh7_w60_8_c0 & bh7_w60_9_c0 & bh7_w60_10_c0;
   bh7_w60_13_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid347_Out0_c0(0);
   bh7_w61_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid347_Out0_c0(1);
   bh7_w62_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid347_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid347: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid347_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid347_Out0_copy348_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid347_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid347_Out0_copy348_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid349_In0_c0 <= "" & bh7_w61_1_c0 & bh7_w61_2_c0 & bh7_w61_6_c0 & bh7_w61_7_c0 & bh7_w61_8_c0 & bh7_w61_9_c0;
   bh7_w61_12_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid349_Out0_c0(0);
   bh7_w62_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid349_Out0_c0(1);
   bh7_w63_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid349_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid349: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid349_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid349_Out0_copy350_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid349_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid349_Out0_copy350_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid351_In0_c0 <= "" & bh7_w62_1_c0 & bh7_w62_5_c0 & bh7_w62_6_c0 & bh7_w62_7_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid351_In1_c0 <= "" & bh7_w63_1_c0;
   bh7_w62_11_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid351_Out0_c0(0);
   bh7_w63_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid351_Out0_c0(1);
   bh7_w64_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid351_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid351: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid351_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid351_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid351_Out0_copy352_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid351_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid351_Out0_copy352_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid353_In0_c0 <= "" & bh7_w63_2_c0 & bh7_w63_6_c0 & bh7_w63_7_c0 & bh7_w63_8_c0 & bh7_w63_9_c0 & bh7_w63_10_c0;
   bh7_w63_13_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid353_Out0_c0(0);
   bh7_w64_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid353_Out0_c0(1);
   bh7_w65_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid353_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid353: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid353_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid353_Out0_copy354_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid353_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid353_Out0_copy354_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid355_In0_c0 <= "" & bh7_w64_1_c0 & bh7_w64_2_c0 & bh7_w64_6_c0 & bh7_w64_7_c0 & bh7_w64_8_c0 & bh7_w64_9_c0;
   bh7_w64_12_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid355_Out0_c0(0);
   bh7_w65_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid355_Out0_c0(1);
   bh7_w66_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid355_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid355: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid355_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid355_Out0_copy356_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid355_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid355_Out0_copy356_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid357_In0_c0 <= "" & bh7_w65_1_c0 & bh7_w65_4_c0 & bh7_w65_5_c0 & bh7_w65_6_c0 & bh7_w65_7_c0 & bh7_w65_8_c0;
   bh7_w65_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid357_Out0_c0(0);
   bh7_w66_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid357_Out0_c0(1);
   bh7_w67_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid357_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid357: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid357_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid357_Out0_copy358_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid357_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid357_Out0_copy358_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid359_In0_c0 <= "" & bh7_w66_1_c0 & bh7_w66_2_c0 & bh7_w66_5_c0 & bh7_w66_6_c0 & bh7_w66_7_c0 & bh7_w66_8_c0;
   bh7_w66_12_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid359_Out0_c0(0);
   bh7_w67_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid359_Out0_c0(1);
   bh7_w68_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid359_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid359: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid359_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid359_Out0_copy360_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid359_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid359_Out0_copy360_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid361_In0_c0 <= "" & bh7_w67_1_c0 & bh7_w67_2_c0 & bh7_w67_5_c0 & bh7_w67_6_c0 & bh7_w67_7_c0 & bh7_w67_8_c0;
   bh7_w67_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid361_Out0_c0(0);
   bh7_w68_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid361_Out0_c0(1);
   bh7_w69_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid361_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid361: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid361_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid361_Out0_copy362_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid361_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid361_Out0_copy362_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid363_In0_c0 <= "" & bh7_w68_1_c0 & bh7_w68_4_c0 & bh7_w68_5_c0 & bh7_w68_6_c0 & bh7_w68_7_c0 & bh7_w68_8_c0;
   bh7_w68_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid363_Out0_c0(0);
   bh7_w69_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid363_Out0_c0(1);
   bh7_w70_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid363_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid363: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid363_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid363_Out0_copy364_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid363_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid363_Out0_copy364_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid365_In0_c0 <= "" & bh7_w69_1_c0 & bh7_w69_2_c0 & bh7_w69_5_c0 & bh7_w69_6_c0 & bh7_w69_7_c0 & bh7_w69_8_c0;
   bh7_w69_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid365_Out0_c0(0);
   bh7_w70_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid365_Out0_c0(1);
   bh7_w71_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid365_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid365: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid365_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid365_Out0_copy366_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid365_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid365_Out0_copy366_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid367_In0_c0 <= "" & bh7_w70_1_c0 & bh7_w70_2_c0 & bh7_w70_5_c0 & bh7_w70_6_c0 & bh7_w70_7_c0 & bh7_w70_8_c0;
   bh7_w70_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid367_Out0_c0(0);
   bh7_w71_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid367_Out0_c0(1);
   bh7_w72_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid367_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid367: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid367_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid367_Out0_copy368_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid367_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid367_Out0_copy368_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid369_In0_c0 <= "" & bh7_w71_1_c0 & bh7_w71_4_c0 & bh7_w71_5_c0 & bh7_w71_6_c0 & bh7_w71_7_c0 & bh7_w71_8_c0;
   bh7_w71_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid369_Out0_c0(0);
   bh7_w72_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid369_Out0_c0(1);
   bh7_w73_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid369_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid369: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid369_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid369_Out0_copy370_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid369_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid369_Out0_copy370_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid371_In0_c0 <= "" & bh7_w72_1_c0 & bh7_w72_2_c0 & bh7_w72_5_c0 & bh7_w72_6_c0 & bh7_w72_7_c0 & bh7_w72_8_c0;
   bh7_w72_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid371_Out0_c0(0);
   bh7_w73_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid371_Out0_c0(1);
   bh7_w74_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid371_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid371: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid371_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid371_Out0_copy372_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid371_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid371_Out0_copy372_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid373_In0_c0 <= "" & bh7_w73_1_c0 & bh7_w73_2_c0 & bh7_w73_5_c0 & bh7_w73_6_c0 & bh7_w73_7_c0 & bh7_w73_8_c0;
   bh7_w73_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid373_Out0_c0(0);
   bh7_w74_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid373_Out0_c0(1);
   bh7_w75_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid373_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid373: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid373_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid373_Out0_copy374_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid373_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid373_Out0_copy374_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid375_In0_c0 <= "" & bh7_w74_1_c0 & bh7_w74_4_c0 & bh7_w74_5_c0 & bh7_w74_6_c0 & bh7_w74_7_c0 & bh7_w74_8_c0;
   bh7_w74_11_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid375_Out0_c0(0);
   bh7_w75_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid375_Out0_c0(1);
   bh7_w76_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid375_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid375: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid375_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid375_Out0_copy376_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid375_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid375_Out0_copy376_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid377_In0_c0 <= "" & bh7_w75_0_c0 & bh7_w75_3_c0 & bh7_w75_4_c0 & bh7_w75_5_c0 & bh7_w75_6_c0 & bh7_w75_7_c0;
   bh7_w75_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid377_Out0_c0(0);
   bh7_w76_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid377_Out0_c0(1);
   bh7_w77_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid377_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid377: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid377_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid377_Out0_copy378_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid377_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid377_Out0_copy378_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid379_In0_c0 <= "" & bh7_w76_0_c0 & bh7_w76_3_c0 & bh7_w76_4_c0 & bh7_w76_5_c0 & bh7_w76_6_c0 & bh7_w76_7_c0;
   bh7_w76_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid379_Out0_c0(0);
   bh7_w77_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid379_Out0_c0(1);
   bh7_w78_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid379_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid379: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid379_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid379_Out0_copy380_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid379_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid379_Out0_copy380_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid381_In0_c0 <= "" & bh7_w77_2_c0 & bh7_w77_3_c0 & bh7_w77_4_c0 & bh7_w77_5_c0 & bh7_w77_6_c0 & bh7_w77_7_c0;
   bh7_w77_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid381_Out0_c0(0);
   bh7_w78_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid381_Out0_c0(1);
   bh7_w79_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid381_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid381: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid381_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid381_Out0_copy382_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid381_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid381_Out0_copy382_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid383_In0_c0 <= "" & bh7_w78_2_c0 & bh7_w78_3_c0 & bh7_w78_4_c0 & bh7_w78_5_c0 & bh7_w78_6_c0 & bh7_w78_7_c0;
   bh7_w78_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid383_Out0_c0(0);
   bh7_w79_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid383_Out0_c0(1);
   bh7_w80_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid383_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid383: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid383_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid383_Out0_copy384_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid383_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid383_Out0_copy384_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid385_In0_c0 <= "" & bh7_w79_2_c0 & bh7_w79_3_c0 & bh7_w79_4_c0 & bh7_w79_5_c0 & bh7_w79_6_c0 & bh7_w79_7_c0;
   bh7_w79_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid385_Out0_c0(0);
   bh7_w80_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid385_Out0_c0(1);
   bh7_w81_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid385_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid385: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid385_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid385_Out0_copy386_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid385_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid385_Out0_copy386_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid387_In0_c0 <= "" & bh7_w80_2_c0 & bh7_w80_3_c0 & bh7_w80_4_c0 & bh7_w80_5_c0 & bh7_w80_6_c0 & bh7_w80_7_c0;
   bh7_w80_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid387_Out0_c0(0);
   bh7_w81_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid387_Out0_c0(1);
   bh7_w82_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid387_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid387: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid387_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid387_Out0_copy388_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid387_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid387_Out0_copy388_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid389_In0_c0 <= "" & bh7_w81_2_c0 & bh7_w81_3_c0 & bh7_w81_4_c0 & bh7_w81_5_c0 & bh7_w81_6_c0 & bh7_w81_7_c0;
   bh7_w81_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid389_Out0_c0(0);
   bh7_w82_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid389_Out0_c0(1);
   bh7_w83_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid389_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid389: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid389_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid389_Out0_copy390_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid389_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid389_Out0_copy390_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid391_In0_c0 <= "" & bh7_w82_1_c0 & bh7_w82_2_c0 & bh7_w82_3_c0 & bh7_w82_4_c0 & bh7_w82_5_c0 & bh7_w82_6_c0;
   bh7_w82_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid391_Out0_c0(0);
   bh7_w83_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid391_Out0_c0(1);
   bh7_w84_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid391_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid391: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid391_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid391_Out0_copy392_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid391_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid391_Out0_copy392_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid393_In0_c0 <= "" & bh7_w83_1_c0 & bh7_w83_2_c0 & bh7_w83_3_c0 & bh7_w83_4_c0 & bh7_w83_5_c0 & bh7_w83_6_c0;
   bh7_w83_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid393_Out0_c0(0);
   bh7_w84_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid393_Out0_c0(1);
   bh7_w85_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid393_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid393: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid393_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid393_Out0_copy394_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid393_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid393_Out0_copy394_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid395_In0_c0 <= "" & bh7_w84_1_c0 & bh7_w84_2_c0 & bh7_w84_3_c0 & bh7_w84_4_c0 & bh7_w84_5_c0 & bh7_w84_6_c0;
   bh7_w84_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid395_Out0_c0(0);
   bh7_w85_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid395_Out0_c0(1);
   bh7_w86_6_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid395_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid395: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid395_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid395_Out0_copy396_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid395_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid395_Out0_copy396_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid397_In0_c0 <= "" & bh7_w85_1_c0 & bh7_w85_2_c0 & bh7_w85_3_c0 & bh7_w85_4_c0 & bh7_w85_5_c0 & bh7_w85_6_c0;
   bh7_w85_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid397_Out0_c0(0);
   bh7_w86_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid397_Out0_c0(1);
   bh7_w87_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid397_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid397: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid397_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid397_Out0_copy398_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid397_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid397_Out0_copy398_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq500_uid400_bh7_uid401_In0_c0 <= "" & bh7_w86_1_c0 & bh7_w86_2_c0 & bh7_w86_3_c0 & bh7_w86_4_c0 & bh7_w86_5_c0;
   bh7_w86_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid401_Out0_c0(0);
   bh7_w87_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid401_Out0_c0(1);
   bh7_w88_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid401_Out0_c0(2);
   Compressor_5_3_Freq500_uid400_uid401: Compressor_5_3_Freq500_uid400
      port map ( X0 => Compressor_5_3_Freq500_uid400_bh7_uid401_In0_c0,
                 R => Compressor_5_3_Freq500_uid400_bh7_uid401_Out0_copy402_c0);
   Compressor_5_3_Freq500_uid400_bh7_uid401_Out0_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid401_Out0_copy402_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid403_In0_c0 <= "" & bh7_w87_1_c0 & bh7_w87_2_c0 & bh7_w87_3_c0 & bh7_w87_4_c0 & bh7_w87_5_c0 & bh7_w87_6_c0;
   bh7_w87_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid403_Out0_c0(0);
   bh7_w88_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid403_Out0_c0(1);
   bh7_w89_6_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid403_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid403: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid403_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid403_Out0_copy404_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid403_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid403_Out0_copy404_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid405_In0_c0 <= "" & bh7_w88_1_c0 & bh7_w88_2_c0 & bh7_w88_3_c0 & bh7_w88_4_c0 & bh7_w88_5_c0 & bh7_w88_6_c0;
   bh7_w88_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid405_Out0_c0(0);
   bh7_w89_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid405_Out0_c0(1);
   bh7_w90_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid405_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid405: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid405_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid405_Out0_copy406_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid405_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid405_Out0_copy406_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq500_uid400_bh7_uid407_In0_c0 <= "" & bh7_w89_1_c0 & bh7_w89_2_c0 & bh7_w89_3_c0 & bh7_w89_4_c0 & bh7_w89_5_c0;
   bh7_w89_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid407_Out0_c0(0);
   bh7_w90_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid407_Out0_c0(1);
   bh7_w91_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid407_Out0_c0(2);
   Compressor_5_3_Freq500_uid400_uid407: Compressor_5_3_Freq500_uid400
      port map ( X0 => Compressor_5_3_Freq500_uid400_bh7_uid407_In0_c0,
                 R => Compressor_5_3_Freq500_uid400_bh7_uid407_Out0_copy408_c0);
   Compressor_5_3_Freq500_uid400_bh7_uid407_Out0_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid407_Out0_copy408_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid409_In0_c0 <= "" & bh7_w90_1_c0 & bh7_w90_2_c0 & bh7_w90_3_c0 & bh7_w90_4_c0 & bh7_w90_5_c0 & bh7_w90_6_c0;
   bh7_w90_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid409_Out0_c0(0);
   bh7_w91_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid409_Out0_c0(1);
   bh7_w92_6_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid409_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid409: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid409_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid409_Out0_copy410_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid409_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid409_Out0_copy410_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid411_In0_c0 <= "" & bh7_w91_1_c0 & bh7_w91_2_c0 & bh7_w91_3_c0 & bh7_w91_4_c0 & bh7_w91_5_c0 & bh7_w91_6_c0;
   bh7_w91_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid411_Out0_c0(0);
   bh7_w92_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid411_Out0_c0(1);
   bh7_w93_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid411_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid411: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid411_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid411_Out0_copy412_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid411_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid411_Out0_copy412_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq500_uid400_bh7_uid413_In0_c0 <= "" & bh7_w92_1_c0 & bh7_w92_2_c0 & bh7_w92_3_c0 & bh7_w92_4_c0 & bh7_w92_5_c0;
   bh7_w92_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid413_Out0_c0(0);
   bh7_w93_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid413_Out0_c0(1);
   bh7_w94_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid413_Out0_c0(2);
   Compressor_5_3_Freq500_uid400_uid413: Compressor_5_3_Freq500_uid400
      port map ( X0 => Compressor_5_3_Freq500_uid400_bh7_uid413_In0_c0,
                 R => Compressor_5_3_Freq500_uid400_bh7_uid413_Out0_copy414_c0);
   Compressor_5_3_Freq500_uid400_bh7_uid413_Out0_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid413_Out0_copy414_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid415_In0_c0 <= "" & bh7_w93_1_c0 & bh7_w93_2_c0 & bh7_w93_3_c0 & bh7_w93_4_c0 & bh7_w93_5_c0 & bh7_w93_6_c0;
   bh7_w93_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid415_Out0_c0(0);
   bh7_w94_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid415_Out0_c0(1);
   bh7_w95_6_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid415_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid415: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid415_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid415_Out0_copy416_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid415_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid415_Out0_copy416_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid417_In0_c0 <= "" & bh7_w94_1_c0 & bh7_w94_2_c0 & bh7_w94_3_c0 & bh7_w94_4_c0 & bh7_w94_5_c0 & bh7_w94_6_c0;
   bh7_w94_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid417_Out0_c0(0);
   bh7_w95_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid417_Out0_c0(1);
   bh7_w96_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid417_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid417: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid417_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid417_Out0_copy418_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid417_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid417_Out0_copy418_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq500_uid400_bh7_uid419_In0_c0 <= "" & bh7_w95_1_c0 & bh7_w95_2_c0 & bh7_w95_3_c0 & bh7_w95_4_c0 & bh7_w95_5_c0;
   bh7_w95_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid419_Out0_c0(0);
   bh7_w96_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid419_Out0_c0(1);
   bh7_w97_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid419_Out0_c0(2);
   Compressor_5_3_Freq500_uid400_uid419: Compressor_5_3_Freq500_uid400
      port map ( X0 => Compressor_5_3_Freq500_uid400_bh7_uid419_In0_c0,
                 R => Compressor_5_3_Freq500_uid400_bh7_uid419_Out0_copy420_c0);
   Compressor_5_3_Freq500_uid400_bh7_uid419_Out0_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid419_Out0_copy420_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid421_In0_c0 <= "" & bh7_w96_1_c0 & bh7_w96_2_c0 & bh7_w96_3_c0 & bh7_w96_4_c0 & bh7_w96_5_c0 & bh7_w96_6_c0;
   bh7_w96_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid421_Out0_c0(0);
   bh7_w97_9_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid421_Out0_c0(1);
   bh7_w98_6_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid421_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid421: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid421_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid421_Out0_copy422_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid421_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid421_Out0_copy422_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid423_In0_c0 <= "" & bh7_w97_1_c0 & bh7_w97_2_c0 & bh7_w97_3_c0 & bh7_w97_4_c0 & bh7_w97_5_c0 & bh7_w97_6_c0;
   bh7_w97_10_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid423_Out0_c0(0);
   bh7_w98_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid423_Out0_c0(1);
   bh7_w99_6_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid423_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid423: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid423_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid423_Out0_copy424_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid423_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid423_Out0_copy424_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq500_uid400_bh7_uid425_In0_c0 <= "" & bh7_w98_1_c0 & bh7_w98_2_c0 & bh7_w98_3_c0 & bh7_w98_4_c0 & bh7_w98_5_c0;
   bh7_w98_8_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid425_Out0_c0(0);
   bh7_w99_7_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid425_Out0_c0(1);
   bh7_w100_6_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid425_Out0_c0(2);
   Compressor_5_3_Freq500_uid400_uid425: Compressor_5_3_Freq500_uid400
      port map ( X0 => Compressor_5_3_Freq500_uid400_bh7_uid425_In0_c0,
                 R => Compressor_5_3_Freq500_uid400_bh7_uid425_Out0_copy426_c0);
   Compressor_5_3_Freq500_uid400_bh7_uid425_Out0_c0 <= Compressor_5_3_Freq500_uid400_bh7_uid425_Out0_copy426_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid427_In0_c0 <= "" & bh7_w99_0_c0 & bh7_w99_1_c0 & bh7_w99_2_c0 & bh7_w99_3_c0 & bh7_w99_4_c0 & bh7_w99_5_c0;
   bh7_w99_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid427_Out0_c0(0);
   bh7_w100_7_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid427_Out0_c0(1);
   bh7_w101_3_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid427_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid427: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid427_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid427_Out0_copy428_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid427_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid427_Out0_copy428_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid429_In0_c0 <= "" & bh7_w100_0_c0 & bh7_w100_1_c0 & bh7_w100_2_c0 & bh7_w100_3_c0 & bh7_w100_4_c0 & bh7_w100_5_c0;
   bh7_w100_8_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid429_Out0_c0(0);
   bh7_w101_4_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid429_Out0_c0(1);
   bh7_w102_4_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid429_Out0_c0(2);
   Compressor_6_3_Freq500_uid334_uid429: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid429_In0_c0,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid429_Out0_copy430_c0);
   Compressor_6_3_Freq500_uid334_bh7_uid429_Out0_c0 <= Compressor_6_3_Freq500_uid334_bh7_uid429_Out0_copy430_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid433_In0_c0 <= "" & bh7_w101_0_c0 & bh7_w101_1_c0 & bh7_w101_2_c0;
   bh7_w101_5_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid433_Out0_c0(0);
   bh7_w102_5_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid433_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid433: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid433_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid433_Out0_copy434_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid433_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid433_Out0_copy434_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid435_In0_c0 <= "" & bh7_w102_0_c0 & bh7_w102_1_c0 & bh7_w102_2_c0 & bh7_w102_3_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid435_In1_c0 <= "" & bh7_w103_0_c0;
   bh7_w102_6_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid435_Out0_c0(0);
   bh7_w103_2_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid435_Out0_c0(1);
   bh7_w104_1_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid435_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid435: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid435_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid435_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid435_Out0_copy436_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid435_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid435_Out0_copy436_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid437_In0_c0 <= "" & bh7_w51_9_c0 & bh7_w51_8_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid437_In1_c0 <= "" & bh7_w52_10_c0 & bh7_w52_9_c0;
   bh7_w51_10_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid437_Out0_c0(0);
   bh7_w52_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid437_Out0_c0(1);
   bh7_w53_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid437_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid437: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid437_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid437_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid437_Out0_copy438_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid437_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid437_Out0_copy438_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid439_In0_c0 <= "" & bh7_w53_11_c0 & bh7_w53_10_c0 & bh7_w53_9_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid439_In1_c0 <= "" & bh7_w54_12_c0 & bh7_w54_11_c0;
   bh7_w53_13_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid439_Out0_c0(0);
   bh7_w54_14_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid439_Out0_c0(1);
   bh7_w55_13_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid439_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid439: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid439_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid439_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid439_Out0_copy440_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid439_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid439_Out0_copy440_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid441_In0_c0 <= "" & bh7_w55_10_c0 & bh7_w55_12_c0 & bh7_w55_11_c0;
   bh7_w55_14_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid441_Out0_c0(0);
   bh7_w56_12_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid441_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid441: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid441_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid441_Out0_copy442_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid441_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid441_Out0_copy442_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid443_In0_c0 <= "" & bh7_w56_8_c0 & bh7_w56_11_c0 & bh7_w56_10_c0 & bh7_w56_9_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid443_In1_c0 <= "" & "0";
   bh7_w56_13_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid443_Out0_c0(0);
   bh7_w57_14_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid443_Out0_c0(1);
   bh7_w58_13_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid443_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid443: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid443_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid443_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid443_Out0_copy444_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid443_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid443_Out0_copy444_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid445_In0_c0 <= "" & bh7_w57_12_c0 & bh7_w57_13_c0 & bh7_w57_11_c0;
   bh7_w57_15_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid445_Out0_c0(0);
   bh7_w58_14_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid445_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid445: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid445_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid445_Out0_copy446_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid445_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid445_Out0_copy446_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid447_In0_c0 <= "" & bh7_w58_10_c0 & bh7_w58_12_c0 & bh7_w58_11_c0;
   bh7_w58_15_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid447_Out0_c0(0);
   bh7_w59_12_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid447_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid447: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid447_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid447_Out0_copy448_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid447_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid447_Out0_copy448_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid449_In0_c0 <= "" & bh7_w59_8_c0 & bh7_w59_11_c0 & bh7_w59_10_c0 & bh7_w59_9_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid449_In1_c0 <= "" & "0";
   bh7_w59_13_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid449_Out0_c0(0);
   bh7_w60_14_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid449_Out0_c0(1);
   bh7_w61_13_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid449_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid449: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid449_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid449_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid449_Out0_copy450_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid449_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid449_Out0_copy450_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid451_In0_c0 <= "" & bh7_w60_12_c0 & bh7_w60_13_c0 & bh7_w60_11_c0;
   bh7_w60_15_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid451_Out0_c0(0);
   bh7_w61_14_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid451_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid451: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid451_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid451_Out0_copy452_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid451_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid451_Out0_copy452_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid453_In0_c0 <= "" & bh7_w61_10_c0 & bh7_w61_12_c0 & bh7_w61_11_c0;
   bh7_w61_15_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid453_Out0_c0(0);
   bh7_w62_12_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid453_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid453: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid453_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid453_Out0_copy454_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid453_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid453_Out0_copy454_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid455_In0_c0 <= "" & bh7_w62_8_c0 & bh7_w62_11_c0 & bh7_w62_10_c0 & bh7_w62_9_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid455_In1_c0 <= "" & "0";
   bh7_w62_13_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid455_Out0_c0(0);
   bh7_w63_14_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid455_Out0_c0(1);
   bh7_w64_13_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid455_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid455: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid455_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid455_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid455_Out0_copy456_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid455_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid455_Out0_copy456_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid457_In0_c0 <= "" & bh7_w63_12_c0 & bh7_w63_13_c0 & bh7_w63_11_c0;
   bh7_w63_15_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid457_Out0_c0(0);
   bh7_w64_14_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid457_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid457: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid457_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid457_Out0_copy458_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid457_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid457_Out0_copy458_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid459_In0_c0 <= "" & bh7_w64_10_c0 & bh7_w64_12_c0 & bh7_w64_11_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid459_In1_c0 <= "" & bh7_w65_11_c0 & bh7_w65_10_c0;
   bh7_w64_15_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid459_Out0_c0(0);
   bh7_w65_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid459_Out0_c0(1);
   bh7_w66_13_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid459_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid459: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid459_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid459_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid459_Out0_copy460_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid459_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid459_Out0_copy460_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid461_In0_c0 <= "" & bh7_w66_9_c0 & bh7_w66_12_c0 & bh7_w66_11_c0 & bh7_w66_10_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid461_In1_c0 <= "" & "0";
   bh7_w66_14_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid461_Out0_c0(0);
   bh7_w67_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid461_Out0_c0(1);
   bh7_w68_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid461_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid461: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid461_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid461_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid461_Out0_copy462_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid461_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid461_Out0_copy462_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid463_In0_c0 <= "" & bh7_w67_11_c0 & bh7_w67_10_c0 & bh7_w67_9_c0;
   bh7_w67_13_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid463_Out0_c0(0);
   bh7_w68_13_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid463_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid463: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid463_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid463_Out0_copy464_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid463_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid463_Out0_copy464_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid465_In0_c0 <= "" & bh7_w68_11_c0 & bh7_w68_10_c0 & bh7_w68_9_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid465_In1_c0 <= "" & bh7_w69_11_c0 & bh7_w69_10_c0;
   bh7_w68_14_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid465_Out0_c0(0);
   bh7_w69_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid465_Out0_c0(1);
   bh7_w70_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid465_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid465: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid465_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid465_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid465_Out0_copy466_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid465_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid465_Out0_copy466_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid467_In0_c0 <= "" & bh7_w70_11_c0 & bh7_w70_10_c0 & bh7_w70_9_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid467_In1_c0 <= "" & bh7_w71_11_c0 & bh7_w71_10_c0;
   bh7_w70_13_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid467_Out0_c0(0);
   bh7_w71_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid467_Out0_c0(1);
   bh7_w72_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid467_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid467: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid467_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid467_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid467_Out0_copy468_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid467_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid467_Out0_copy468_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid469_In0_c0 <= "" & bh7_w72_11_c0 & bh7_w72_10_c0 & bh7_w72_9_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid469_In1_c0 <= "" & bh7_w73_11_c0 & bh7_w73_10_c0;
   bh7_w72_13_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid469_Out0_c0(0);
   bh7_w73_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid469_Out0_c0(1);
   bh7_w74_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid469_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid469: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid469_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid469_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid469_Out0_copy470_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid469_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid469_Out0_copy470_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid471_In0_c0 <= "" & bh7_w74_11_c0 & bh7_w74_10_c0 & bh7_w74_9_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid471_In1_c0 <= "" & bh7_w75_10_c0 & bh7_w75_9_c0;
   bh7_w74_13_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid471_Out0_c0(0);
   bh7_w75_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid471_Out0_c0(1);
   bh7_w76_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid471_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid471: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid471_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid471_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid471_Out0_copy472_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid471_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid471_Out0_copy472_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid473_In0_c0 <= "" & bh7_w76_10_c0 & bh7_w76_9_c0 & bh7_w76_8_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid473_In1_c0 <= "" & bh7_w77_10_c0 & bh7_w77_9_c0;
   bh7_w76_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid473_Out0_c0(0);
   bh7_w77_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid473_Out0_c0(1);
   bh7_w78_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid473_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid473: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid473_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid473_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid473_Out0_copy474_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid473_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid473_Out0_copy474_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid475_In0_c0 <= "" & bh7_w78_10_c0 & bh7_w78_9_c0 & bh7_w78_8_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid475_In1_c0 <= "" & bh7_w79_10_c0 & bh7_w79_9_c0;
   bh7_w78_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid475_Out0_c0(0);
   bh7_w79_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid475_Out0_c0(1);
   bh7_w80_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid475_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid475: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid475_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid475_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid475_Out0_copy476_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid475_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid475_Out0_copy476_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid477_In0_c0 <= "" & bh7_w80_10_c0 & bh7_w80_9_c0 & bh7_w80_8_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid477_In1_c0 <= "" & bh7_w81_10_c0 & bh7_w81_9_c0;
   bh7_w80_12_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid477_Out0_c0(0);
   bh7_w81_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid477_Out0_c0(1);
   bh7_w82_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid477_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid477: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid477_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid477_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid477_Out0_copy478_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid477_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid477_Out0_copy478_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid479_In0_c0 <= "" & bh7_w82_7_c0 & bh7_w82_10_c0 & bh7_w82_9_c0 & bh7_w82_8_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid479_In1_c0 <= "" & "0";
   bh7_w82_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid479_Out0_c0(0);
   bh7_w83_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid479_Out0_c0(1);
   bh7_w84_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid479_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid479: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid479_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid479_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid479_Out0_copy480_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid479_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid479_Out0_copy480_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid481_In0_c0 <= "" & bh7_w83_9_c0 & bh7_w83_8_c0 & bh7_w83_7_c0;
   bh7_w83_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid481_Out0_c0(0);
   bh7_w84_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid481_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid481: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid481_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid481_Out0_copy482_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid481_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid481_Out0_copy482_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid483_In0_c0 <= "" & bh7_w84_9_c0 & bh7_w84_8_c0 & bh7_w84_7_c0;
   bh7_w84_12_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid483_Out0_c0(0);
   bh7_w85_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid483_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid483: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid483_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid483_Out0_copy484_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid483_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid483_Out0_copy484_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid485_In0_c0 <= "" & bh7_w85_7_c0 & bh7_w85_10_c0 & bh7_w85_9_c0 & bh7_w85_8_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid485_In1_c0 <= "" & "0";
   bh7_w85_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid485_Out0_c0(0);
   bh7_w86_9_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid485_Out0_c0(1);
   bh7_w87_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid485_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid485: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid485_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid485_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid485_Out0_copy486_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid485_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid485_Out0_copy486_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid487_In0_c0 <= "" & bh7_w86_8_c0 & bh7_w86_7_c0 & bh7_w86_6_c0;
   bh7_w86_10_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid487_Out0_c0(0);
   bh7_w87_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid487_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid487: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid487_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid487_Out0_copy488_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid487_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid487_Out0_copy488_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid489_In0_c0 <= "" & bh7_w87_8_c0 & bh7_w87_9_c0 & bh7_w87_7_c0;
   bh7_w87_12_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid489_Out0_c0(0);
   bh7_w88_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid489_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid489: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid489_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid489_Out0_copy490_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid489_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid489_Out0_copy490_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid491_In0_c0 <= "" & bh7_w88_7_c0 & bh7_w88_8_c0 & bh7_w88_10_c0 & bh7_w88_9_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid491_In1_c0 <= "" & "0";
   bh7_w88_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid491_Out0_c0(0);
   bh7_w89_9_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid491_Out0_c0(1);
   bh7_w90_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid491_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid491: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid491_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid491_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid491_Out0_copy492_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid491_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid491_Out0_copy492_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid493_In0_c0 <= "" & bh7_w89_8_c0 & bh7_w89_7_c0 & bh7_w89_6_c0;
   bh7_w89_10_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid493_Out0_c0(0);
   bh7_w90_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid493_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid493: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid493_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid493_Out0_copy494_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid493_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid493_Out0_copy494_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid495_In0_c0 <= "" & bh7_w90_8_c0 & bh7_w90_9_c0 & bh7_w90_7_c0;
   bh7_w90_12_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid495_Out0_c0(0);
   bh7_w91_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid495_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid495: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid495_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid495_Out0_copy496_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid495_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid495_Out0_copy496_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid497_In0_c0 <= "" & bh7_w91_7_c0 & bh7_w91_8_c0 & bh7_w91_10_c0 & bh7_w91_9_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid497_In1_c0 <= "" & "0";
   bh7_w91_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid497_Out0_c0(0);
   bh7_w92_9_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid497_Out0_c0(1);
   bh7_w93_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid497_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid497: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid497_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid497_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid497_Out0_copy498_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid497_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid497_Out0_copy498_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid499_In0_c0 <= "" & bh7_w92_8_c0 & bh7_w92_7_c0 & bh7_w92_6_c0;
   bh7_w92_10_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid499_Out0_c0(0);
   bh7_w93_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid499_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid499: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid499_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid499_Out0_copy500_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid499_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid499_Out0_copy500_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid501_In0_c0 <= "" & bh7_w93_8_c0 & bh7_w93_9_c0 & bh7_w93_7_c0;
   bh7_w93_12_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid501_Out0_c0(0);
   bh7_w94_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid501_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid501: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid501_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid501_Out0_copy502_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid501_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid501_Out0_copy502_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid503_In0_c0 <= "" & bh7_w94_7_c0 & bh7_w94_8_c0 & bh7_w94_10_c0 & bh7_w94_9_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid503_In1_c0 <= "" & "0";
   bh7_w94_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid503_Out0_c0(0);
   bh7_w95_9_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid503_Out0_c0(1);
   bh7_w96_10_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid503_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid503: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid503_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid503_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid503_Out0_copy504_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid503_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid503_Out0_copy504_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid505_In0_c0 <= "" & bh7_w95_8_c0 & bh7_w95_7_c0 & bh7_w95_6_c0;
   bh7_w95_10_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid505_Out0_c0(0);
   bh7_w96_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid505_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid505: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid505_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid505_Out0_copy506_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid505_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid505_Out0_copy506_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid507_In0_c0 <= "" & bh7_w96_8_c0 & bh7_w96_9_c0 & bh7_w96_7_c0;
   bh7_w96_12_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid507_Out0_c0(0);
   bh7_w97_11_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid507_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid507: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid507_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid507_Out0_copy508_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid507_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid507_Out0_copy508_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid509_In0_c0 <= "" & bh7_w97_7_c0 & bh7_w97_8_c0 & bh7_w97_10_c0 & bh7_w97_9_c0;
   Compressor_14_3_Freq500_uid326_bh7_uid509_In1_c0 <= "" & "0";
   bh7_w97_12_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid509_Out0_c0(0);
   bh7_w98_9_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid509_Out0_c0(1);
   bh7_w99_9_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid509_Out0_c0(2);
   Compressor_14_3_Freq500_uid326_uid509: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid509_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid509_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid509_Out0_copy510_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid509_Out0_c0 <= Compressor_14_3_Freq500_uid326_bh7_uid509_Out0_copy510_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid511_In0_c0 <= "" & bh7_w98_8_c0 & bh7_w98_7_c0 & bh7_w98_6_c0;
   bh7_w98_10_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid511_Out0_c0(0);
   bh7_w99_10_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid511_Out0_c0(1);
   Compressor_3_2_Freq500_uid432_uid511: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid511_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid511_Out0_copy512_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid511_Out0_c0 <= Compressor_3_2_Freq500_uid432_bh7_uid511_Out0_copy512_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid513_In0_c0 <= "" & bh7_w99_7_c0 & bh7_w99_8_c0 & bh7_w99_6_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid513_In1_c0 <= "" & bh7_w100_6_c0 & bh7_w100_8_c0;
   bh7_w99_11_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid513_Out0_c0(0);
   bh7_w100_9_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid513_Out0_c0(1);
   bh7_w101_6_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid513_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid513: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid513_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid513_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid513_Out0_copy514_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid513_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid513_Out0_copy514_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid515_In0_c0 <= "" & bh7_w101_5_c0 & bh7_w101_4_c0 & bh7_w101_3_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid515_In1_c0 <= "" & bh7_w102_6_c0 & bh7_w102_5_c0;
   bh7_w101_7_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid515_Out0_c0(0);
   bh7_w102_7_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid515_Out0_c0(1);
   bh7_w103_3_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid515_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid515: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid515_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid515_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid515_Out0_copy516_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid515_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid515_Out0_copy516_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid517_In0_c0 <= "" & bh7_w103_1_c0 & bh7_w103_2_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid517_In1_c0 <= "" & bh7_w104_0_c0 & bh7_w104_1_c0;
   bh7_w103_4_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid517_Out0_c0(0);
   bh7_w104_2_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid517_Out0_c0(1);
   bh7_w105_1_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid517_Out0_c0(2);
   Compressor_23_3_Freq500_uid322_uid517: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid517_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid517_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid517_Out0_copy518_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid517_Out0_c0 <= Compressor_23_3_Freq500_uid322_bh7_uid517_Out0_copy518_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid519_In0_c0 <= "" & bh7_w53_13_c0 & bh7_w53_12_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid519_In1_c0 <= "" & bh7_w54_13_c0 & bh7_w54_14_c0;
   bh7_w53_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_c1(0);
   bh7_w54_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_c1(1);
   bh7_w55_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid519: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid519_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid519_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_copy520_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid519_Out0_copy520_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid521_In0_c0 <= "" & bh7_w55_13_c0 & bh7_w55_14_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid521_In1_c0 <= "" & bh7_w56_13_c0 & bh7_w56_12_c0;
   bh7_w55_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_c1(0);
   bh7_w56_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_c1(1);
   bh7_w57_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid521: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid521_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid521_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_copy522_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid521_Out0_copy522_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid523_In0_c0 <= "" & bh7_w57_14_c0 & bh7_w57_15_c0 & "0";
   bh7_w57_17_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_c1(0);
   bh7_w58_16_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid523: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid523_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_copy524_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid523_Out0_copy524_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid525_In0_c0 <= "" & bh7_w58_13_c0 & bh7_w58_15_c0 & bh7_w58_14_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid525_In1_c0 <= "" & bh7_w59_13_c0 & bh7_w59_12_c0;
   bh7_w58_17_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_c1(0);
   bh7_w59_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_c1(1);
   bh7_w60_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid525: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid525_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid525_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_copy526_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid525_Out0_copy526_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid527_In0_c0 <= "" & bh7_w60_14_c0 & bh7_w60_15_c0 & "0";
   bh7_w60_17_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_c1(0);
   bh7_w61_16_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid527: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid527_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_copy528_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid527_Out0_copy528_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid529_In0_c0 <= "" & bh7_w61_13_c0 & bh7_w61_15_c0 & bh7_w61_14_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid529_In1_c0 <= "" & bh7_w62_13_c0 & bh7_w62_12_c0;
   bh7_w61_17_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_c1(0);
   bh7_w62_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_c1(1);
   bh7_w63_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid529: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid529_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid529_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_copy530_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid529_Out0_copy530_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid531_In0_c0 <= "" & bh7_w63_14_c0 & bh7_w63_15_c0 & "0";
   bh7_w63_17_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_c1(0);
   bh7_w64_16_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid531: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid531_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_copy532_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid531_Out0_copy532_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid533_In0_c0 <= "" & bh7_w64_13_c0 & bh7_w64_15_c0 & bh7_w64_14_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid533_In1_c0 <= "" & bh7_w65_9_c0 & bh7_w65_12_c0;
   bh7_w64_17_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_c1(0);
   bh7_w65_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_c1(1);
   bh7_w66_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid533: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid533_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid533_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_copy534_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid533_Out0_copy534_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid535_In0_c0 <= "" & bh7_w66_14_c0 & bh7_w66_13_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid535_In1_c0 <= "" & bh7_w67_12_c0 & bh7_w67_13_c0;
   bh7_w66_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_c1(0);
   bh7_w67_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_c1(1);
   bh7_w68_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid535: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid535_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid535_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_copy536_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid535_Out0_copy536_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid537_In0_c0 <= "" & bh7_w68_12_c0 & bh7_w68_14_c0 & bh7_w68_13_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid537_In1_c0 <= "" & bh7_w69_9_c0 & bh7_w69_12_c0;
   bh7_w68_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_c1(0);
   bh7_w69_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_c1(1);
   bh7_w70_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid537: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid537_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid537_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_copy538_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid537_Out0_copy538_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid539_In0_c0 <= "" & bh7_w70_13_c0 & bh7_w70_12_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid539_In1_c0 <= "" & bh7_w71_9_c0 & bh7_w71_12_c0;
   bh7_w70_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_c1(0);
   bh7_w71_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_c1(1);
   bh7_w72_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid539: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid539_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid539_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_copy540_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid539_Out0_copy540_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid541_In0_c0 <= "" & bh7_w72_13_c0 & bh7_w72_12_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid541_In1_c0 <= "" & bh7_w73_9_c0 & bh7_w73_12_c0;
   bh7_w72_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_c1(0);
   bh7_w73_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_c1(1);
   bh7_w74_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid541: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid541_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid541_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_copy542_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid541_Out0_copy542_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid543_In0_c0 <= "" & bh7_w74_13_c0 & bh7_w74_12_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid543_In1_c0 <= "" & bh7_w75_8_c0 & bh7_w75_11_c0;
   bh7_w74_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_c1(0);
   bh7_w75_12_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_c1(1);
   bh7_w76_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid543: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid543_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid543_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_copy544_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid543_Out0_copy544_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid545_In0_c0 <= "" & bh7_w76_12_c0 & bh7_w76_11_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid545_In1_c0 <= "" & bh7_w77_8_c0 & bh7_w77_11_c0;
   bh7_w76_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_c1(0);
   bh7_w77_12_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_c1(1);
   bh7_w78_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid545: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid545_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid545_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_copy546_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid545_Out0_copy546_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid547_In0_c0 <= "" & bh7_w78_12_c0 & bh7_w78_11_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid547_In1_c0 <= "" & bh7_w79_8_c0 & bh7_w79_11_c0;
   bh7_w78_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_c1(0);
   bh7_w79_12_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_c1(1);
   bh7_w80_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid547: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid547_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid547_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_copy548_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid547_Out0_copy548_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid549_In0_c0 <= "" & bh7_w80_12_c0 & bh7_w80_11_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid549_In1_c0 <= "" & bh7_w81_8_c0 & bh7_w81_11_c0;
   bh7_w80_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_c1(0);
   bh7_w81_12_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_c1(1);
   bh7_w82_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid549: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid549_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid549_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_copy550_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid549_Out0_copy550_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid551_In0_c0 <= "" & bh7_w82_12_c0 & bh7_w82_11_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid551_In1_c0 <= "" & bh7_w83_10_c0 & bh7_w83_11_c0;
   bh7_w82_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_c1(0);
   bh7_w83_12_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_c1(1);
   bh7_w84_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid551: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid551_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid551_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_copy552_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid551_Out0_copy552_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid553_In0_c0 <= "" & bh7_w84_10_c0 & bh7_w84_12_c0 & bh7_w84_11_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid553_In1_c0 <= "" & bh7_w85_12_c0 & bh7_w85_11_c0;
   bh7_w84_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_c1(0);
   bh7_w85_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_c1(1);
   bh7_w86_11_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid553: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid553_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid553_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_copy554_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid553_Out0_copy554_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid555_In0_c0 <= "" & bh7_w86_9_c0 & bh7_w86_10_c0 & "0";
   bh7_w86_12_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_c1(0);
   bh7_w87_13_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid555: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid555_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_copy556_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid555_Out0_copy556_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid557_In0_c0 <= "" & bh7_w87_10_c0 & bh7_w87_12_c0 & bh7_w87_11_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid557_In1_c0 <= "" & bh7_w88_12_c0 & bh7_w88_11_c0;
   bh7_w87_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_c1(0);
   bh7_w88_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_c1(1);
   bh7_w89_11_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid557: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid557_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid557_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_copy558_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid557_Out0_copy558_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid559_In0_c0 <= "" & bh7_w89_9_c0 & bh7_w89_10_c0 & "0";
   bh7_w89_12_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_c1(0);
   bh7_w90_13_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid559: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid559_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_copy560_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid559_Out0_copy560_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid561_In0_c0 <= "" & bh7_w90_10_c0 & bh7_w90_12_c0 & bh7_w90_11_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid561_In1_c0 <= "" & bh7_w91_12_c0 & bh7_w91_11_c0;
   bh7_w90_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_c1(0);
   bh7_w91_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_c1(1);
   bh7_w92_11_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid561: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid561_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid561_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_copy562_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid561_Out0_copy562_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid563_In0_c0 <= "" & bh7_w92_9_c0 & bh7_w92_10_c0 & "0";
   bh7_w92_12_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_c1(0);
   bh7_w93_13_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid563: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid563_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_copy564_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid563_Out0_copy564_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid565_In0_c0 <= "" & bh7_w93_10_c0 & bh7_w93_12_c0 & bh7_w93_11_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid565_In1_c0 <= "" & bh7_w94_12_c0 & bh7_w94_11_c0;
   bh7_w93_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_c1(0);
   bh7_w94_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_c1(1);
   bh7_w95_11_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid565: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid565_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid565_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_copy566_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid565_Out0_copy566_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid567_In0_c0 <= "" & bh7_w95_9_c0 & bh7_w95_10_c0 & "0";
   bh7_w95_12_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_c1(0);
   bh7_w96_13_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid567: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid567_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_copy568_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid567_Out0_copy568_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid569_In0_c0 <= "" & bh7_w96_10_c0 & bh7_w96_12_c0 & bh7_w96_11_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid569_In1_c0 <= "" & bh7_w97_12_c0 & bh7_w97_11_c0;
   bh7_w96_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_c1(0);
   bh7_w97_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_c1(1);
   bh7_w98_11_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid569: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid569_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid569_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_copy570_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid569_Out0_copy570_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid571_In0_c0 <= "" & bh7_w98_9_c0 & bh7_w98_10_c0 & "0";
   bh7_w98_12_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_c1(0);
   bh7_w99_12_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid571: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid571_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_copy572_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid571_Out0_copy572_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid573_In0_c0 <= "" & bh7_w99_9_c0 & bh7_w99_11_c0 & bh7_w99_10_c0;
   Compressor_23_3_Freq500_uid322_bh7_uid573_In1_c0 <= "" & bh7_w100_7_c0 & bh7_w100_9_c0;
   bh7_w99_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_c1(0);
   bh7_w100_10_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_c1(1);
   bh7_w101_8_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid573: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid573_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid573_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_copy574_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid573_Out0_copy574_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid575_In0_c0 <= "" & bh7_w101_7_c0 & bh7_w101_6_c0 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid575_In1_c0 <= "" & bh7_w102_4_c0 & bh7_w102_7_c0;
   bh7_w101_9_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_c1(0);
   bh7_w102_8_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_c1(1);
   bh7_w103_5_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid575: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid575_In0_c0,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid575_In1_c0,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_copy576_c0);
   Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid575_Out0_copy576_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid577_In0_c0 <= "" & bh7_w103_4_c0 & bh7_w103_3_c0 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid577_In1_c0 <= "" & bh7_w104_2_c0;
   bh7_w103_6_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_c1(0);
   bh7_w104_3_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_c1(1);
   bh7_w105_2_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid577: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid577_In0_c0,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid577_In1_c0,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_copy578_c0);
   Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid577_Out0_copy578_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid579_In0_c0 <= "" & bh7_w105_0_c0 & bh7_w105_1_c0 & "0";
   bh7_w105_3_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid579_Out0_c1(0);
   Compressor_3_2_Freq500_uid432_uid579: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid579_In0_c0,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid579_Out0_copy580_c0);
   Compressor_3_2_Freq500_uid432_bh7_uid579_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid579_Out0_copy580_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid581_In0_c1 <= "" & bh7_w55_16_c1 & bh7_w55_15_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid581_In1_c1 <= "" & bh7_w56_14_c1;
   bh7_w55_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid581_Out0_c1(0);
   bh7_w56_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid581_Out0_c1(1);
   bh7_w57_18_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid581_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid581: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid581_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid581_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid581_Out0_copy582_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid581_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid581_Out0_copy582_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid583_In0_c1 <= "" & bh7_w57_16_c1 & bh7_w57_17_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid583_In1_c1 <= "" & bh7_w58_16_c1 & bh7_w58_17_c1;
   bh7_w57_19_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid583_Out0_c1(0);
   bh7_w58_18_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid583_Out0_c1(1);
   bh7_w59_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid583_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid583: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid583_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid583_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid583_Out0_copy584_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid583_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid583_Out0_copy584_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid585_In0_c1 <= "" & bh7_w60_16_c1 & bh7_w60_17_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid585_In1_c1 <= "" & bh7_w61_16_c1 & bh7_w61_17_c1;
   bh7_w60_18_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid585_Out0_c1(0);
   bh7_w61_18_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid585_Out0_c1(1);
   bh7_w62_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid585_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid585: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid585_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid585_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid585_Out0_copy586_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid585_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid585_Out0_copy586_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid587_In0_c1 <= "" & bh7_w63_16_c1 & bh7_w63_17_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid587_In1_c1 <= "" & bh7_w64_16_c1 & bh7_w64_17_c1;
   bh7_w63_18_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid587_Out0_c1(0);
   bh7_w64_18_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid587_Out0_c1(1);
   bh7_w65_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid587_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid587: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid587_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid587_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid587_Out0_copy588_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid587_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid587_Out0_copy588_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid589_In0_c1 <= "" & bh7_w66_15_c1 & bh7_w66_16_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid589_In1_c1 <= "" & bh7_w67_14_c1;
   bh7_w66_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid589_Out0_c1(0);
   bh7_w67_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid589_Out0_c1(1);
   bh7_w68_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid589_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid589: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid589_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid589_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid589_Out0_copy590_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid589_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid589_Out0_copy590_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid591_In0_c1 <= "" & bh7_w68_15_c1 & bh7_w68_16_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid591_In1_c1 <= "" & bh7_w69_13_c1;
   bh7_w68_18_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid591_Out0_c1(0);
   bh7_w69_14_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid591_Out0_c1(1);
   bh7_w70_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid591_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid591: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid591_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid591_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid591_Out0_copy592_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid591_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid591_Out0_copy592_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid593_In0_c1 <= "" & bh7_w70_14_c1 & bh7_w70_15_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid593_In1_c1 <= "" & bh7_w71_13_c1;
   bh7_w70_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid593_Out0_c1(0);
   bh7_w71_14_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid593_Out0_c1(1);
   bh7_w72_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid593_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid593: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid593_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid593_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid593_Out0_copy594_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid593_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid593_Out0_copy594_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid595_In0_c1 <= "" & bh7_w72_15_c1 & bh7_w72_14_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid595_In1_c1 <= "" & bh7_w73_13_c1;
   bh7_w72_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid595_Out0_c1(0);
   bh7_w73_14_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid595_Out0_c1(1);
   bh7_w74_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid595_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid595: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid595_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid595_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid595_Out0_copy596_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid595_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid595_Out0_copy596_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid597_In0_c1 <= "" & bh7_w74_15_c1 & bh7_w74_14_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid597_In1_c1 <= "" & bh7_w75_12_c1;
   bh7_w74_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid597_Out0_c1(0);
   bh7_w75_13_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid597_Out0_c1(1);
   bh7_w76_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid597_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid597: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid597_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid597_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid597_Out0_copy598_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid597_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid597_Out0_copy598_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid599_In0_c1 <= "" & bh7_w76_14_c1 & bh7_w76_13_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid599_In1_c1 <= "" & bh7_w77_12_c1;
   bh7_w76_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid599_Out0_c1(0);
   bh7_w77_13_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid599_Out0_c1(1);
   bh7_w78_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid599_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid599: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid599_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid599_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid599_Out0_copy600_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid599_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid599_Out0_copy600_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid601_In0_c1 <= "" & bh7_w78_14_c1 & bh7_w78_13_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid601_In1_c1 <= "" & bh7_w79_12_c1;
   bh7_w78_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid601_Out0_c1(0);
   bh7_w79_13_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid601_Out0_c1(1);
   bh7_w80_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid601_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid601: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid601_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid601_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid601_Out0_copy602_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid601_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid601_Out0_copy602_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid603_In0_c1 <= "" & bh7_w80_14_c1 & bh7_w80_13_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid603_In1_c1 <= "" & bh7_w81_12_c1;
   bh7_w80_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid603_Out0_c1(0);
   bh7_w81_13_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid603_Out0_c1(1);
   bh7_w82_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid603_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid603: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid603_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid603_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid603_Out0_copy604_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid603_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid603_Out0_copy604_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid605_In0_c1 <= "" & bh7_w82_14_c1 & bh7_w82_13_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid605_In1_c1 <= "" & bh7_w83_12_c1;
   bh7_w82_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid605_Out0_c1(0);
   bh7_w83_13_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid605_Out0_c1(1);
   bh7_w84_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid605_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid605: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid605_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid605_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid605_Out0_copy606_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid605_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid605_Out0_copy606_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid607_In0_c1 <= "" & bh7_w84_13_c1 & bh7_w84_14_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid607_In1_c1 <= "" & bh7_w85_13_c1;
   bh7_w84_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid607_Out0_c1(0);
   bh7_w85_14_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid607_Out0_c1(1);
   bh7_w86_13_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid607_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid607: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid607_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid607_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid607_Out0_copy608_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid607_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid607_Out0_copy608_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid609_In0_c1 <= "" & bh7_w86_11_c1 & bh7_w86_12_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid609_In1_c1 <= "" & bh7_w87_13_c1 & bh7_w87_14_c1;
   bh7_w86_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid609_Out0_c1(0);
   bh7_w87_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid609_Out0_c1(1);
   bh7_w88_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid609_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid609: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid609_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid609_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid609_Out0_copy610_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid609_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid609_Out0_copy610_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid611_In0_c1 <= "" & bh7_w89_11_c1 & bh7_w89_12_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid611_In1_c1 <= "" & bh7_w90_13_c1 & bh7_w90_14_c1;
   bh7_w89_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid611_Out0_c1(0);
   bh7_w90_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid611_Out0_c1(1);
   bh7_w91_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid611_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid611: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid611_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid611_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid611_Out0_copy612_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid611_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid611_Out0_copy612_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid613_In0_c1 <= "" & bh7_w92_11_c1 & bh7_w92_12_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid613_In1_c1 <= "" & bh7_w93_13_c1 & bh7_w93_14_c1;
   bh7_w92_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid613_Out0_c1(0);
   bh7_w93_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid613_Out0_c1(1);
   bh7_w94_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid613_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid613: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid613_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid613_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid613_Out0_copy614_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid613_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid613_Out0_copy614_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid615_In0_c1 <= "" & bh7_w95_11_c1 & bh7_w95_12_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid615_In1_c1 <= "" & bh7_w96_13_c1 & bh7_w96_14_c1;
   bh7_w95_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid615_Out0_c1(0);
   bh7_w96_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid615_Out0_c1(1);
   bh7_w97_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid615_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid615: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid615_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid615_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid615_Out0_copy616_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid615_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid615_Out0_copy616_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid617_In0_c1 <= "" & bh7_w98_11_c1 & bh7_w98_12_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid617_In1_c1 <= "" & bh7_w99_12_c1 & bh7_w99_13_c1;
   bh7_w98_13_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid617_Out0_c1(0);
   bh7_w99_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid617_Out0_c1(1);
   bh7_w100_11_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid617_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid617: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid617_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid617_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid617_Out0_copy618_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid617_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid617_Out0_copy618_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid619_In0_c1 <= "" & bh7_w101_8_c1 & bh7_w101_9_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid619_In1_c1 <= "" & bh7_w102_8_c1;
   bh7_w101_10_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid619_Out0_c1(0);
   bh7_w102_9_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid619_Out0_c1(1);
   bh7_w103_7_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid619_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid619: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid619_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid619_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid619_Out0_copy620_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid619_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid619_Out0_copy620_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid621_In0_c1 <= "" & bh7_w103_6_c1 & bh7_w103_5_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid621_In1_c1 <= "" & bh7_w104_3_c1;
   bh7_w103_8_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid621_Out0_c1(0);
   bh7_w104_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid621_Out0_c1(1);
   bh7_w105_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid621_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid621: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid621_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid621_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid621_Out0_copy622_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid621_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid621_Out0_copy622_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid623_In0_c1 <= "" & bh7_w105_3_c1 & bh7_w105_2_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid623_In1_c0 <= "" & "0";
   bh7_w105_5_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid623_Out0_c1(0);
   Compressor_14_3_Freq500_uid326_uid623: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid623_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid623_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid623_Out0_copy624_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid623_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid623_Out0_copy624_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid625_In0_c1 <= "" & bh7_w17_0_c1 & bh7_w17_1_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid625_In1_c1 <= "" & bh7_w18_0_c1 & bh7_w18_1_c1;
   bh7_w17_2_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid625_Out0_c1(0);
   bh7_w18_2_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid625_Out0_c1(1);
   bh7_w19_2_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid625_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid625: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid625_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid625_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid625_Out0_copy626_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid625_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid625_Out0_copy626_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid627_In0_c1 <= "" & bh7_w19_0_c1 & bh7_w19_1_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid627_In1_c1 <= "" & bh7_w20_0_c1 & bh7_w20_1_c1;
   bh7_w19_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid627_Out0_c1(0);
   bh7_w20_2_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid627_Out0_c1(1);
   bh7_w21_2_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid627_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid627: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid627_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid627_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid627_Out0_copy628_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid627_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid627_Out0_copy628_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid629_In0_c1 <= "" & bh7_w21_0_c1 & bh7_w21_1_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid629_In1_c1 <= "" & bh7_w22_0_c1 & bh7_w22_1_c1;
   bh7_w21_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid629_Out0_c1(0);
   bh7_w22_2_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid629_Out0_c1(1);
   bh7_w23_2_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid629_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid629: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid629_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid629_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid629_Out0_copy630_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid629_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid629_Out0_copy630_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid631_In0_c1 <= "" & bh7_w23_0_c1 & bh7_w23_1_c1 & "0";
   bh7_w23_3_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid631_Out0_c1(0);
   bh7_w24_3_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid631_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid631: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid631_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid631_Out0_copy632_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid631_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid631_Out0_copy632_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid633_In0_c1 <= "" & bh7_w24_0_c1 & bh7_w24_1_c1 & bh7_w24_2_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid633_In1_c1 <= "" & bh7_w25_0_c1 & bh7_w25_1_c1;
   bh7_w24_4_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid633_Out0_c1(0);
   bh7_w25_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid633_Out0_c1(1);
   bh7_w26_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid633_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid633: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid633_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid633_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid633_Out0_copy634_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid633_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid633_Out0_copy634_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid635_In0_c1 <= "" & bh7_w26_0_c1 & bh7_w26_1_c1 & bh7_w26_2_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid635_In1_c1 <= "" & bh7_w27_0_c1 & bh7_w27_1_c1;
   bh7_w26_4_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid635_Out0_c1(0);
   bh7_w27_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid635_Out0_c1(1);
   bh7_w28_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid635_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid635: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid635_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid635_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid635_Out0_copy636_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid635_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid635_Out0_copy636_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid637_In0_c1 <= "" & bh7_w28_0_c1 & bh7_w28_1_c1 & bh7_w28_2_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid637_In1_c1 <= "" & bh7_w29_0_c1 & bh7_w29_1_c1;
   bh7_w28_4_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid637_Out0_c1(0);
   bh7_w29_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid637_Out0_c1(1);
   bh7_w30_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid637_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid637: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid637_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid637_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid637_Out0_copy638_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid637_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid637_Out0_copy638_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid639_In0_c1 <= "" & bh7_w30_0_c1 & bh7_w30_1_c1 & bh7_w30_2_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid639_In1_c1 <= "" & bh7_w31_0_c1 & bh7_w31_1_c1;
   bh7_w30_4_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid639_Out0_c1(0);
   bh7_w31_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid639_Out0_c1(1);
   bh7_w32_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid639_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid639: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid639_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid639_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid639_Out0_copy640_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid639_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid639_Out0_copy640_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid641_In0_c1 <= "" & bh7_w32_0_c1 & bh7_w32_1_c1 & bh7_w32_2_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid641_In1_c1 <= "" & bh7_w33_0_c1 & bh7_w33_1_c1;
   bh7_w32_4_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid641_Out0_c1(0);
   bh7_w33_3_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid641_Out0_c1(1);
   bh7_w34_4_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid641_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid641: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid641_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid641_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid641_Out0_copy642_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid641_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid641_Out0_copy642_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid643_In0_c1 <= "" & bh7_w34_0_c1 & bh7_w34_1_c1 & bh7_w34_2_c1 & bh7_w34_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid643_In1_c1 <= "" & bh7_w35_0_c1;
   bh7_w34_5_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid643_Out0_c1(0);
   bh7_w35_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid643_Out0_c1(1);
   bh7_w36_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid643_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid643: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid643_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid643_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid643_Out0_copy644_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid643_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid643_Out0_copy644_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid645_In0_c1 <= "" & bh7_w35_1_c1 & bh7_w35_2_c1 & bh7_w35_3_c1;
   bh7_w35_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid645_Out0_c1(0);
   bh7_w36_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid645_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid645: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid645_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid645_Out0_copy646_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid645_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid645_Out0_copy646_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid647_In0_c1 <= "" & bh7_w36_0_c1 & bh7_w36_1_c1 & bh7_w36_2_c1 & bh7_w36_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid647_In1_c1 <= "" & bh7_w37_0_c1;
   bh7_w36_6_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid647_Out0_c1(0);
   bh7_w37_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid647_Out0_c1(1);
   bh7_w38_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid647_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid647: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid647_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid647_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid647_Out0_copy648_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid647_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid647_Out0_copy648_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid649_In0_c1 <= "" & bh7_w37_1_c1 & bh7_w37_2_c1 & bh7_w37_3_c1;
   bh7_w37_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid649_Out0_c1(0);
   bh7_w38_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid649_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid649: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid649_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid649_Out0_copy650_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid649_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid649_Out0_copy650_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid651_In0_c1 <= "" & bh7_w38_0_c1 & bh7_w38_1_c1 & bh7_w38_2_c1 & bh7_w38_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid651_In1_c1 <= "" & bh7_w39_0_c1;
   bh7_w38_6_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid651_Out0_c1(0);
   bh7_w39_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid651_Out0_c1(1);
   bh7_w40_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid651_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid651: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid651_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid651_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid651_Out0_copy652_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid651_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid651_Out0_copy652_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid653_In0_c1 <= "" & bh7_w39_1_c1 & bh7_w39_2_c1 & bh7_w39_3_c1;
   bh7_w39_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid653_Out0_c1(0);
   bh7_w40_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid653_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid653: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid653_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid653_Out0_copy654_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid653_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid653_Out0_copy654_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid655_In0_c1 <= "" & bh7_w40_0_c1 & bh7_w40_1_c1 & bh7_w40_2_c1 & bh7_w40_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid655_In1_c1 <= "" & bh7_w41_0_c1;
   bh7_w40_6_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid655_Out0_c1(0);
   bh7_w41_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid655_Out0_c1(1);
   bh7_w42_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid655_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid655: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid655_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid655_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid655_Out0_copy656_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid655_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid655_Out0_copy656_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid657_In0_c1 <= "" & bh7_w41_1_c1 & bh7_w41_2_c1 & bh7_w41_3_c1;
   bh7_w41_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid657_Out0_c1(0);
   bh7_w42_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid657_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid657: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid657_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid657_Out0_copy658_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid657_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid657_Out0_copy658_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid659_In0_c1 <= "" & bh7_w42_0_c1 & bh7_w42_1_c1 & bh7_w42_2_c1 & bh7_w42_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid659_In1_c1 <= "" & bh7_w43_0_c1;
   bh7_w42_6_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid659_Out0_c1(0);
   bh7_w43_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid659_Out0_c1(1);
   bh7_w44_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid659_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid659: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid659_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid659_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid659_Out0_copy660_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid659_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid659_Out0_copy660_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid661_In0_c1 <= "" & bh7_w43_1_c1 & bh7_w43_2_c1 & bh7_w43_3_c1;
   bh7_w43_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid661_Out0_c1(0);
   bh7_w44_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid661_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid661: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid661_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid661_Out0_copy662_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid661_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid661_Out0_copy662_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid663_In0_c1 <= "" & bh7_w44_0_c1 & bh7_w44_1_c1 & bh7_w44_2_c1 & bh7_w44_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid663_In1_c1 <= "" & bh7_w45_0_c1;
   bh7_w44_6_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid663_Out0_c1(0);
   bh7_w45_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid663_Out0_c1(1);
   bh7_w46_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid663_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid663: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid663_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid663_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid663_Out0_copy664_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid663_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid663_Out0_copy664_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid665_In0_c1 <= "" & bh7_w45_1_c1 & bh7_w45_2_c1 & bh7_w45_3_c1;
   bh7_w45_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid665_Out0_c1(0);
   bh7_w46_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid665_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid665: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid665_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid665_Out0_copy666_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid665_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid665_Out0_copy666_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid667_In0_c1 <= "" & bh7_w46_0_c1 & bh7_w46_1_c1 & bh7_w46_2_c1 & bh7_w46_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid667_In1_c1 <= "" & bh7_w47_0_c1;
   bh7_w46_6_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid667_Out0_c1(0);
   bh7_w47_4_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid667_Out0_c1(1);
   bh7_w48_5_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid667_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid667: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid667_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid667_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid667_Out0_copy668_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid667_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid667_Out0_copy668_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid669_In0_c1 <= "" & bh7_w47_1_c1 & bh7_w47_2_c1 & bh7_w47_3_c1;
   bh7_w47_5_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid669_Out0_c1(0);
   bh7_w48_6_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid669_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid669: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid669_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid669_Out0_copy670_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid669_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid669_Out0_copy670_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid671_In0_c1 <= "" & bh7_w48_4_c1 & bh7_w48_0_c1 & bh7_w48_1_c1 & bh7_w48_2_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid671_In1_c0 <= "" & bh7_w49_5_c0;
   bh7_w48_7_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid671_Out0_c1(0);
   bh7_w49_6_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid671_Out0_c1(1);
   bh7_w50_7_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid671_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid671: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid671_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid671_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid671_Out0_copy672_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid671_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid671_Out0_copy672_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid673_In0_c1 <= "" & bh7_w49_0_c1 & bh7_w49_1_c1 & bh7_w49_2_c1 & bh7_w49_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid673_In1_c0 <= "" & bh7_w50_6_c0;
   bh7_w49_7_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid673_Out0_c1(0);
   bh7_w50_8_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid673_Out0_c1(1);
   bh7_w51_11_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid673_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid673: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid673_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid673_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid673_Out0_copy674_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid673_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid673_Out0_copy674_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid675_In0_c1 <= "" & bh7_w50_0_c1 & bh7_w50_1_c1 & bh7_w50_2_c1 & bh7_w50_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid675_In1_c0 <= "" & bh7_w51_10_c0;
   bh7_w50_9_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid675_Out0_c1(0);
   bh7_w51_12_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid675_Out0_c1(1);
   bh7_w52_12_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid675_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid675: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid675_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid675_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid675_Out0_copy676_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid675_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid675_Out0_copy676_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid677_In0_c1 <= "" & bh7_w51_0_c1 & bh7_w51_1_c1 & bh7_w51_3_c1 & bh7_w51_4_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid677_In1_c0 <= "" & bh7_w52_11_c0;
   bh7_w51_13_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid677_Out0_c1(0);
   bh7_w52_13_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid677_Out0_c1(1);
   bh7_w53_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid677_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid677: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid677_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid677_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid677_Out0_copy678_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid677_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid677_Out0_copy678_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid679_In0_c1 <= "" & bh7_w52_0_c1 & bh7_w52_1_c1 & bh7_w52_3_c1 & bh7_w52_4_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid679_In1_c1 <= "" & bh7_w53_14_c1;
   bh7_w52_14_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid679_Out0_c1(0);
   bh7_w53_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid679_Out0_c1(1);
   bh7_w54_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid679_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid679: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid679_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid679_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid679_Out0_copy680_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid679_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid679_Out0_copy680_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid681_In0_c1 <= "" & bh7_w53_0_c1 & bh7_w53_1_c1 & bh7_w53_3_c1 & bh7_w53_4_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid681_In1_c1 <= "" & bh7_w54_15_c1;
   bh7_w53_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid681_Out0_c1(0);
   bh7_w54_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid681_Out0_c1(1);
   bh7_w55_18_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid681_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid681: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid681_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid681_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid681_Out0_copy682_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid681_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid681_Out0_copy682_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid683_In0_c1 <= "" & bh7_w54_0_c1 & bh7_w54_1_c1 & bh7_w54_4_c1 & bh7_w54_5_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid683_In1_c1 <= "" & bh7_w55_17_c1;
   bh7_w54_18_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid683_Out0_c1(0);
   bh7_w55_19_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid683_Out0_c1(1);
   bh7_w56_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid683_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid683: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid683_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid683_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid683_Out0_copy684_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid683_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid683_Out0_copy684_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid685_In0_c1 <= "" & bh7_w55_0_c1 & bh7_w55_1_c1 & bh7_w55_4_c1 & bh7_w55_5_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid685_In1_c1 <= "" & bh7_w56_15_c1;
   bh7_w55_20_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid685_Out0_c1(0);
   bh7_w56_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid685_Out0_c1(1);
   bh7_w57_20_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid685_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid685: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid685_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid685_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid685_Out0_copy686_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid685_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid685_Out0_copy686_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid687_In0_c1 <= "" & bh7_w56_0_c1 & bh7_w56_1_c1 & bh7_w56_3_c1;
   bh7_w56_18_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid687_Out0_c1(0);
   bh7_w57_21_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid687_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid687: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid687_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid687_Out0_copy688_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid687_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid687_Out0_copy688_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid689_In0_c1 <= "" & bh7_w57_18_c1 & bh7_w57_19_c1 & bh7_w57_0_c1 & bh7_w57_1_c1 & bh7_w57_4_c1 & bh7_w57_5_c1;
   bh7_w57_22_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid689_Out0_c1(0);
   bh7_w58_19_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid689_Out0_c1(1);
   bh7_w59_16_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid689_Out0_c1(2);
   Compressor_6_3_Freq500_uid334_uid689: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid689_In0_c1,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid689_Out0_copy690_c1);
   Compressor_6_3_Freq500_uid334_bh7_uid689_Out0_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid689_Out0_copy690_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq500_uid400_bh7_uid691_In0_c1 <= "" & bh7_w58_18_c1 & bh7_w58_0_c1 & bh7_w58_3_c1 & bh7_w58_4_c1 & bh7_w58_5_c1;
   bh7_w58_20_c1 <= Compressor_5_3_Freq500_uid400_bh7_uid691_Out0_c1(0);
   bh7_w59_17_c1 <= Compressor_5_3_Freq500_uid400_bh7_uid691_Out0_c1(1);
   bh7_w60_19_c1 <= Compressor_5_3_Freq500_uid400_bh7_uid691_Out0_c1(2);
   Compressor_5_3_Freq500_uid400_uid691: Compressor_5_3_Freq500_uid400
      port map ( X0 => Compressor_5_3_Freq500_uid400_bh7_uid691_In0_c1,
                 R => Compressor_5_3_Freq500_uid400_bh7_uid691_Out0_copy692_c1);
   Compressor_5_3_Freq500_uid400_bh7_uid691_Out0_c1 <= Compressor_5_3_Freq500_uid400_bh7_uid691_Out0_copy692_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid693_In0_c1 <= "" & bh7_w59_14_c1 & bh7_w59_15_c1 & bh7_w59_0_c1 & bh7_w59_2_c1 & bh7_w59_3_c1 & bh7_w59_4_c1;
   bh7_w59_18_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid693_Out0_c1(0);
   bh7_w60_20_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid693_Out0_c1(1);
   bh7_w61_19_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid693_Out0_c1(2);
   Compressor_6_3_Freq500_uid334_uid693: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid693_In0_c1,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid693_Out0_copy694_c1);
   Compressor_6_3_Freq500_uid334_bh7_uid693_Out0_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid693_Out0_copy694_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid695_In0_c1 <= "" & bh7_w60_18_c1 & bh7_w60_0_c1 & bh7_w60_3_c1 & bh7_w60_4_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid695_In1_c1 <= "" & bh7_w61_18_c1;
   bh7_w60_21_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid695_Out0_c1(0);
   bh7_w61_20_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid695_Out0_c1(1);
   bh7_w62_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid695_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid695: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid695_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid695_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid695_Out0_copy696_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid695_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid695_Out0_copy696_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid697_In0_c1 <= "" & bh7_w61_0_c1 & bh7_w61_3_c1 & bh7_w61_4_c1;
   bh7_w61_21_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid697_Out0_c1(0);
   bh7_w62_17_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid697_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid697: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid697_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid697_Out0_copy698_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid697_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid697_Out0_copy698_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq500_uid334_bh7_uid699_In0_c1 <= "" & bh7_w62_14_c1 & bh7_w62_15_c1 & bh7_w62_0_c1 & bh7_w62_2_c1 & bh7_w62_3_c1 & bh7_w62_4_c1;
   bh7_w62_18_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid699_Out0_c1(0);
   bh7_w63_19_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid699_Out0_c1(1);
   bh7_w64_19_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid699_Out0_c1(2);
   Compressor_6_3_Freq500_uid334_uid699: Compressor_6_3_Freq500_uid334
      port map ( X0 => Compressor_6_3_Freq500_uid334_bh7_uid699_In0_c1,
                 R => Compressor_6_3_Freq500_uid334_bh7_uid699_Out0_copy700_c1);
   Compressor_6_3_Freq500_uid334_bh7_uid699_Out0_c1 <= Compressor_6_3_Freq500_uid334_bh7_uid699_Out0_copy700_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid701_In0_c1 <= "" & bh7_w63_18_c1 & bh7_w63_0_c1 & bh7_w63_3_c1 & bh7_w63_4_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid701_In1_c1 <= "" & bh7_w64_18_c1;
   bh7_w63_20_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid701_Out0_c1(0);
   bh7_w64_20_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid701_Out0_c1(1);
   bh7_w65_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid701_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid701: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid701_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid701_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid701_Out0_copy702_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid701_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid701_Out0_copy702_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid703_In0_c1 <= "" & bh7_w64_0_c1 & bh7_w64_3_c1 & bh7_w64_4_c1 & bh7_w64_5_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid703_In1_c1 <= "" & bh7_w65_13_c1;
   bh7_w64_21_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid703_Out0_c1(0);
   bh7_w65_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid703_Out0_c1(1);
   bh7_w66_18_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid703_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid703: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid703_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid703_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid703_Out0_copy704_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid703_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid703_Out0_copy704_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid705_In0_c1 <= "" & bh7_w65_14_c1 & bh7_w65_0_c1 & bh7_w65_2_c1 & bh7_w65_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid705_In1_c1 <= "" & bh7_w66_17_c1;
   bh7_w65_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid705_Out0_c1(0);
   bh7_w66_19_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid705_Out0_c1(1);
   bh7_w67_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid705_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid705: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid705_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid705_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid705_Out0_copy706_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid705_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid705_Out0_copy706_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid707_In0_c1 <= "" & bh7_w66_0_c1 & bh7_w66_3_c1 & bh7_w66_4_c1;
   bh7_w66_20_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid707_Out0_c1(0);
   bh7_w67_17_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid707_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid707: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid707_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid707_Out0_copy708_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid707_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid707_Out0_copy708_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid709_In0_c1 <= "" & bh7_w67_15_c1 & bh7_w67_0_c1 & bh7_w67_3_c1 & bh7_w67_4_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid709_In1_c1 <= "" & bh7_w68_17_c1;
   bh7_w67_18_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid709_Out0_c1(0);
   bh7_w68_19_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid709_Out0_c1(1);
   bh7_w69_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid709_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid709: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid709_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid709_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid709_Out0_copy710_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid709_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid709_Out0_copy710_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid711_In0_c1 <= "" & bh7_w68_18_c1 & bh7_w68_0_c1 & bh7_w68_2_c1 & bh7_w68_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid711_In1_c1 <= "" & bh7_w69_14_c1;
   bh7_w68_20_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid711_Out0_c1(0);
   bh7_w69_16_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid711_Out0_c1(1);
   bh7_w70_18_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid711_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid711: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid711_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid711_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid711_Out0_copy712_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid711_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid711_Out0_copy712_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid713_In0_c1 <= "" & bh7_w69_0_c1 & bh7_w69_3_c1 & bh7_w69_4_c1;
   bh7_w69_17_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid713_Out0_c1(0);
   bh7_w70_19_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid713_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid713: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid713_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid713_Out0_copy714_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid713_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid713_Out0_copy714_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid715_In0_c1 <= "" & bh7_w70_16_c1 & bh7_w70_17_c1 & bh7_w70_0_c1 & bh7_w70_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid715_In1_c1 <= "" & bh7_w71_14_c1;
   bh7_w70_20_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid715_Out0_c1(0);
   bh7_w71_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid715_Out0_c1(1);
   bh7_w72_18_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid715_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid715: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid715_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid715_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid715_Out0_copy716_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid715_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid715_Out0_copy716_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid717_In0_c1 <= "" & bh7_w71_0_c1 & bh7_w71_2_c1 & bh7_w71_3_c1;
   bh7_w71_16_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid717_Out0_c1(0);
   bh7_w72_19_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid717_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid717: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid717_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid717_Out0_copy718_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid717_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid717_Out0_copy718_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid719_In0_c1 <= "" & bh7_w72_16_c1 & bh7_w72_17_c1 & bh7_w72_0_c1 & bh7_w72_3_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid719_In1_c1 <= "" & bh7_w73_14_c1;
   bh7_w72_20_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid719_Out0_c1(0);
   bh7_w73_15_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid719_Out0_c1(1);
   bh7_w74_18_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid719_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid719: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid719_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid719_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid719_Out0_copy720_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid719_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid719_Out0_copy720_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid721_In0_c1 <= "" & bh7_w73_0_c1 & bh7_w73_3_c1 & bh7_w73_4_c1;
   bh7_w73_16_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid721_Out0_c1(0);
   bh7_w74_19_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid721_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid721: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid721_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid721_Out0_copy722_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid721_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid721_Out0_copy722_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid723_In0_c1 <= "" & bh7_w74_17_c1 & bh7_w74_16_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid723_In1_c1 <= "" & bh7_w75_13_c1;
   bh7_w74_20_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid723_Out0_c1(0);
   bh7_w75_14_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid723_Out0_c1(1);
   bh7_w76_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid723_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid723: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid723_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid723_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid723_Out0_copy724_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid723_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid723_Out0_copy724_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid725_In0_c1 <= "" & bh7_w74_0_c1 & bh7_w74_2_c1 & bh7_w74_3_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid725_In1_c1 <= "" & bh7_w75_1_c1 & bh7_w75_2_c1;
   bh7_w74_21_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid725_Out0_c1(0);
   bh7_w75_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid725_Out0_c1(1);
   bh7_w76_18_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid725_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid725: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid725_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid725_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid725_Out0_copy726_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid725_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid725_Out0_copy726_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid727_In0_c1 <= "" & bh7_w76_16_c1 & bh7_w76_15_c1 & bh7_w76_1_c1 & bh7_w76_2_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid727_In1_c0 <= "" & "0";
   bh7_w76_19_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid727_Out0_c1(0);
   bh7_w77_14_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid727_Out0_c1(1);
   bh7_w78_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid727_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid727: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid727_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid727_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid727_Out0_copy728_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid727_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid727_Out0_copy728_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid729_In0_c1 <= "" & bh7_w77_13_c1 & bh7_w77_0_c1 & bh7_w77_1_c1;
   bh7_w77_15_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid729_Out0_c1(0);
   bh7_w78_18_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid729_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid729: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid729_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid729_Out0_copy730_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid729_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid729_Out0_copy730_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid731_In0_c1 <= "" & bh7_w78_16_c1 & bh7_w78_15_c1 & bh7_w78_0_c1 & bh7_w78_1_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid731_In1_c0 <= "" & "0";
   bh7_w78_19_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid731_Out0_c1(0);
   bh7_w79_14_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid731_Out0_c1(1);
   bh7_w80_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid731_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid731: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid731_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid731_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid731_Out0_copy732_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid731_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid731_Out0_copy732_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid733_In0_c1 <= "" & bh7_w79_13_c1 & bh7_w79_0_c1 & bh7_w79_1_c1;
   bh7_w79_15_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid733_Out0_c1(0);
   bh7_w80_18_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid733_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid733: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid733_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid733_Out0_copy734_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid733_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid733_Out0_copy734_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid735_In0_c1 <= "" & bh7_w80_16_c1 & bh7_w80_15_c1 & bh7_w80_0_c1 & bh7_w80_1_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid735_In1_c0 <= "" & "0";
   bh7_w80_19_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid735_Out0_c1(0);
   bh7_w81_14_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid735_Out0_c1(1);
   bh7_w82_17_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid735_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid735: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid735_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid735_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid735_Out0_copy736_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid735_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid735_Out0_copy736_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid737_In0_c1 <= "" & bh7_w81_13_c1 & bh7_w81_0_c1 & bh7_w81_1_c1;
   bh7_w81_15_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid737_Out0_c1(0);
   bh7_w82_18_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid737_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid737: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid737_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid737_Out0_copy738_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid737_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid737_Out0_copy738_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid739_In0_c1 <= "" & bh7_w82_16_c1 & bh7_w82_15_c1 & bh7_w82_0_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid739_In1_c1 <= "" & bh7_w83_13_c1 & bh7_w83_0_c1;
   bh7_w82_19_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid739_Out0_c1(0);
   bh7_w83_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid739_Out0_c1(1);
   bh7_w84_17_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid739_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid739: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid739_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid739_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid739_Out0_copy740_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid739_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid739_Out0_copy740_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid741_In0_c1 <= "" & bh7_w84_15_c1 & bh7_w84_16_c1 & bh7_w84_0_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid741_In1_c1 <= "" & bh7_w85_14_c1 & bh7_w85_0_c1;
   bh7_w84_18_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid741_Out0_c1(0);
   bh7_w85_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid741_Out0_c1(1);
   bh7_w86_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid741_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid741: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid741_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid741_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid741_Out0_copy742_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid741_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid741_Out0_copy742_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid743_In0_c1 <= "" & bh7_w86_13_c1 & bh7_w86_14_c1 & bh7_w86_0_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid743_In1_c1 <= "" & bh7_w87_15_c1 & bh7_w87_0_c1;
   bh7_w86_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid743_Out0_c1(0);
   bh7_w87_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid743_Out0_c1(1);
   bh7_w88_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid743_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid743: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid743_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid743_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid743_Out0_copy744_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid743_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid743_Out0_copy744_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid745_In0_c1 <= "" & bh7_w88_13_c1 & bh7_w88_14_c1 & bh7_w88_0_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid745_In1_c1 <= "" & bh7_w89_13_c1 & bh7_w89_0_c1;
   bh7_w88_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid745_Out0_c1(0);
   bh7_w89_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid745_Out0_c1(1);
   bh7_w90_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid745_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid745: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid745_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid745_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid745_Out0_copy746_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid745_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid745_Out0_copy746_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid747_In0_c1 <= "" & bh7_w90_15_c1 & bh7_w90_0_c1 & "0";
   bh7_w90_17_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid747_Out0_c1(0);
   bh7_w91_15_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid747_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid747: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid747_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid747_Out0_copy748_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid747_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid747_Out0_copy748_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid749_In0_c1 <= "" & bh7_w91_13_c1 & bh7_w91_14_c1 & bh7_w91_0_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid749_In1_c1 <= "" & bh7_w92_13_c1 & bh7_w92_0_c1;
   bh7_w91_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid749_Out0_c1(0);
   bh7_w92_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid749_Out0_c1(1);
   bh7_w93_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid749_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid749: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid749_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid749_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid749_Out0_copy750_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid749_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid749_Out0_copy750_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid751_In0_c1 <= "" & bh7_w93_15_c1 & bh7_w93_0_c1 & "0";
   bh7_w93_17_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid751_Out0_c1(0);
   bh7_w94_15_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid751_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid751: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid751_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid751_Out0_copy752_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid751_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid751_Out0_copy752_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid753_In0_c1 <= "" & bh7_w94_13_c1 & bh7_w94_14_c1 & bh7_w94_0_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid753_In1_c1 <= "" & bh7_w95_13_c1 & bh7_w95_0_c1;
   bh7_w94_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid753_Out0_c1(0);
   bh7_w95_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid753_Out0_c1(1);
   bh7_w96_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid753_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid753: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid753_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid753_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid753_Out0_copy754_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid753_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid753_Out0_copy754_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid755_In0_c1 <= "" & bh7_w96_15_c1 & bh7_w96_0_c1 & "0";
   bh7_w96_17_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid755_Out0_c1(0);
   bh7_w97_15_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid755_Out0_c1(1);
   Compressor_3_2_Freq500_uid432_uid755: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid755_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid755_Out0_copy756_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid755_Out0_c1 <= Compressor_3_2_Freq500_uid432_bh7_uid755_Out0_copy756_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid757_In0_c1 <= "" & bh7_w97_13_c1 & bh7_w97_14_c1 & bh7_w97_0_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid757_In1_c1 <= "" & bh7_w98_13_c1 & bh7_w98_0_c1;
   bh7_w97_16_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid757_Out0_c1(0);
   bh7_w98_14_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid757_Out0_c1(1);
   bh7_w99_15_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid757_Out0_c1(2);
   Compressor_23_3_Freq500_uid322_uid757: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid757_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid757_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid757_Out0_copy758_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid757_Out0_c1 <= Compressor_23_3_Freq500_uid322_bh7_uid757_Out0_copy758_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid759_In0_c1 <= "" & bh7_w100_10_c1 & bh7_w100_11_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid759_In1_c1 <= "" & bh7_w101_10_c1;
   bh7_w100_12_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid759_Out0_c1(0);
   bh7_w101_11_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid759_Out0_c1(1);
   bh7_w102_10_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid759_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid759: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid759_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid759_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid759_Out0_copy760_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid759_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid759_Out0_copy760_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid761_In0_c1 <= "" & bh7_w103_7_c1 & bh7_w103_8_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid761_In1_c1 <= "" & bh7_w104_4_c1;
   bh7_w103_9_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid761_Out0_c1(0);
   bh7_w104_5_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid761_Out0_c1(1);
   bh7_w105_6_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid761_Out0_c1(2);
   Compressor_14_3_Freq500_uid326_uid761: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid761_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid761_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid761_Out0_copy762_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid761_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid761_Out0_copy762_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid763_In0_c1 <= "" & bh7_w105_5_c1 & bh7_w105_4_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid763_In1_c0 <= "" & "0";
   bh7_w105_7_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid763_Out0_c1(0);
   Compressor_14_3_Freq500_uid326_uid763: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid763_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid763_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid763_Out0_copy764_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid763_Out0_c1 <= Compressor_14_3_Freq500_uid326_bh7_uid763_Out0_copy764_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid765_In0_c1 <= "" & bh7_w19_3_c1 & bh7_w19_2_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid765_In1_c1 <= "" & bh7_w20_2_c1;
   bh7_w19_4_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_c2(0);
   bh7_w20_3_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_c2(1);
   bh7_w21_4_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid765: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid765_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid765_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_copy766_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid765_Out0_copy766_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid767_In0_c1 <= "" & bh7_w21_3_c1 & bh7_w21_2_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid767_In1_c1 <= "" & bh7_w22_2_c1;
   bh7_w21_5_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_c2(0);
   bh7_w22_3_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_c2(1);
   bh7_w23_4_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid767: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid767_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid767_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_copy768_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid767_Out0_copy768_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid769_In0_c1 <= "" & bh7_w23_3_c1 & bh7_w23_2_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid769_In1_c1 <= "" & bh7_w24_4_c1 & bh7_w24_3_c1;
   bh7_w23_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_c2(0);
   bh7_w24_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_c2(1);
   bh7_w25_4_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid769: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid769_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid769_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_copy770_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid769_Out0_copy770_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid771_In0_c1 <= "" & bh7_w25_2_c1 & bh7_w25_3_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid771_In1_c1 <= "" & bh7_w26_4_c1 & bh7_w26_3_c1;
   bh7_w25_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_c2(0);
   bh7_w26_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_c2(1);
   bh7_w27_4_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid771: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid771_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid771_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_copy772_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid771_Out0_copy772_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid773_In0_c1 <= "" & bh7_w27_2_c1 & bh7_w27_3_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid773_In1_c1 <= "" & bh7_w28_4_c1 & bh7_w28_3_c1;
   bh7_w27_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_c2(0);
   bh7_w28_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_c2(1);
   bh7_w29_4_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid773: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid773_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid773_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_copy774_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid773_Out0_copy774_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid775_In0_c1 <= "" & bh7_w29_2_c1 & bh7_w29_3_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid775_In1_c1 <= "" & bh7_w30_4_c1 & bh7_w30_3_c1;
   bh7_w29_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_c2(0);
   bh7_w30_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_c2(1);
   bh7_w31_4_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid775: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid775_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid775_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_copy776_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid775_Out0_copy776_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid777_In0_c1 <= "" & bh7_w31_2_c1 & bh7_w31_3_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid777_In1_c1 <= "" & bh7_w32_4_c1 & bh7_w32_3_c1;
   bh7_w31_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_c2(0);
   bh7_w32_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_c2(1);
   bh7_w33_4_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid777: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid777_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid777_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_copy778_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid777_Out0_copy778_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid779_In0_c1 <= "" & bh7_w33_2_c1 & bh7_w33_3_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid779_In1_c1 <= "" & bh7_w34_5_c1 & bh7_w34_4_c1;
   bh7_w33_5_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_c2(0);
   bh7_w34_6_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_c2(1);
   bh7_w35_6_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid779: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid779_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid779_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_copy780_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid779_Out0_copy780_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid781_In0_c1 <= "" & bh7_w35_5_c1 & bh7_w35_4_c1 & "0";
   bh7_w35_7_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_c2(0);
   bh7_w36_7_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_c2(1);
   Compressor_3_2_Freq500_uid432_uid781: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid781_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_copy782_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid781_Out0_copy782_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid783_In0_c1 <= "" & bh7_w36_6_c1 & bh7_w36_5_c1 & bh7_w36_4_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid783_In1_c1 <= "" & bh7_w37_5_c1 & bh7_w37_4_c1;
   bh7_w36_8_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_c2(0);
   bh7_w37_6_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_c2(1);
   bh7_w38_7_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid783: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid783_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid783_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_copy784_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid783_Out0_copy784_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid785_In0_c1 <= "" & bh7_w38_6_c1 & bh7_w38_5_c1 & bh7_w38_4_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid785_In1_c1 <= "" & bh7_w39_5_c1 & bh7_w39_4_c1;
   bh7_w38_8_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_c2(0);
   bh7_w39_6_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_c2(1);
   bh7_w40_7_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid785: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid785_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid785_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_copy786_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid785_Out0_copy786_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid787_In0_c1 <= "" & bh7_w40_6_c1 & bh7_w40_5_c1 & bh7_w40_4_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid787_In1_c1 <= "" & bh7_w41_5_c1 & bh7_w41_4_c1;
   bh7_w40_8_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_c2(0);
   bh7_w41_6_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_c2(1);
   bh7_w42_7_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid787: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid787_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid787_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_copy788_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid787_Out0_copy788_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid789_In0_c1 <= "" & bh7_w42_6_c1 & bh7_w42_5_c1 & bh7_w42_4_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid789_In1_c1 <= "" & bh7_w43_5_c1 & bh7_w43_4_c1;
   bh7_w42_8_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_c2(0);
   bh7_w43_6_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_c2(1);
   bh7_w44_7_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid789: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid789_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid789_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_copy790_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid789_Out0_copy790_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid791_In0_c1 <= "" & bh7_w44_6_c1 & bh7_w44_5_c1 & bh7_w44_4_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid791_In1_c1 <= "" & bh7_w45_5_c1 & bh7_w45_4_c1;
   bh7_w44_8_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_c2(0);
   bh7_w45_6_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_c2(1);
   bh7_w46_7_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid791: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid791_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid791_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_copy792_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid791_Out0_copy792_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid793_In0_c1 <= "" & bh7_w46_6_c1 & bh7_w46_5_c1 & bh7_w46_4_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid793_In1_c1 <= "" & bh7_w47_5_c1 & bh7_w47_4_c1;
   bh7_w46_8_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_c2(0);
   bh7_w47_6_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_c2(1);
   bh7_w48_8_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid793: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid793_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid793_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_copy794_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid793_Out0_copy794_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid795_In0_c1 <= "" & bh7_w48_3_c1 & bh7_w48_7_c1 & bh7_w48_6_c1 & bh7_w48_5_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid795_In1_c1 <= "" & bh7_w49_7_c1;
   bh7_w48_9_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_c2(0);
   bh7_w49_8_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_c2(1);
   bh7_w50_10_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid795: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid795_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid795_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_copy796_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid795_Out0_copy796_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid797_In0_c1 <= "" & bh7_w50_9_c1 & bh7_w50_8_c1 & bh7_w50_7_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid797_In1_c1 <= "" & bh7_w51_13_c1 & bh7_w51_12_c1;
   bh7_w50_11_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_c2(0);
   bh7_w51_14_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_c2(1);
   bh7_w52_15_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid797: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid797_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid797_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_copy798_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid797_Out0_copy798_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid799_In0_c1 <= "" & bh7_w52_14_c1 & bh7_w52_13_c1 & bh7_w52_12_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid799_In1_c1 <= "" & bh7_w53_17_c1 & bh7_w53_16_c1;
   bh7_w52_16_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_c2(0);
   bh7_w53_18_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_c2(1);
   bh7_w54_19_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid799: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid799_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid799_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_copy800_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid799_Out0_copy800_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid801_In0_c1 <= "" & bh7_w54_18_c1 & bh7_w54_17_c1 & bh7_w54_16_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid801_In1_c1 <= "" & bh7_w55_19_c1 & bh7_w55_20_c1;
   bh7_w54_20_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_c2(0);
   bh7_w55_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_c2(1);
   bh7_w56_19_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid801: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid801_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid801_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_copy802_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid801_Out0_copy802_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid803_In0_c1 <= "" & bh7_w56_16_c1 & bh7_w56_17_c1 & bh7_w56_4_c1 & bh7_w56_18_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid803_In1_c0 <= "" & "0";
   bh7_w56_20_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_c2(0);
   bh7_w57_23_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_c2(1);
   bh7_w58_21_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid803: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid803_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid803_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_copy804_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid803_Out0_copy804_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid805_In0_c1 <= "" & bh7_w57_20_c1 & bh7_w57_22_c1 & bh7_w57_21_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid805_In1_c1 <= "" & bh7_w58_19_c1 & bh7_w58_20_c1;
   bh7_w57_24_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_c2(0);
   bh7_w58_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_c2(1);
   bh7_w59_19_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid805: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid805_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid805_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_copy806_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid805_Out0_copy806_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid807_In0_c1 <= "" & bh7_w59_16_c1 & bh7_w59_17_c1 & bh7_w59_18_c1;
   bh7_w59_20_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_c2(0);
   bh7_w60_22_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_c2(1);
   Compressor_3_2_Freq500_uid432_uid807: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid807_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_copy808_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid807_Out0_copy808_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid809_In0_c1 <= "" & bh7_w60_19_c1 & bh7_w60_20_c1 & bh7_w60_21_c1 & bh7_w60_5_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid809_In1_c1 <= "" & bh7_w61_19_c1;
   bh7_w60_23_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_c2(0);
   bh7_w61_22_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_c2(1);
   bh7_w62_19_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid809: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid809_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid809_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_copy810_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid809_Out0_copy810_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid811_In0_c1 <= "" & bh7_w61_20_c1 & bh7_w61_5_c1 & bh7_w61_21_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid811_In1_c1 <= "" & bh7_w62_16_c1 & bh7_w62_18_c1;
   bh7_w61_23_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_c2(0);
   bh7_w62_20_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_c2(1);
   bh7_w63_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid811: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid811_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid811_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_copy812_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid811_Out0_copy812_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid813_In0_c1 <= "" & bh7_w63_19_c1 & bh7_w63_20_c1 & bh7_w63_5_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid813_In1_c1 <= "" & bh7_w64_19_c1 & bh7_w64_20_c1;
   bh7_w63_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_c2(0);
   bh7_w64_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_c2(1);
   bh7_w65_18_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid813: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid813_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid813_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_copy814_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid813_Out0_copy814_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid815_In0_c1 <= "" & bh7_w65_15_c1 & bh7_w65_16_c1 & bh7_w65_17_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid815_In1_c1 <= "" & bh7_w66_18_c1 & bh7_w66_19_c1;
   bh7_w65_19_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_c2(0);
   bh7_w66_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_c2(1);
   bh7_w67_19_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid815: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid815_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid815_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_copy816_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid815_Out0_copy816_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid817_In0_c1 <= "" & bh7_w67_16_c1 & bh7_w67_18_c1 & bh7_w67_17_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid817_In1_c1 <= "" & bh7_w68_19_c1 & bh7_w68_20_c1;
   bh7_w67_20_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_c2(0);
   bh7_w68_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_c2(1);
   bh7_w69_18_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid817: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid817_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid817_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_copy818_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid817_Out0_copy818_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid819_In0_c1 <= "" & bh7_w69_15_c1 & bh7_w69_16_c1 & bh7_w69_17_c1;
   bh7_w69_19_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_c2(0);
   bh7_w70_21_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_c2(1);
   Compressor_3_2_Freq500_uid432_uid819: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid819_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_copy820_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid819_Out0_copy820_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid821_In0_c1 <= "" & bh7_w70_18_c1 & bh7_w70_20_c1 & bh7_w70_4_c1 & bh7_w70_19_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid821_In1_c1 <= "" & bh7_w71_15_c1;
   bh7_w70_22_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_c2(0);
   bh7_w71_17_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_c2(1);
   bh7_w72_21_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid821: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid821_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid821_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_copy822_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid821_Out0_copy822_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid823_In0_c1 <= "" & bh7_w72_18_c1 & bh7_w72_20_c1 & bh7_w72_4_c1 & bh7_w72_19_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid823_In1_c1 <= "" & bh7_w73_15_c1;
   bh7_w72_22_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_c2(0);
   bh7_w73_17_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_c2(1);
   bh7_w74_22_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid823: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid823_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid823_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_copy824_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid823_Out0_copy824_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid825_In0_c1 <= "" & bh7_w74_18_c1 & bh7_w74_20_c1 & bh7_w74_21_c1 & bh7_w74_19_c1;
   Compressor_14_3_Freq500_uid326_bh7_uid825_In1_c1 <= "" & bh7_w75_14_c1;
   bh7_w74_23_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_c2(0);
   bh7_w75_16_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_c2(1);
   bh7_w76_20_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid825: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid825_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid825_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_copy826_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid825_Out0_copy826_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid827_In0_c1 <= "" & bh7_w76_19_c1 & bh7_w76_17_c1 & bh7_w76_18_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid827_In1_c1 <= "" & bh7_w77_14_c1 & bh7_w77_15_c1;
   bh7_w76_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_c2(0);
   bh7_w77_16_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_c2(1);
   bh7_w78_20_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid827: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid827_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid827_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_copy828_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid827_Out0_copy828_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid829_In0_c1 <= "" & bh7_w78_17_c1 & bh7_w78_19_c1 & bh7_w78_18_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid829_In1_c1 <= "" & bh7_w79_14_c1 & bh7_w79_15_c1;
   bh7_w78_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_c2(0);
   bh7_w79_16_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_c2(1);
   bh7_w80_20_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid829: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid829_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid829_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_copy830_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid829_Out0_copy830_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid831_In0_c1 <= "" & bh7_w80_17_c1 & bh7_w80_19_c1 & bh7_w80_18_c1;
   Compressor_23_3_Freq500_uid322_bh7_uid831_In1_c1 <= "" & bh7_w81_14_c1 & bh7_w81_15_c1;
   bh7_w80_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_c2(0);
   bh7_w81_16_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_c2(1);
   bh7_w82_20_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid831: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid831_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid831_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_copy832_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid831_Out0_copy832_c2; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq500_uid432_bh7_uid833_In0_c1 <= "" & bh7_w82_17_c1 & bh7_w82_19_c1 & bh7_w82_18_c1;
   bh7_w82_21_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_c2(0);
   bh7_w83_15_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_c2(1);
   Compressor_3_2_Freq500_uid432_uid833: Compressor_3_2_Freq500_uid432
      port map ( X0 => Compressor_3_2_Freq500_uid432_bh7_uid833_In0_c1,
                 R => Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_copy834_c1);
   Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_c2 <= Compressor_3_2_Freq500_uid432_bh7_uid833_Out0_copy834_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid835_In0_c1 <= "" & bh7_w84_17_c1 & bh7_w84_18_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid835_In1_c1 <= "" & bh7_w85_15_c1;
   bh7_w84_19_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_c2(0);
   bh7_w85_16_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_c2(1);
   bh7_w86_17_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid835: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid835_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid835_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_copy836_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid835_Out0_copy836_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid837_In0_c1 <= "" & bh7_w86_15_c1 & bh7_w86_16_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid837_In1_c1 <= "" & bh7_w87_16_c1;
   bh7_w86_18_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_c2(0);
   bh7_w87_17_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_c2(1);
   bh7_w88_17_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid837: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid837_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid837_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_copy838_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid837_Out0_copy838_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid839_In0_c1 <= "" & bh7_w88_15_c1 & bh7_w88_16_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid839_In1_c1 <= "" & bh7_w89_14_c1;
   bh7_w88_18_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_c2(0);
   bh7_w89_15_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_c2(1);
   bh7_w90_18_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid839: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid839_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid839_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_copy840_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid839_Out0_copy840_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid841_In0_c1 <= "" & bh7_w90_16_c1 & bh7_w90_17_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid841_In1_c1 <= "" & bh7_w91_15_c1 & bh7_w91_16_c1;
   bh7_w90_19_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_c2(0);
   bh7_w91_17_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_c2(1);
   bh7_w92_15_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid841: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid841_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid841_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_copy842_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid841_Out0_copy842_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid843_In0_c1 <= "" & bh7_w93_16_c1 & bh7_w93_17_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid843_In1_c1 <= "" & bh7_w94_15_c1 & bh7_w94_16_c1;
   bh7_w93_18_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_c2(0);
   bh7_w94_17_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_c2(1);
   bh7_w95_15_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid843: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid843_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid843_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_copy844_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid843_Out0_copy844_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid845_In0_c1 <= "" & bh7_w96_16_c1 & bh7_w96_17_c1 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid845_In1_c1 <= "" & bh7_w97_15_c1 & bh7_w97_16_c1;
   bh7_w96_18_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_c2(0);
   bh7_w97_17_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_c2(1);
   bh7_w98_15_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid845: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid845_In0_c1,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid845_In1_c1,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_copy846_c1);
   Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid845_Out0_copy846_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid847_In0_c1 <= "" & bh7_w99_14_c1 & bh7_w99_15_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid847_In1_c1 <= "" & bh7_w100_12_c1;
   bh7_w99_16_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_c2(0);
   bh7_w100_13_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_c2(1);
   bh7_w101_12_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid847: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid847_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid847_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_copy848_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid847_Out0_copy848_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid849_In0_c1 <= "" & bh7_w102_9_c1 & bh7_w102_10_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid849_In1_c1 <= "" & bh7_w103_9_c1;
   bh7_w102_11_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_c2(0);
   bh7_w103_10_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_c2(1);
   bh7_w104_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid849: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid849_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid849_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_copy850_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid849_Out0_copy850_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid851_In0_c1 <= "" & bh7_w105_6_c1 & bh7_w105_7_c1 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid851_In1_c0 <= "" & "0";
   bh7_w105_8_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid851_Out0_c2(0);
   Compressor_14_3_Freq500_uid326_uid851: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid851_In0_c1,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid851_In1_c1,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid851_Out0_copy852_c1);
   Compressor_14_3_Freq500_uid326_bh7_uid851_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid851_Out0_copy852_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid853_In0_c2 <= "" & bh7_w21_5_c2 & bh7_w21_4_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid853_In1_c2 <= "" & bh7_w22_3_c2;
   bh7_w21_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid853_Out0_c2(0);
   bh7_w22_4_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid853_Out0_c2(1);
   bh7_w23_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid853_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid853: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid853_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid853_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid853_Out0_copy854_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid853_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid853_Out0_copy854_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid855_In0_c2 <= "" & bh7_w23_5_c2 & bh7_w23_4_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid855_In1_c2 <= "" & bh7_w24_5_c2;
   bh7_w23_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid855_Out0_c2(0);
   bh7_w24_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid855_Out0_c2(1);
   bh7_w25_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid855_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid855: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid855_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid855_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid855_Out0_copy856_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid855_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid855_Out0_copy856_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid857_In0_c2 <= "" & bh7_w25_5_c2 & bh7_w25_4_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid857_In1_c2 <= "" & bh7_w26_5_c2;
   bh7_w25_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid857_Out0_c2(0);
   bh7_w26_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid857_Out0_c2(1);
   bh7_w27_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid857_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid857: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid857_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid857_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid857_Out0_copy858_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid857_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid857_Out0_copy858_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid859_In0_c2 <= "" & bh7_w27_5_c2 & bh7_w27_4_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid859_In1_c2 <= "" & bh7_w28_5_c2;
   bh7_w27_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid859_Out0_c2(0);
   bh7_w28_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid859_Out0_c2(1);
   bh7_w29_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid859_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid859: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid859_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid859_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid859_Out0_copy860_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid859_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid859_Out0_copy860_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid861_In0_c2 <= "" & bh7_w29_5_c2 & bh7_w29_4_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid861_In1_c2 <= "" & bh7_w30_5_c2;
   bh7_w29_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid861_Out0_c2(0);
   bh7_w30_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid861_Out0_c2(1);
   bh7_w31_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid861_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid861: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid861_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid861_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid861_Out0_copy862_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid861_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid861_Out0_copy862_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid863_In0_c2 <= "" & bh7_w31_5_c2 & bh7_w31_4_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid863_In1_c2 <= "" & bh7_w32_5_c2;
   bh7_w31_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid863_Out0_c2(0);
   bh7_w32_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid863_Out0_c2(1);
   bh7_w33_6_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid863_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid863: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid863_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid863_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid863_Out0_copy864_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid863_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid863_Out0_copy864_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid865_In0_c2 <= "" & bh7_w33_5_c2 & bh7_w33_4_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid865_In1_c2 <= "" & bh7_w34_6_c2;
   bh7_w33_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid865_Out0_c2(0);
   bh7_w34_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid865_Out0_c2(1);
   bh7_w35_8_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid865_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid865: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid865_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid865_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid865_Out0_copy866_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid865_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid865_Out0_copy866_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid867_In0_c2 <= "" & bh7_w35_7_c2 & bh7_w35_6_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid867_In1_c2 <= "" & bh7_w36_8_c2 & bh7_w36_7_c2;
   bh7_w35_9_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid867_Out0_c2(0);
   bh7_w36_9_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid867_Out0_c2(1);
   bh7_w37_7_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid867_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid867: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid867_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid867_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid867_Out0_copy868_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid867_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid867_Out0_copy868_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid869_In0_c2 <= "" & bh7_w38_8_c2 & bh7_w38_7_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid869_In1_c2 <= "" & bh7_w39_6_c2;
   bh7_w38_9_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid869_Out0_c2(0);
   bh7_w39_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid869_Out0_c2(1);
   bh7_w40_9_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid869_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid869: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid869_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid869_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid869_Out0_copy870_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid869_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid869_Out0_copy870_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid871_In0_c2 <= "" & bh7_w40_8_c2 & bh7_w40_7_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid871_In1_c2 <= "" & bh7_w41_6_c2;
   bh7_w40_10_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid871_Out0_c2(0);
   bh7_w41_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid871_Out0_c2(1);
   bh7_w42_9_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid871_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid871: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid871_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid871_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid871_Out0_copy872_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid871_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid871_Out0_copy872_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid873_In0_c2 <= "" & bh7_w42_8_c2 & bh7_w42_7_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid873_In1_c2 <= "" & bh7_w43_6_c2;
   bh7_w42_10_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid873_Out0_c2(0);
   bh7_w43_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid873_Out0_c2(1);
   bh7_w44_9_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid873_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid873: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid873_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid873_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid873_Out0_copy874_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid873_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid873_Out0_copy874_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid875_In0_c2 <= "" & bh7_w44_8_c2 & bh7_w44_7_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid875_In1_c2 <= "" & bh7_w45_6_c2;
   bh7_w44_10_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid875_Out0_c2(0);
   bh7_w45_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid875_Out0_c2(1);
   bh7_w46_9_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid875_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid875: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid875_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid875_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid875_Out0_copy876_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid875_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid875_Out0_copy876_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid877_In0_c2 <= "" & bh7_w46_8_c2 & bh7_w46_7_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid877_In1_c2 <= "" & bh7_w47_6_c2;
   bh7_w46_10_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid877_Out0_c2(0);
   bh7_w47_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid877_Out0_c2(1);
   bh7_w48_10_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid877_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid877: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid877_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid877_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid877_Out0_copy878_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid877_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid877_Out0_copy878_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid879_In0_c2 <= "" & bh7_w48_9_c2 & bh7_w48_8_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid879_In1_c2 <= "" & bh7_w49_6_c2 & bh7_w49_8_c2;
   bh7_w48_11_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid879_Out0_c2(0);
   bh7_w49_9_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid879_Out0_c2(1);
   bh7_w50_12_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid879_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid879: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid879_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid879_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid879_Out0_copy880_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid879_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid879_Out0_copy880_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid881_In0_c2 <= "" & bh7_w50_11_c2 & bh7_w50_10_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid881_In1_c2 <= "" & bh7_w51_11_c2 & bh7_w51_14_c2;
   bh7_w50_13_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid881_Out0_c2(0);
   bh7_w51_15_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid881_Out0_c2(1);
   bh7_w52_17_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid881_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid881: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid881_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid881_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid881_Out0_copy882_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid881_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid881_Out0_copy882_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid883_In0_c2 <= "" & bh7_w52_16_c2 & bh7_w52_15_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid883_In1_c2 <= "" & bh7_w53_15_c2 & bh7_w53_18_c2;
   bh7_w52_18_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid883_Out0_c2(0);
   bh7_w53_19_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid883_Out0_c2(1);
   bh7_w54_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid883_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid883: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid883_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid883_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid883_Out0_copy884_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid883_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid883_Out0_copy884_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid885_In0_c2 <= "" & bh7_w54_20_c2 & bh7_w54_19_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid885_In1_c2 <= "" & bh7_w55_21_c2 & bh7_w55_18_c2;
   bh7_w54_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid885_Out0_c2(0);
   bh7_w55_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid885_Out0_c2(1);
   bh7_w56_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid885_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid885: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid885_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid885_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid885_Out0_copy886_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid885_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid885_Out0_copy886_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid887_In0_c2 <= "" & bh7_w56_19_c2 & bh7_w56_20_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid887_In1_c2 <= "" & bh7_w57_23_c2 & bh7_w57_24_c2;
   bh7_w56_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid887_Out0_c2(0);
   bh7_w57_25_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid887_Out0_c2(1);
   bh7_w58_23_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid887_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid887: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid887_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid887_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid887_Out0_copy888_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid887_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid887_Out0_copy888_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid889_In0_c2 <= "" & bh7_w58_21_c2 & bh7_w58_22_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid889_In1_c2 <= "" & bh7_w59_19_c2 & bh7_w59_20_c2;
   bh7_w58_24_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid889_Out0_c2(0);
   bh7_w59_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid889_Out0_c2(1);
   bh7_w60_24_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid889_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid889: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid889_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid889_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid889_Out0_copy890_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid889_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid889_Out0_copy890_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid891_In0_c2 <= "" & bh7_w60_22_c2 & bh7_w60_23_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid891_In1_c2 <= "" & bh7_w61_22_c2 & bh7_w61_23_c2;
   bh7_w60_25_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid891_Out0_c2(0);
   bh7_w61_24_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid891_Out0_c2(1);
   bh7_w62_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid891_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid891: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid891_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid891_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid891_Out0_copy892_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid891_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid891_Out0_copy892_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid893_In0_c2 <= "" & bh7_w62_19_c2 & bh7_w62_20_c2 & bh7_w62_17_c2;
   Compressor_23_3_Freq500_uid322_bh7_uid893_In1_c2 <= "" & bh7_w63_21_c2 & bh7_w63_22_c2;
   bh7_w62_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid893_Out0_c2(0);
   bh7_w63_23_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid893_Out0_c2(1);
   bh7_w64_23_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid893_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid893: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid893_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid893_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid893_Out0_copy894_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid893_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid893_Out0_copy894_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid895_In0_c2 <= "" & bh7_w64_21_c2 & bh7_w64_22_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid895_In1_c2 <= "" & bh7_w65_18_c2 & bh7_w65_19_c2;
   bh7_w64_24_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid895_Out0_c2(0);
   bh7_w65_20_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid895_Out0_c2(1);
   bh7_w66_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid895_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid895: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid895_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid895_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid895_Out0_copy896_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid895_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid895_Out0_copy896_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid897_In0_c2 <= "" & bh7_w66_21_c2 & bh7_w66_20_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid897_In1_c2 <= "" & bh7_w67_19_c2 & bh7_w67_20_c2;
   bh7_w66_23_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid897_Out0_c2(0);
   bh7_w67_21_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid897_Out0_c2(1);
   bh7_w68_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid897_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid897: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid897_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid897_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid897_Out0_copy898_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid897_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid897_Out0_copy898_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid899_In0_c2 <= "" & bh7_w69_18_c2 & bh7_w69_19_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid899_In1_c2 <= "" & bh7_w70_21_c2 & bh7_w70_22_c2;
   bh7_w69_20_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid899_Out0_c2(0);
   bh7_w70_23_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid899_Out0_c2(1);
   bh7_w71_18_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid899_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid899: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid899_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid899_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid899_Out0_copy900_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid899_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid899_Out0_copy900_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid901_In0_c2 <= "" & bh7_w71_17_c2 & bh7_w71_16_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid901_In1_c2 <= "" & bh7_w72_21_c2 & bh7_w72_22_c2;
   bh7_w71_19_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid901_Out0_c2(0);
   bh7_w72_23_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid901_Out0_c2(1);
   bh7_w73_18_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid901_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid901: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid901_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid901_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid901_Out0_copy902_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid901_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid901_Out0_copy902_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid903_In0_c2 <= "" & bh7_w73_17_c2 & bh7_w73_16_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid903_In1_c2 <= "" & bh7_w74_22_c2 & bh7_w74_23_c2;
   bh7_w73_19_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid903_Out0_c2(0);
   bh7_w74_24_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid903_Out0_c2(1);
   bh7_w75_17_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid903_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid903: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid903_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid903_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid903_Out0_copy904_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid903_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid903_Out0_copy904_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid905_In0_c2 <= "" & bh7_w75_16_c2 & bh7_w75_15_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid905_In1_c2 <= "" & bh7_w76_20_c2 & bh7_w76_21_c2;
   bh7_w75_18_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid905_Out0_c2(0);
   bh7_w76_22_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid905_Out0_c2(1);
   bh7_w77_17_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid905_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid905: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid905_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid905_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid905_Out0_copy906_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid905_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid905_Out0_copy906_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid907_In0_c2 <= "" & bh7_w78_20_c2 & bh7_w78_21_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid907_In1_c2 <= "" & bh7_w79_16_c2;
   bh7_w78_22_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid907_Out0_c2(0);
   bh7_w79_17_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid907_Out0_c2(1);
   bh7_w80_22_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid907_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid907: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid907_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid907_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid907_Out0_copy908_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid907_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid907_Out0_copy908_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid909_In0_c2 <= "" & bh7_w80_20_c2 & bh7_w80_21_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid909_In1_c2 <= "" & bh7_w81_16_c2;
   bh7_w80_23_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid909_Out0_c2(0);
   bh7_w81_17_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid909_Out0_c2(1);
   bh7_w82_22_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid909_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid909: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid909_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid909_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid909_Out0_copy910_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid909_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid909_Out0_copy910_c2; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq500_uid322_bh7_uid911_In0_c2 <= "" & bh7_w82_20_c2 & bh7_w82_21_c2 & "0";
   Compressor_23_3_Freq500_uid322_bh7_uid911_In1_c2 <= "" & bh7_w83_14_c2 & bh7_w83_15_c2;
   bh7_w82_23_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid911_Out0_c2(0);
   bh7_w83_16_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid911_Out0_c2(1);
   bh7_w84_20_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid911_Out0_c2(2);
   Compressor_23_3_Freq500_uid322_uid911: Compressor_23_3_Freq500_uid322
      port map ( X0 => Compressor_23_3_Freq500_uid322_bh7_uid911_In0_c2,
                 X1 => Compressor_23_3_Freq500_uid322_bh7_uid911_In1_c2,
                 R => Compressor_23_3_Freq500_uid322_bh7_uid911_Out0_copy912_c2);
   Compressor_23_3_Freq500_uid322_bh7_uid911_Out0_c2 <= Compressor_23_3_Freq500_uid322_bh7_uid911_Out0_copy912_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid913_In0_c2 <= "" & bh7_w86_17_c2 & bh7_w86_18_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid913_In1_c2 <= "" & bh7_w87_17_c2;
   bh7_w86_19_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid913_Out0_c2(0);
   bh7_w87_18_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid913_Out0_c2(1);
   bh7_w88_19_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid913_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid913: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid913_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid913_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid913_Out0_copy914_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid913_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid913_Out0_copy914_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid915_In0_c2 <= "" & bh7_w88_17_c2 & bh7_w88_18_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid915_In1_c2 <= "" & bh7_w89_15_c2;
   bh7_w88_20_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid915_Out0_c2(0);
   bh7_w89_16_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid915_Out0_c2(1);
   bh7_w90_20_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid915_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid915: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid915_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid915_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid915_Out0_copy916_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid915_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid915_Out0_copy916_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid917_In0_c2 <= "" & bh7_w90_18_c2 & bh7_w90_19_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid917_In1_c2 <= "" & bh7_w91_17_c2;
   bh7_w90_21_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid917_Out0_c2(0);
   bh7_w91_18_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid917_Out0_c2(1);
   bh7_w92_16_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid917_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid917: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid917_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid917_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid917_Out0_copy918_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid917_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid917_Out0_copy918_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid919_In0_c2 <= "" & bh7_w92_14_c2 & bh7_w92_15_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid919_In1_c2 <= "" & bh7_w93_18_c2;
   bh7_w92_17_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid919_Out0_c2(0);
   bh7_w93_19_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid919_Out0_c2(1);
   bh7_w94_18_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid919_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid919: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid919_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid919_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid919_Out0_copy920_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid919_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid919_Out0_copy920_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid921_In0_c2 <= "" & bh7_w95_14_c2 & bh7_w95_15_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid921_In1_c2 <= "" & bh7_w96_18_c2;
   bh7_w95_16_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid921_Out0_c2(0);
   bh7_w96_19_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid921_Out0_c2(1);
   bh7_w97_18_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid921_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid921: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid921_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid921_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid921_Out0_copy922_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid921_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid921_Out0_copy922_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid923_In0_c2 <= "" & bh7_w98_14_c2 & bh7_w98_15_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid923_In1_c2 <= "" & bh7_w99_16_c2;
   bh7_w98_16_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid923_Out0_c2(0);
   bh7_w99_17_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid923_Out0_c2(1);
   bh7_w100_14_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid923_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid923: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid923_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid923_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid923_Out0_copy924_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid923_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid923_Out0_copy924_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid925_In0_c2 <= "" & bh7_w101_11_c2 & bh7_w101_12_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid925_In1_c2 <= "" & bh7_w102_11_c2;
   bh7_w101_13_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid925_Out0_c2(0);
   bh7_w102_12_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid925_Out0_c2(1);
   bh7_w103_11_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid925_Out0_c2(2);
   Compressor_14_3_Freq500_uid326_uid925: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid925_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid925_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid925_Out0_copy926_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid925_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid925_Out0_copy926_c2; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq500_uid326_bh7_uid927_In0_c2 <= "" & bh7_w104_5_c2 & bh7_w104_6_c2 & "0" & "0";
   Compressor_14_3_Freq500_uid326_bh7_uid927_In1_c2 <= "" & bh7_w105_8_c2;
   bh7_w104_7_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid927_Out0_c2(0);
   bh7_w105_9_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid927_Out0_c2(1);
   Compressor_14_3_Freq500_uid326_uid927: Compressor_14_3_Freq500_uid326
      port map ( X0 => Compressor_14_3_Freq500_uid326_bh7_uid927_In0_c2,
                 X1 => Compressor_14_3_Freq500_uid326_bh7_uid927_In1_c2,
                 R => Compressor_14_3_Freq500_uid326_bh7_uid927_Out0_copy928_c2);
   Compressor_14_3_Freq500_uid326_bh7_uid927_Out0_c2 <= Compressor_14_3_Freq500_uid326_bh7_uid927_Out0_copy928_c2; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh7_22_c2 <= bh7_w22_4_c2 & bh7_w21_6_c2 & bh7_w20_3_c2 & bh7_w19_4_c2 & bh7_w18_2_c2 & bh7_w17_2_c2 & bh7_w16_0_c2 & bh7_w15_0_c2 & bh7_w14_0_c2 & bh7_w13_0_c2 & bh7_w12_0_c2 & bh7_w11_0_c2 & bh7_w10_0_c2 & bh7_w9_0_c2 & bh7_w8_0_c2 & bh7_w7_0_c2 & bh7_w6_0_c2 & bh7_w5_0_c2 & bh7_w4_0_c2 & bh7_w3_0_c2 & bh7_w2_0_c2 & bh7_w1_0_c2 & bh7_w0_0_c2;

   bitheapFinalAdd_bh7_In0_c2 <= "0" & bh7_w105_9_c2 & bh7_w104_7_c2 & bh7_w103_10_c2 & bh7_w102_12_c2 & bh7_w101_13_c2 & bh7_w100_13_c2 & bh7_w99_17_c2 & bh7_w98_16_c2 & bh7_w97_17_c2 & bh7_w96_19_c2 & bh7_w95_16_c2 & bh7_w94_17_c2 & bh7_w93_19_c2 & bh7_w92_16_c2 & bh7_w91_18_c2 & bh7_w90_20_c2 & bh7_w89_16_c2 & bh7_w88_19_c2 & bh7_w87_18_c2 & bh7_w86_19_c2 & bh7_w85_16_c2 & bh7_w84_19_c2 & bh7_w83_16_c2 & bh7_w82_22_c2 & bh7_w81_17_c2 & bh7_w80_22_c2 & bh7_w79_17_c2 & bh7_w78_22_c2 & bh7_w77_16_c2 & bh7_w76_22_c2 & bh7_w75_17_c2 & bh7_w74_24_c2 & bh7_w73_18_c2 & bh7_w72_23_c2 & bh7_w71_18_c2 & bh7_w70_23_c2 & bh7_w69_20_c2 & bh7_w68_21_c2 & bh7_w67_21_c2 & bh7_w66_22_c2 & bh7_w65_20_c2 & bh7_w64_23_c2 & bh7_w63_23_c2 & bh7_w62_21_c2 & bh7_w61_24_c2 & bh7_w60_24_c2 & bh7_w59_21_c2 & bh7_w58_23_c2 & bh7_w57_25_c2 & bh7_w56_21_c2 & bh7_w55_22_c2 & bh7_w54_22_c2 & bh7_w53_19_c2 & bh7_w52_18_c2 & bh7_w51_15_c2 & bh7_w50_13_c2 & bh7_w49_9_c2 & bh7_w48_11_c2 & bh7_w47_7_c2 & bh7_w46_10_c2 & bh7_w45_7_c2 & bh7_w44_10_c2 & bh7_w43_7_c2 & bh7_w42_10_c2 & bh7_w41_7_c2 & bh7_w40_10_c2 & bh7_w39_7_c2 & bh7_w38_9_c2 & bh7_w37_6_c2 & bh7_w36_9_c2 & bh7_w35_9_c2 & bh7_w34_7_c2 & bh7_w33_7_c2 & bh7_w32_6_c2 & bh7_w31_7_c2 & bh7_w30_6_c2 & bh7_w29_7_c2 & bh7_w28_6_c2 & bh7_w27_7_c2 & bh7_w26_6_c2 & bh7_w25_7_c2 & bh7_w24_6_c2 & bh7_w23_7_c2;
   bitheapFinalAdd_bh7_In1_c2 <= "0" & "0" & "0" & bh7_w103_11_c2 & "0" & "0" & bh7_w100_14_c2 & "0" & "0" & bh7_w97_18_c2 & "0" & "0" & bh7_w94_18_c2 & "0" & bh7_w92_17_c2 & "0" & bh7_w90_21_c2 & "0" & bh7_w88_20_c2 & "0" & "0" & "0" & bh7_w84_20_c2 & "0" & bh7_w82_23_c2 & "0" & bh7_w80_23_c2 & "0" & "0" & bh7_w77_17_c2 & "0" & bh7_w75_18_c2 & "0" & bh7_w73_19_c2 & "0" & bh7_w71_19_c2 & "0" & "0" & bh7_w68_22_c2 & "0" & bh7_w66_23_c2 & "0" & bh7_w64_24_c2 & "0" & bh7_w62_22_c2 & "0" & bh7_w60_25_c2 & "0" & bh7_w58_24_c2 & "0" & bh7_w56_22_c2 & "0" & bh7_w54_21_c2 & "0" & bh7_w52_17_c2 & "0" & bh7_w50_12_c2 & "0" & bh7_w48_10_c2 & "0" & bh7_w46_9_c2 & "0" & bh7_w44_9_c2 & "0" & bh7_w42_9_c2 & "0" & bh7_w40_9_c2 & "0" & "0" & bh7_w37_7_c2 & "0" & bh7_w35_8_c2 & "0" & bh7_w33_6_c2 & "0" & bh7_w31_6_c2 & "0" & bh7_w29_6_c2 & "0" & bh7_w27_6_c2 & "0" & bh7_w25_6_c2 & "0" & bh7_w23_6_c2;
   bitheapFinalAdd_bh7_Cin_c0 <= '0';

   bitheapFinalAdd_bh7: IntAdder_84_Freq500_uid930
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 Cin => bitheapFinalAdd_bh7_Cin_c0,
                 X => bitheapFinalAdd_bh7_In0_c2,
                 Y => bitheapFinalAdd_bh7_In1_c2,
                 R => bitheapFinalAdd_bh7_Out_c4);
   bitheapResult_bh7_c4 <= bitheapFinalAdd_bh7_Out_c4(82 downto 0) & tmp_bitheapResult_bh7_22_c4;
   R <= bitheapResult_bh7_c4(105 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_65_Freq500_uid933
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_65_Freq500_uid933 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(64 downto 0);
          Y : in  std_logic_vector(64 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(64 downto 0)   );
end entity;

architecture arch of IntAdder_65_Freq500_uid933 is
signal Cin_0_c5, Cin_0_c6 :  std_logic;
signal X_0_c4, X_0_c5, X_0_c6 :  std_logic_vector(27 downto 0);
signal Y_0_c0, Y_0_c1, Y_0_c2, Y_0_c3, Y_0_c4, Y_0_c5, Y_0_c6 :  std_logic_vector(27 downto 0);
signal S_0_c6 :  std_logic_vector(27 downto 0);
signal R_0_c6 :  std_logic_vector(26 downto 0);
signal Cin_1_c6 :  std_logic;
signal X_1_c4, X_1_c5, X_1_c6 :  std_logic_vector(38 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3, Y_1_c4, Y_1_c5, Y_1_c6 :  std_logic_vector(38 downto 0);
signal S_1_c6 :  std_logic_vector(38 downto 0);
signal R_1_c6 :  std_logic_vector(37 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_0_c1 <= Y_0_c0;
               Y_1_c1 <= Y_1_c0;
            end if;
            if ce_2 = '1' then
               Y_0_c2 <= Y_0_c1;
               Y_1_c2 <= Y_1_c1;
            end if;
            if ce_3 = '1' then
               Y_0_c3 <= Y_0_c2;
               Y_1_c3 <= Y_1_c2;
            end if;
            if ce_4 = '1' then
               Y_0_c4 <= Y_0_c3;
               Y_1_c4 <= Y_1_c3;
            end if;
            if ce_5 = '1' then
               X_0_c5 <= X_0_c4;
               Y_0_c5 <= Y_0_c4;
               X_1_c5 <= X_1_c4;
               Y_1_c5 <= Y_1_c4;
            end if;
            if ce_6 = '1' then
               Cin_0_c6 <= Cin_0_c5;
               X_0_c6 <= X_0_c5;
               Y_0_c6 <= Y_0_c5;
               X_1_c6 <= X_1_c5;
               Y_1_c6 <= Y_1_c5;
            end if;
         end if;
      end process;
   Cin_0_c5 <= Cin;
   X_0_c4 <= '0' & X(26 downto 0);
   Y_0_c0 <= '0' & Y(26 downto 0);
   S_0_c6 <= X_0_c6 + Y_0_c6 + Cin_0_c6;
   R_0_c6 <= S_0_c6(26 downto 0);
   Cin_1_c6 <= S_0_c6(27);
   X_1_c4 <= '0' & X(64 downto 27);
   Y_1_c0 <= '0' & Y(64 downto 27);
   S_1_c6 <= X_1_c6 + Y_1_c6 + Cin_1_c6;
   R_1_c6 <= S_1_c6(37 downto 0);
   R <= R_1_c6 & R_0_c6 ;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointMultiplier
--                      (FPMult_11_52_uid2_Freq500_uid3)
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointMultiplier_64_2_758000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointMultiplier_64_2_758000 is
   component IntMultiplier_53x53_106_Freq500_uid5 is
      port ( clk, ce_1, ce_2, ce_3, ce_4 : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             Y : in  std_logic_vector(52 downto 0);
             R : out  std_logic_vector(105 downto 0)   );
   end component;

   component IntAdder_65_Freq500_uid933 is
      port ( clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
             X : in  std_logic_vector(64 downto 0);
             Y : in  std_logic_vector(64 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(64 downto 0)   );
   end component;

signal sign_c0, sign_c1, sign_c2, sign_c3, sign_c4, sign_c5, sign_c6 :  std_logic;
signal expX_c0 :  std_logic_vector(10 downto 0);
signal expY_c0 :  std_logic_vector(10 downto 0);
signal expSumPreSub_c0, expSumPreSub_c1 :  std_logic_vector(12 downto 0);
signal bias_c0, bias_c1 :  std_logic_vector(12 downto 0);
signal expSum_c1, expSum_c2, expSum_c3, expSum_c4 :  std_logic_vector(12 downto 0);
signal sigX_c0 :  std_logic_vector(52 downto 0);
signal sigY_c0 :  std_logic_vector(52 downto 0);
signal sigProd_c4 :  std_logic_vector(105 downto 0);
signal excSel_c0 :  std_logic_vector(3 downto 0);
signal exc_c0, exc_c1, exc_c2, exc_c3, exc_c4, exc_c5, exc_c6 :  std_logic_vector(1 downto 0);
signal norm_c4 :  std_logic;
signal expPostNorm_c4 :  std_logic_vector(12 downto 0);
signal sigProdExt_c4, sigProdExt_c5 :  std_logic_vector(105 downto 0);
signal expSig_c4 :  std_logic_vector(64 downto 0);
signal sticky_c4, sticky_c5 :  std_logic;
signal guard_c4, guard_c5 :  std_logic;
signal round_c5 :  std_logic;
signal expSigPostRound_c6 :  std_logic_vector(64 downto 0);
signal excPostNorm_c6 :  std_logic_vector(1 downto 0);
signal finalExc_c6 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               sign_c1 <= sign_c0;
               expSumPreSub_c1 <= expSumPreSub_c0;
               bias_c1 <= bias_c0;
               exc_c1 <= exc_c0;
            end if;
            if ce_2 = '1' then
               sign_c2 <= sign_c1;
               expSum_c2 <= expSum_c1;
               exc_c2 <= exc_c1;
            end if;
            if ce_3 = '1' then
               sign_c3 <= sign_c2;
               expSum_c3 <= expSum_c2;
               exc_c3 <= exc_c2;
            end if;
            if ce_4 = '1' then
               sign_c4 <= sign_c3;
               expSum_c4 <= expSum_c3;
               exc_c4 <= exc_c3;
            end if;
            if ce_5 = '1' then
               sign_c5 <= sign_c4;
               exc_c5 <= exc_c4;
               sigProdExt_c5 <= sigProdExt_c4;
               sticky_c5 <= sticky_c4;
               guard_c5 <= guard_c4;
            end if;
            if ce_6 = '1' then
               sign_c6 <= sign_c5;
               exc_c6 <= exc_c5;
            end if;
         end if;
      end process;
   sign_c0 <= X(63) xor Y(63);
   expX_c0 <= X(62 downto 52);
   expY_c0 <= Y(62 downto 52);
   expSumPreSub_c0 <= ("00" & expX_c0) + ("00" & expY_c0);
   bias_c0 <= CONV_STD_LOGIC_VECTOR(1023,13);
   expSum_c1 <= expSumPreSub_c1 - bias_c1;
   sigX_c0 <= "1" & X(51 downto 0);
   sigY_c0 <= "1" & Y(51 downto 0);
   SignificandMultiplication: IntMultiplier_53x53_106_Freq500_uid5
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 X => sigX_c0,
                 Y => sigY_c0,
                 R => sigProd_c4);
   excSel_c0 <= X(65 downto 64) & Y(65 downto 64);
   with excSel_c0  select  
   exc_c0 <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm_c4 <= sigProd_c4(105);
   -- exponent update
   expPostNorm_c4 <= expSum_c4 + ("000000000000" & norm_c4);
   -- significand normalization shift
   sigProdExt_c4 <= sigProd_c4(104 downto 0) & "0" when norm_c4='1' else
                         sigProd_c4(103 downto 0) & "00";
   expSig_c4 <= expPostNorm_c4 & sigProdExt_c4(105 downto 54);
   sticky_c4 <= sigProdExt_c4(53);
   guard_c4 <= '0' when sigProdExt_c4(52 downto 0)="00000000000000000000000000000000000000000000000000000" else '1';
   round_c5 <= sticky_c5 and ( (guard_c5 and not(sigProdExt_c5(54))) or (sigProdExt_c5(54) ))  ;
   RoundingAdder: IntAdder_65_Freq500_uid933
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 ce_4=> ce_4,
                 ce_5=> ce_5,
                 ce_6=> ce_6,
                 Cin => round_c5,
                 X => expSig_c4,
                 Y => "00000000000000000000000000000000000000000000000000000000000000000",
                 R => expSigPostRound_c6);
   with expSigPostRound_c6(64 downto 63)  select 
   excPostNorm_c6 <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_c6  select  
   finalExc_c6 <= exc_c6 when  "11"|"10"|"00",
                       excPostNorm_c6 when others; 
   R <= finalExc_c6 & sign_c6 & expSigPostRound_c6(62 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid17
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid17 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid17 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid22
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid22 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid22 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid27
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid27 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid27 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid32
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid32 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid32 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid37
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid37 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid37 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid42
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid42 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid42 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid47
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid47 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid47 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid52
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid52 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid52 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid63
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid63 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid63 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid68
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid68 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid68 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid73
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid73 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid73 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid78
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid78 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid78 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid83
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid83 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid83 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid88
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid88 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid88 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid93
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid93 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid93 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid98
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid98 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid98 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid113
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid113 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid113 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid118
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid118 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid118 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid123
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid123 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid123 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid128
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid128 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid128 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid133
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid133 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid133 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid138
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid138 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid138 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid143
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid143 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid143 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid148
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid148 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid148 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid153
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid153 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid153 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid158
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid158 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid158 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid163
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid163 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid163 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid168
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid168 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid168 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid183
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid183 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid183 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid188
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid188 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid188 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid193
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid193 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid193 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid198
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid198 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid198 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid203
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid203 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid203 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid208
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid208 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid208 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid213
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid213 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid213 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid218
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid218 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid218 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid223
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid223 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid223 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid228
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid228 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid228 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid233
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid233 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid233 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid238
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid238 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid238 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid253
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid253 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid253 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid258
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid258 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid258 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid263
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid263 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid263 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid268
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid268 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid268 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid273
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid273 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid273 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid278
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid278 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid278 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid283
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid283 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid283 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid288
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid288 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid288 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid293
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid293 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid293 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid298
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid298 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid298 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid303
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid303 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid303 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid308
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid308 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid308 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00000" when "00101",
      "00000" when "00110",
      "00000" when "00111",
      "00000" when "01000",
      "00001" when "01001",
      "00010" when "01010",
      "00011" when "01011",
      "00100" when "01100",
      "00101" when "01101",
      "00110" when "01110",
      "00111" when "01111",
      "00000" when "10000",
      "00010" when "10001",
      "00100" when "10010",
      "00110" when "10011",
      "01000" when "10100",
      "01010" when "10101",
      "01100" when "10110",
      "01110" when "10111",
      "00000" when "11000",
      "00011" when "11001",
      "00110" when "11010",
      "01001" when "11011",
      "01100" when "11100",
      "01111" when "11101",
      "10010" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid313
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid313 is
    port (X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid313 is
signal Y0 :  std_logic_vector(3 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(3 downto 0);
begin
   with X  select  Y0 <= 
      "0000" when "0000",
      "0000" when "0001",
      "0000" when "0010",
      "0000" when "0011",
      "0000" when "0100",
      "0001" when "0101",
      "0010" when "0110",
      "0011" when "0111",
      "0000" when "1000",
      "0010" when "1001",
      "0100" when "1010",
      "0110" when "1011",
      "0000" when "1100",
      "0011" when "1101",
      "0110" when "1110",
      "1001" when "1111",
      "----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          MultTable_Freq300_uid318
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity MultTable_Freq300_uid318 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of MultTable_Freq300_uid318 is
signal Y0 :  std_logic_vector(4 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(4 downto 0);
begin
   with X  select  Y0 <= 
      "00000" when "00000",
      "00000" when "00001",
      "00000" when "00010",
      "00000" when "00011",
      "00000" when "00100",
      "00001" when "00101",
      "00010" when "00110",
      "00011" when "00111",
      "00000" when "01000",
      "00010" when "01001",
      "00100" when "01010",
      "00110" when "01011",
      "00000" when "01100",
      "00011" when "01101",
      "00110" when "01110",
      "01001" when "01111",
      "00000" when "10000",
      "00100" when "10001",
      "01000" when "10010",
      "01100" when "10011",
      "00000" when "10100",
      "00101" when "10101",
      "01010" when "10110",
      "01111" when "10111",
      "00000" when "11000",
      "00110" when "11001",
      "01100" when "11010",
      "10010" when "11011",
      "00000" when "11100",
      "00111" when "11101",
      "01110" when "11110",
      "10101" when "11111",
      "-----" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq300_uid322
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq300_uid322 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq300_uid322 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq300_uid326
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq300_uid326 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq300_uid326 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_6_3_Freq300_uid334
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_Freq300_uid334 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_Freq300_uid334 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_5_3_Freq300_uid400
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3_Freq300_uid400 is
    port (X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3_Freq300_uid400 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000" | "10000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100" | "11000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "100" when "01111" | "10111" | "11011" | "11101" | "11110",
      "101" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_3_2_Freq300_uid432
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_Freq300_uid432 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_Freq300_uid432 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid9
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid9 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid9 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid11
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid11 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid11 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid13
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid13 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid13 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid15
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid15 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid15 is
   component MultTable_Freq300_uid17 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy18_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid17
      port map ( X => Xtable_c0,
                 Y => Y1_copy18_c0);
   Y1_c0 <= Y1_copy18_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid20
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid20 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid20 is
   component MultTable_Freq300_uid22 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy23_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid22
      port map ( X => Xtable_c0,
                 Y => Y1_copy23_c0);
   Y1_c0 <= Y1_copy23_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid25
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid25 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid25 is
   component MultTable_Freq300_uid27 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy28_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid27
      port map ( X => Xtable_c0,
                 Y => Y1_copy28_c0);
   Y1_c0 <= Y1_copy28_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid30
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid30 is
   component MultTable_Freq300_uid32 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy33_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid32
      port map ( X => Xtable_c0,
                 Y => Y1_copy33_c0);
   Y1_c0 <= Y1_copy33_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid35
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid35 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid35 is
   component MultTable_Freq300_uid37 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy38_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid37
      port map ( X => Xtable_c0,
                 Y => Y1_copy38_c0);
   Y1_c0 <= Y1_copy38_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid40
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid40 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid40 is
   component MultTable_Freq300_uid42 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy43_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid42
      port map ( X => Xtable_c0,
                 Y => Y1_copy43_c0);
   Y1_c0 <= Y1_copy43_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid45
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid45 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid45 is
   component MultTable_Freq300_uid47 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy48_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid47
      port map ( X => Xtable_c0,
                 Y => Y1_copy48_c0);
   Y1_c0 <= Y1_copy48_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid50
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid50 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid50 is
   component MultTable_Freq300_uid52 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy53_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid52
      port map ( X => Xtable_c0,
                 Y => Y1_copy53_c0);
   Y1_c0 <= Y1_copy53_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid55
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid55 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid55 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid57
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid57 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid57 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                        DSPBlock_17x24_Freq300_uid59
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_Freq300_uid59 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_Freq300_uid59 is
signal Mfull_c0 :  std_logic_vector(40 downto 0);
signal M_c0 :  std_logic_vector(40 downto 0);
begin
   Mfull_c0 <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M_c0 <= Mfull_c0(40 downto 0);
   R <= M_c0;
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid61
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid61 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid61 is
   component MultTable_Freq300_uid63 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy64_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid63
      port map ( X => Xtable_c0,
                 Y => Y1_copy64_c0);
   Y1_c0 <= Y1_copy64_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid66
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid66 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid66 is
   component MultTable_Freq300_uid68 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy69_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid68
      port map ( X => Xtable_c0,
                 Y => Y1_copy69_c0);
   Y1_c0 <= Y1_copy69_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid71
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid71 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid71 is
   component MultTable_Freq300_uid73 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy74_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid73
      port map ( X => Xtable_c0,
                 Y => Y1_copy74_c0);
   Y1_c0 <= Y1_copy74_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid76
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid76 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid76 is
   component MultTable_Freq300_uid78 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy79_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid78
      port map ( X => Xtable_c0,
                 Y => Y1_copy79_c0);
   Y1_c0 <= Y1_copy79_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid81
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid81 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid81 is
   component MultTable_Freq300_uid83 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy84_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid83
      port map ( X => Xtable_c0,
                 Y => Y1_copy84_c0);
   Y1_c0 <= Y1_copy84_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid86
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid86 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid86 is
   component MultTable_Freq300_uid88 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy89_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid88
      port map ( X => Xtable_c0,
                 Y => Y1_copy89_c0);
   Y1_c0 <= Y1_copy89_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid91
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid91 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid91 is
   component MultTable_Freq300_uid93 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy94_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid93
      port map ( X => Xtable_c0,
                 Y => Y1_copy94_c0);
   Y1_c0 <= Y1_copy94_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                     IntMultiplierLUT_2x3_Freq300_uid96
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid96 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid96 is
   component MultTable_Freq300_uid98 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy99_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid98
      port map ( X => Xtable_c0,
                 Y => Y1_copy99_c0);
   Y1_c0 <= Y1_copy99_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid101
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid101 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid101 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid103
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid103 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid103 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid105
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid105 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid105 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid107
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid107 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid107 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid109
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid109 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid109 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid111
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid111 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid111 is
   component MultTable_Freq300_uid113 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy114_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid113
      port map ( X => Xtable_c0,
                 Y => Y1_copy114_c0);
   Y1_c0 <= Y1_copy114_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid116
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid116 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid116 is
   component MultTable_Freq300_uid118 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy119_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid118
      port map ( X => Xtable_c0,
                 Y => Y1_copy119_c0);
   Y1_c0 <= Y1_copy119_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid121
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid121 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid121 is
   component MultTable_Freq300_uid123 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy124_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid123
      port map ( X => Xtable_c0,
                 Y => Y1_copy124_c0);
   Y1_c0 <= Y1_copy124_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid126
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid126 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid126 is
   component MultTable_Freq300_uid128 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy129_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid128
      port map ( X => Xtable_c0,
                 Y => Y1_copy129_c0);
   Y1_c0 <= Y1_copy129_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid131
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid131 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid131 is
   component MultTable_Freq300_uid133 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy134_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid133
      port map ( X => Xtable_c0,
                 Y => Y1_copy134_c0);
   Y1_c0 <= Y1_copy134_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid136
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid136 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid136 is
   component MultTable_Freq300_uid138 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy139_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid138
      port map ( X => Xtable_c0,
                 Y => Y1_copy139_c0);
   Y1_c0 <= Y1_copy139_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid141
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid141 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid141 is
   component MultTable_Freq300_uid143 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy144_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid143
      port map ( X => Xtable_c0,
                 Y => Y1_copy144_c0);
   Y1_c0 <= Y1_copy144_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid146
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid146 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid146 is
   component MultTable_Freq300_uid148 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy149_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid148
      port map ( X => Xtable_c0,
                 Y => Y1_copy149_c0);
   Y1_c0 <= Y1_copy149_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid151
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid151 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid151 is
   component MultTable_Freq300_uid153 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy154_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid153
      port map ( X => Xtable_c0,
                 Y => Y1_copy154_c0);
   Y1_c0 <= Y1_copy154_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid156
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid156 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid156 is
   component MultTable_Freq300_uid158 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy159_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid158
      port map ( X => Xtable_c0,
                 Y => Y1_copy159_c0);
   Y1_c0 <= Y1_copy159_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid161
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid161 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid161 is
   component MultTable_Freq300_uid163 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy164_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid163
      port map ( X => Xtable_c0,
                 Y => Y1_copy164_c0);
   Y1_c0 <= Y1_copy164_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid166
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid166 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid166 is
   component MultTable_Freq300_uid168 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy169_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid168
      port map ( X => Xtable_c0,
                 Y => Y1_copy169_c0);
   Y1_c0 <= Y1_copy169_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid171
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid171 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid171 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid173
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid173 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid173 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid175
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid175 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid175 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid177
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid177 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid177 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid179
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid179 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid179 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid181
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid181 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid181 is
   component MultTable_Freq300_uid183 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy184_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid183
      port map ( X => Xtable_c0,
                 Y => Y1_copy184_c0);
   Y1_c0 <= Y1_copy184_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid186
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid186 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid186 is
   component MultTable_Freq300_uid188 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy189_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid188
      port map ( X => Xtable_c0,
                 Y => Y1_copy189_c0);
   Y1_c0 <= Y1_copy189_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid191
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid191 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid191 is
   component MultTable_Freq300_uid193 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy194_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid193
      port map ( X => Xtable_c0,
                 Y => Y1_copy194_c0);
   Y1_c0 <= Y1_copy194_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid196
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid196 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid196 is
   component MultTable_Freq300_uid198 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy199_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid198
      port map ( X => Xtable_c0,
                 Y => Y1_copy199_c0);
   Y1_c0 <= Y1_copy199_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid201
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid201 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid201 is
   component MultTable_Freq300_uid203 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy204_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid203
      port map ( X => Xtable_c0,
                 Y => Y1_copy204_c0);
   Y1_c0 <= Y1_copy204_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid206
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid206 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid206 is
   component MultTable_Freq300_uid208 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy209_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid208
      port map ( X => Xtable_c0,
                 Y => Y1_copy209_c0);
   Y1_c0 <= Y1_copy209_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid211
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid211 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid211 is
   component MultTable_Freq300_uid213 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy214_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid213
      port map ( X => Xtable_c0,
                 Y => Y1_copy214_c0);
   Y1_c0 <= Y1_copy214_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid216
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid216 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid216 is
   component MultTable_Freq300_uid218 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy219_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid218
      port map ( X => Xtable_c0,
                 Y => Y1_copy219_c0);
   Y1_c0 <= Y1_copy219_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid221
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid221 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid221 is
   component MultTable_Freq300_uid223 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy224_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid223
      port map ( X => Xtable_c0,
                 Y => Y1_copy224_c0);
   Y1_c0 <= Y1_copy224_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid226
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid226 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid226 is
   component MultTable_Freq300_uid228 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy229_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid228
      port map ( X => Xtable_c0,
                 Y => Y1_copy229_c0);
   Y1_c0 <= Y1_copy229_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid231
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid231 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid231 is
   component MultTable_Freq300_uid233 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy234_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid233
      port map ( X => Xtable_c0,
                 Y => Y1_copy234_c0);
   Y1_c0 <= Y1_copy234_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid236
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid236 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid236 is
   component MultTable_Freq300_uid238 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy239_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid238
      port map ( X => Xtable_c0,
                 Y => Y1_copy239_c0);
   Y1_c0 <= Y1_copy239_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_1x1_Freq300_uid241
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_1x1_Freq300_uid241 is
    port (clk : in std_logic;
          X : in  std_logic_vector(0 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(0 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_1x1_Freq300_uid241 is
signal replicated_c0 :  std_logic_vector(0 downto 0);
signal prod_c0 :  std_logic_vector(0 downto 0);
begin
   replicated_c0 <= (0 downto 0 => X(0));
   prod_c0 <= Y and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid243
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid243 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid243 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid245
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid245 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid245 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid247
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid247 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid247 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_4x1_Freq300_uid249
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_4x1_Freq300_uid249 is
    port (clk : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_4x1_Freq300_uid249 is
signal replicated_c0 :  std_logic_vector(3 downto 0);
signal prod_c0 :  std_logic_vector(3 downto 0);
begin
   replicated_c0 <= (3 downto 0 => Y(0));
   prod_c0 <= X and replicated_c0;
   R <= prod_c0;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid251
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid251 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid251 is
   component MultTable_Freq300_uid253 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy254_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid253
      port map ( X => Xtable_c0,
                 Y => Y1_copy254_c0);
   Y1_c0 <= Y1_copy254_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid256
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid256 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid256 is
   component MultTable_Freq300_uid258 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy259_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid258
      port map ( X => Xtable_c0,
                 Y => Y1_copy259_c0);
   Y1_c0 <= Y1_copy259_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid261
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid261 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid261 is
   component MultTable_Freq300_uid263 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy264_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid263
      port map ( X => Xtable_c0,
                 Y => Y1_copy264_c0);
   Y1_c0 <= Y1_copy264_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid266
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid266 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid266 is
   component MultTable_Freq300_uid268 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy269_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid268
      port map ( X => Xtable_c0,
                 Y => Y1_copy269_c0);
   Y1_c0 <= Y1_copy269_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid271
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid271 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid271 is
   component MultTable_Freq300_uid273 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy274_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid273
      port map ( X => Xtable_c0,
                 Y => Y1_copy274_c0);
   Y1_c0 <= Y1_copy274_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid276
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid276 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid276 is
   component MultTable_Freq300_uid278 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy279_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid278
      port map ( X => Xtable_c0,
                 Y => Y1_copy279_c0);
   Y1_c0 <= Y1_copy279_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid281
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid281 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid281 is
   component MultTable_Freq300_uid283 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy284_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid283
      port map ( X => Xtable_c0,
                 Y => Y1_copy284_c0);
   Y1_c0 <= Y1_copy284_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid286
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid286 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid286 is
   component MultTable_Freq300_uid288 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy289_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid288
      port map ( X => Xtable_c0,
                 Y => Y1_copy289_c0);
   Y1_c0 <= Y1_copy289_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid291
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid291 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid291 is
   component MultTable_Freq300_uid293 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy294_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid293
      port map ( X => Xtable_c0,
                 Y => Y1_copy294_c0);
   Y1_c0 <= Y1_copy294_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid296
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid296 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid296 is
   component MultTable_Freq300_uid298 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy299_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid298
      port map ( X => Xtable_c0,
                 Y => Y1_copy299_c0);
   Y1_c0 <= Y1_copy299_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid301
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid301 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid301 is
   component MultTable_Freq300_uid303 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy304_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid303
      port map ( X => Xtable_c0,
                 Y => Y1_copy304_c0);
   Y1_c0 <= Y1_copy304_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_3x2_Freq300_uid306
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_3x2_Freq300_uid306 is
    port (clk : in std_logic;
          X : in  std_logic_vector(2 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_3x2_Freq300_uid306 is
   component MultTable_Freq300_uid308 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy309_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid308
      port map ( X => Xtable_c0,
                 Y => Y1_copy309_c0);
   Y1_c0 <= Y1_copy309_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x2_Freq300_uid311
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x2_Freq300_uid311 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x2_Freq300_uid311 is
   component MultTable_Freq300_uid313 is
      port ( X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(3 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(3 downto 0);
signal Y1_c0 :  std_logic_vector(3 downto 0);
signal Y1_copy314_c0 :  std_logic_vector(3 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid313
      port map ( X => Xtable_c0,
                 Y => Y1_copy314_c0);
   Y1_c0 <= Y1_copy314_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplierLUT_2x3_Freq300_uid316
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntMultiplierLUT_2x3_Freq300_uid316 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1 downto 0);
          Y : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(4 downto 0)   );
end entity;

architecture arch of IntMultiplierLUT_2x3_Freq300_uid316 is
   component MultTable_Freq300_uid318 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(4 downto 0)   );
   end component;

signal Xtable_c0 :  std_logic_vector(4 downto 0);
signal Y1_c0 :  std_logic_vector(4 downto 0);
signal Y1_copy319_c0 :  std_logic_vector(4 downto 0);
begin
Xtable_c0 <= Y & X;
   R <= Y1_c0;
   TableMult: MultTable_Freq300_uid318
      port map ( X => Xtable_c0,
                 Y => Y1_copy319_c0);
   Y1_c0 <= Y1_copy319_c0; -- output copy to hold a pipeline register if needed
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_84_Freq300_uid972
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_84_Freq300_uid972 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(83 downto 0);
          Y : in  std_logic_vector(83 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(83 downto 0)   );
end entity;

architecture arch of IntAdder_84_Freq300_uid972 is
signal Rtmp_c2 :  std_logic_vector(83 downto 0);
signal X_c2 :  std_logic_vector(83 downto 0);
signal Y_c2 :  std_logic_vector(83 downto 0);
signal Cin_c1, Cin_c2 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Cin_c1 <= Cin;
            end if;
            if ce_2 = '1' then
               X_c2 <= X;
               Y_c2 <= Y;
               Cin_c2 <= Cin_c1;
            end if;
         end if;
      end process;
   Rtmp_c2 <= X_c2 + Y_c2 + Cin_c2;
   R <= Rtmp_c2;
end architecture;

--------------------------------------------------------------------------------
--                    IntMultiplier_53x53_106_Freq300_uid5
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012-
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_53x53_106_Freq300_uid5 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(52 downto 0);
          Y : in  std_logic_vector(52 downto 0);
          R : out  std_logic_vector(105 downto 0)   );
end entity;

architecture arch of IntMultiplier_53x53_106_Freq300_uid5 is
   component DSPBlock_17x24_Freq300_uid9 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid11 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid13 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid15 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid20 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid25 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid35 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid40 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid45 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid50 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid55 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid57 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_Freq300_uid59 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid61 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid66 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid71 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid76 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid81 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid86 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid91 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid96 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid101 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid103 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid105 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid107 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid109 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid111 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid116 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid121 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid126 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid131 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid136 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid141 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid146 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid151 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid156 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid161 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid166 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid171 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid173 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid175 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid177 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid179 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid181 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid186 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid191 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid196 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid201 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid206 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid211 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid216 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid221 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid226 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid231 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid236 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_1x1_Freq300_uid241 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(0 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(0 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid243 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid245 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid247 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_4x1_Freq300_uid249 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid251 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid256 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid261 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid266 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid271 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid276 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid281 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid286 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid291 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid296 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid301 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_3x2_Freq300_uid306 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(2 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component IntMultiplierLUT_2x2_Freq300_uid311 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(3 downto 0)   );
   end component;

   component IntMultiplierLUT_2x3_Freq300_uid316 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1 downto 0);
             Y : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(4 downto 0)   );
   end component;

   component Compressor_23_3_Freq300_uid322 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq300_uid326 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_Freq300_uid334 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3_Freq300_uid400 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_Freq300_uid432 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component IntAdder_84_Freq300_uid972 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(83 downto 0);
             Y : in  std_logic_vector(83 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(83 downto 0)   );
   end component;

signal XX_m6_c0 :  std_logic_vector(52 downto 0);
signal YY_m6_c0 :  std_logic_vector(52 downto 0);
signal tile_0_X_c0 :  std_logic_vector(16 downto 0);
signal tile_0_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_0_output_c0 :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w0_0_c0, bh7_w0_0_c1 :  std_logic;
signal bh7_w1_0_c0, bh7_w1_0_c1 :  std_logic;
signal bh7_w2_0_c0, bh7_w2_0_c1 :  std_logic;
signal bh7_w3_0_c0, bh7_w3_0_c1 :  std_logic;
signal bh7_w4_0_c0, bh7_w4_0_c1 :  std_logic;
signal bh7_w5_0_c0, bh7_w5_0_c1 :  std_logic;
signal bh7_w6_0_c0, bh7_w6_0_c1 :  std_logic;
signal bh7_w7_0_c0, bh7_w7_0_c1 :  std_logic;
signal bh7_w8_0_c0, bh7_w8_0_c1 :  std_logic;
signal bh7_w9_0_c0, bh7_w9_0_c1 :  std_logic;
signal bh7_w10_0_c0, bh7_w10_0_c1 :  std_logic;
signal bh7_w11_0_c0, bh7_w11_0_c1 :  std_logic;
signal bh7_w12_0_c0, bh7_w12_0_c1 :  std_logic;
signal bh7_w13_0_c0, bh7_w13_0_c1 :  std_logic;
signal bh7_w14_0_c0, bh7_w14_0_c1 :  std_logic;
signal bh7_w15_0_c0, bh7_w15_0_c1 :  std_logic;
signal bh7_w16_0_c0, bh7_w16_0_c1 :  std_logic;
signal bh7_w17_0_c0 :  std_logic;
signal bh7_w18_0_c0 :  std_logic;
signal bh7_w19_0_c0 :  std_logic;
signal bh7_w20_0_c0 :  std_logic;
signal bh7_w21_0_c0 :  std_logic;
signal bh7_w22_0_c0 :  std_logic;
signal bh7_w23_0_c0 :  std_logic;
signal bh7_w24_0_c0 :  std_logic;
signal bh7_w25_0_c0 :  std_logic;
signal bh7_w26_0_c0 :  std_logic;
signal bh7_w27_0_c0 :  std_logic;
signal bh7_w28_0_c0 :  std_logic;
signal bh7_w29_0_c0 :  std_logic;
signal bh7_w30_0_c0 :  std_logic;
signal bh7_w31_0_c0 :  std_logic;
signal bh7_w32_0_c0 :  std_logic;
signal bh7_w33_0_c0 :  std_logic;
signal bh7_w34_0_c0 :  std_logic;
signal bh7_w35_0_c0 :  std_logic;
signal bh7_w36_0_c0 :  std_logic;
signal bh7_w37_0_c0 :  std_logic;
signal bh7_w38_0_c0 :  std_logic;
signal bh7_w39_0_c0 :  std_logic;
signal bh7_w40_0_c0 :  std_logic;
signal tile_1_X_c0 :  std_logic_vector(16 downto 0);
signal tile_1_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_1_output_c0 :  std_logic_vector(40 downto 0);
signal tile_1_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w17_1_c0 :  std_logic;
signal bh7_w18_1_c0 :  std_logic;
signal bh7_w19_1_c0 :  std_logic;
signal bh7_w20_1_c0 :  std_logic;
signal bh7_w21_1_c0 :  std_logic;
signal bh7_w22_1_c0 :  std_logic;
signal bh7_w23_1_c0 :  std_logic;
signal bh7_w24_1_c0 :  std_logic;
signal bh7_w25_1_c0 :  std_logic;
signal bh7_w26_1_c0 :  std_logic;
signal bh7_w27_1_c0 :  std_logic;
signal bh7_w28_1_c0 :  std_logic;
signal bh7_w29_1_c0 :  std_logic;
signal bh7_w30_1_c0 :  std_logic;
signal bh7_w31_1_c0 :  std_logic;
signal bh7_w32_1_c0 :  std_logic;
signal bh7_w33_1_c0 :  std_logic;
signal bh7_w34_1_c0 :  std_logic;
signal bh7_w35_1_c0 :  std_logic;
signal bh7_w36_1_c0 :  std_logic;
signal bh7_w37_1_c0 :  std_logic;
signal bh7_w38_1_c0 :  std_logic;
signal bh7_w39_1_c0 :  std_logic;
signal bh7_w40_1_c0 :  std_logic;
signal bh7_w41_0_c0 :  std_logic;
signal bh7_w42_0_c0 :  std_logic;
signal bh7_w43_0_c0 :  std_logic;
signal bh7_w44_0_c0 :  std_logic;
signal bh7_w45_0_c0 :  std_logic;
signal bh7_w46_0_c0 :  std_logic;
signal bh7_w47_0_c0 :  std_logic;
signal bh7_w48_0_c0 :  std_logic;
signal bh7_w49_0_c0 :  std_logic;
signal bh7_w50_0_c0 :  std_logic;
signal bh7_w51_0_c0 :  std_logic;
signal bh7_w52_0_c0 :  std_logic;
signal bh7_w53_0_c0 :  std_logic;
signal bh7_w54_0_c0 :  std_logic;
signal bh7_w55_0_c0 :  std_logic;
signal bh7_w56_0_c0 :  std_logic;
signal bh7_w57_0_c0 :  std_logic;
signal tile_2_X_c0 :  std_logic_vector(16 downto 0);
signal tile_2_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_2_output_c0 :  std_logic_vector(40 downto 0);
signal tile_2_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w34_2_c0 :  std_logic;
signal bh7_w35_2_c0 :  std_logic;
signal bh7_w36_2_c0 :  std_logic;
signal bh7_w37_2_c0 :  std_logic;
signal bh7_w38_2_c0 :  std_logic;
signal bh7_w39_2_c0 :  std_logic;
signal bh7_w40_2_c0 :  std_logic;
signal bh7_w41_1_c0 :  std_logic;
signal bh7_w42_1_c0 :  std_logic;
signal bh7_w43_1_c0 :  std_logic;
signal bh7_w44_1_c0 :  std_logic;
signal bh7_w45_1_c0 :  std_logic;
signal bh7_w46_1_c0 :  std_logic;
signal bh7_w47_1_c0 :  std_logic;
signal bh7_w48_1_c0 :  std_logic;
signal bh7_w49_1_c0 :  std_logic;
signal bh7_w50_1_c0 :  std_logic;
signal bh7_w51_1_c0 :  std_logic;
signal bh7_w52_1_c0 :  std_logic;
signal bh7_w53_1_c0 :  std_logic;
signal bh7_w54_1_c0 :  std_logic;
signal bh7_w55_1_c0 :  std_logic;
signal bh7_w56_1_c0 :  std_logic;
signal bh7_w57_1_c0 :  std_logic;
signal bh7_w58_0_c0 :  std_logic;
signal bh7_w59_0_c0, bh7_w59_0_c1 :  std_logic;
signal bh7_w60_0_c0, bh7_w60_0_c1 :  std_logic;
signal bh7_w61_0_c0, bh7_w61_0_c1 :  std_logic;
signal bh7_w62_0_c0, bh7_w62_0_c1 :  std_logic;
signal bh7_w63_0_c0 :  std_logic;
signal bh7_w64_0_c0, bh7_w64_0_c1 :  std_logic;
signal bh7_w65_0_c0, bh7_w65_0_c1 :  std_logic;
signal bh7_w66_0_c0 :  std_logic;
signal bh7_w67_0_c0, bh7_w67_0_c1 :  std_logic;
signal bh7_w68_0_c0 :  std_logic;
signal bh7_w69_0_c0, bh7_w69_0_c1 :  std_logic;
signal bh7_w70_0_c0, bh7_w70_0_c1 :  std_logic;
signal bh7_w71_0_c0 :  std_logic;
signal bh7_w72_0_c0, bh7_w72_0_c1 :  std_logic;
signal bh7_w73_0_c0 :  std_logic;
signal bh7_w74_0_c0, bh7_w74_0_c1 :  std_logic;
signal tile_3_X_c0 :  std_logic_vector(1 downto 0);
signal tile_3_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_3_output_c0 :  std_logic_vector(4 downto 0);
signal tile_3_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w72_1_c0 :  std_logic;
signal bh7_w73_1_c0 :  std_logic;
signal bh7_w74_1_c0 :  std_logic;
signal bh7_w75_0_c0 :  std_logic;
signal bh7_w76_0_c0 :  std_logic;
signal tile_4_X_c0 :  std_logic_vector(1 downto 0);
signal tile_4_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_4_output_c0 :  std_logic_vector(4 downto 0);
signal tile_4_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w69_1_c0 :  std_logic;
signal bh7_w70_1_c0 :  std_logic;
signal bh7_w71_1_c0 :  std_logic;
signal bh7_w72_2_c0 :  std_logic;
signal bh7_w73_2_c0 :  std_logic;
signal tile_5_X_c0 :  std_logic_vector(1 downto 0);
signal tile_5_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_5_output_c0 :  std_logic_vector(4 downto 0);
signal tile_5_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w66_1_c0 :  std_logic;
signal bh7_w67_1_c0 :  std_logic;
signal bh7_w68_1_c0 :  std_logic;
signal bh7_w69_2_c0 :  std_logic;
signal bh7_w70_2_c0 :  std_logic;
signal tile_6_X_c0 :  std_logic_vector(1 downto 0);
signal tile_6_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_6_output_c0 :  std_logic_vector(4 downto 0);
signal tile_6_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w63_1_c0 :  std_logic;
signal bh7_w64_1_c0 :  std_logic;
signal bh7_w65_1_c0 :  std_logic;
signal bh7_w66_2_c0 :  std_logic;
signal bh7_w67_2_c0 :  std_logic;
signal tile_7_X_c0 :  std_logic_vector(1 downto 0);
signal tile_7_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_7_output_c0 :  std_logic_vector(4 downto 0);
signal tile_7_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_1_c0 :  std_logic;
signal bh7_w61_1_c0 :  std_logic;
signal bh7_w62_1_c0 :  std_logic;
signal bh7_w63_2_c0 :  std_logic;
signal bh7_w64_2_c0 :  std_logic;
signal tile_8_X_c0 :  std_logic_vector(1 downto 0);
signal tile_8_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_8_output_c0 :  std_logic_vector(4 downto 0);
signal tile_8_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_2_c0 :  std_logic;
signal bh7_w58_1_c0 :  std_logic;
signal bh7_w59_1_c0 :  std_logic;
signal bh7_w60_2_c0 :  std_logic;
signal bh7_w61_2_c0 :  std_logic;
signal tile_9_X_c0 :  std_logic_vector(1 downto 0);
signal tile_9_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_9_output_c0 :  std_logic_vector(4 downto 0);
signal tile_9_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_2_c0 :  std_logic;
signal bh7_w55_2_c0 :  std_logic;
signal bh7_w56_2_c0 :  std_logic;
signal bh7_w57_3_c0 :  std_logic;
signal bh7_w58_2_c0 :  std_logic;
signal tile_10_X_c0 :  std_logic_vector(1 downto 0);
signal tile_10_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_10_output_c0 :  std_logic_vector(4 downto 0);
signal tile_10_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_2_c0 :  std_logic;
signal bh7_w52_2_c0 :  std_logic;
signal bh7_w53_2_c0 :  std_logic;
signal bh7_w54_3_c0 :  std_logic;
signal bh7_w55_3_c0 :  std_logic;
signal tile_11_X_c0 :  std_logic_vector(16 downto 0);
signal tile_11_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_11_output_c0 :  std_logic_vector(40 downto 0);
signal tile_11_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w24_2_c0 :  std_logic;
signal bh7_w25_2_c0, bh7_w25_2_c1 :  std_logic;
signal bh7_w26_2_c0 :  std_logic;
signal bh7_w27_2_c0, bh7_w27_2_c1 :  std_logic;
signal bh7_w28_2_c0 :  std_logic;
signal bh7_w29_2_c0, bh7_w29_2_c1 :  std_logic;
signal bh7_w30_2_c0 :  std_logic;
signal bh7_w31_2_c0, bh7_w31_2_c1 :  std_logic;
signal bh7_w32_2_c0 :  std_logic;
signal bh7_w33_2_c0, bh7_w33_2_c1 :  std_logic;
signal bh7_w34_3_c0 :  std_logic;
signal bh7_w35_3_c0 :  std_logic;
signal bh7_w36_3_c0 :  std_logic;
signal bh7_w37_3_c0 :  std_logic;
signal bh7_w38_3_c0 :  std_logic;
signal bh7_w39_3_c0 :  std_logic;
signal bh7_w40_3_c0 :  std_logic;
signal bh7_w41_2_c0 :  std_logic;
signal bh7_w42_2_c0 :  std_logic;
signal bh7_w43_2_c0 :  std_logic;
signal bh7_w44_2_c0 :  std_logic;
signal bh7_w45_2_c0 :  std_logic;
signal bh7_w46_2_c0 :  std_logic;
signal bh7_w47_2_c0 :  std_logic;
signal bh7_w48_2_c0 :  std_logic;
signal bh7_w49_2_c0 :  std_logic;
signal bh7_w50_2_c0 :  std_logic;
signal bh7_w51_3_c0 :  std_logic;
signal bh7_w52_3_c0 :  std_logic;
signal bh7_w53_3_c0 :  std_logic;
signal bh7_w54_4_c0 :  std_logic;
signal bh7_w55_4_c0 :  std_logic;
signal bh7_w56_3_c0 :  std_logic;
signal bh7_w57_4_c0 :  std_logic;
signal bh7_w58_3_c0 :  std_logic;
signal bh7_w59_2_c0, bh7_w59_2_c1 :  std_logic;
signal bh7_w60_3_c0, bh7_w60_3_c1 :  std_logic;
signal bh7_w61_3_c0, bh7_w61_3_c1 :  std_logic;
signal bh7_w62_2_c0, bh7_w62_2_c1 :  std_logic;
signal bh7_w63_3_c0 :  std_logic;
signal bh7_w64_3_c0, bh7_w64_3_c1 :  std_logic;
signal tile_12_X_c0 :  std_logic_vector(16 downto 0);
signal tile_12_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_12_output_c0 :  std_logic_vector(40 downto 0);
signal tile_12_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w41_3_c0 :  std_logic;
signal bh7_w42_3_c0 :  std_logic;
signal bh7_w43_3_c0 :  std_logic;
signal bh7_w44_3_c0 :  std_logic;
signal bh7_w45_3_c0 :  std_logic;
signal bh7_w46_3_c0 :  std_logic;
signal bh7_w47_3_c0 :  std_logic;
signal bh7_w48_3_c0, bh7_w48_3_c1 :  std_logic;
signal bh7_w49_3_c0 :  std_logic;
signal bh7_w50_3_c0 :  std_logic;
signal bh7_w51_4_c0 :  std_logic;
signal bh7_w52_4_c0 :  std_logic;
signal bh7_w53_4_c0 :  std_logic;
signal bh7_w54_5_c0 :  std_logic;
signal bh7_w55_5_c0 :  std_logic;
signal bh7_w56_4_c0 :  std_logic;
signal bh7_w57_5_c0 :  std_logic;
signal bh7_w58_4_c0 :  std_logic;
signal bh7_w59_3_c0, bh7_w59_3_c1 :  std_logic;
signal bh7_w60_4_c0, bh7_w60_4_c1 :  std_logic;
signal bh7_w61_4_c0, bh7_w61_4_c1 :  std_logic;
signal bh7_w62_3_c0, bh7_w62_3_c1 :  std_logic;
signal bh7_w63_4_c0 :  std_logic;
signal bh7_w64_4_c0, bh7_w64_4_c1 :  std_logic;
signal bh7_w65_2_c0, bh7_w65_2_c1 :  std_logic;
signal bh7_w66_3_c0 :  std_logic;
signal bh7_w67_3_c0, bh7_w67_3_c1 :  std_logic;
signal bh7_w68_2_c0 :  std_logic;
signal bh7_w69_3_c0, bh7_w69_3_c1 :  std_logic;
signal bh7_w70_3_c0, bh7_w70_3_c1 :  std_logic;
signal bh7_w71_2_c0 :  std_logic;
signal bh7_w72_3_c0, bh7_w72_3_c1 :  std_logic;
signal bh7_w73_3_c0 :  std_logic;
signal bh7_w74_2_c0, bh7_w74_2_c1 :  std_logic;
signal bh7_w75_1_c0 :  std_logic;
signal bh7_w76_1_c0, bh7_w76_1_c1 :  std_logic;
signal bh7_w77_0_c0, bh7_w77_0_c1 :  std_logic;
signal bh7_w78_0_c0, bh7_w78_0_c1 :  std_logic;
signal bh7_w79_0_c0, bh7_w79_0_c1 :  std_logic;
signal bh7_w80_0_c0, bh7_w80_0_c1 :  std_logic;
signal bh7_w81_0_c0, bh7_w81_0_c1 :  std_logic;
signal tile_13_X_c0 :  std_logic_vector(16 downto 0);
signal tile_13_Y_c0 :  std_logic_vector(23 downto 0);
signal tile_13_output_c0 :  std_logic_vector(40 downto 0);
signal tile_13_filtered_output_c0 :  unsigned(40-0 downto 0);
signal bh7_w58_5_c0, bh7_w58_5_c1 :  std_logic;
signal bh7_w59_4_c0, bh7_w59_4_c1 :  std_logic;
signal bh7_w60_5_c0, bh7_w60_5_c1 :  std_logic;
signal bh7_w61_5_c0, bh7_w61_5_c1 :  std_logic;
signal bh7_w62_4_c0, bh7_w62_4_c1 :  std_logic;
signal bh7_w63_5_c0, bh7_w63_5_c1 :  std_logic;
signal bh7_w64_5_c0, bh7_w64_5_c1 :  std_logic;
signal bh7_w65_3_c0, bh7_w65_3_c1 :  std_logic;
signal bh7_w66_4_c0 :  std_logic;
signal bh7_w67_4_c0, bh7_w67_4_c1 :  std_logic;
signal bh7_w68_3_c0 :  std_logic;
signal bh7_w69_4_c0, bh7_w69_4_c1 :  std_logic;
signal bh7_w70_4_c0, bh7_w70_4_c1 :  std_logic;
signal bh7_w71_3_c0 :  std_logic;
signal bh7_w72_4_c0, bh7_w72_4_c1 :  std_logic;
signal bh7_w73_4_c0 :  std_logic;
signal bh7_w74_3_c0, bh7_w74_3_c1 :  std_logic;
signal bh7_w75_2_c0, bh7_w75_2_c1 :  std_logic;
signal bh7_w76_2_c0, bh7_w76_2_c1 :  std_logic;
signal bh7_w77_1_c0, bh7_w77_1_c1 :  std_logic;
signal bh7_w78_1_c0, bh7_w78_1_c1 :  std_logic;
signal bh7_w79_1_c0, bh7_w79_1_c1 :  std_logic;
signal bh7_w80_1_c0, bh7_w80_1_c1 :  std_logic;
signal bh7_w81_1_c0, bh7_w81_1_c1 :  std_logic;
signal bh7_w82_0_c0, bh7_w82_0_c1 :  std_logic;
signal bh7_w83_0_c0, bh7_w83_0_c1 :  std_logic;
signal bh7_w84_0_c0, bh7_w84_0_c1 :  std_logic;
signal bh7_w85_0_c0, bh7_w85_0_c1 :  std_logic;
signal bh7_w86_0_c0, bh7_w86_0_c1 :  std_logic;
signal bh7_w87_0_c0, bh7_w87_0_c1 :  std_logic;
signal bh7_w88_0_c0, bh7_w88_0_c1 :  std_logic;
signal bh7_w89_0_c0, bh7_w89_0_c1 :  std_logic;
signal bh7_w90_0_c0, bh7_w90_0_c1 :  std_logic;
signal bh7_w91_0_c0, bh7_w91_0_c1 :  std_logic;
signal bh7_w92_0_c0, bh7_w92_0_c1 :  std_logic;
signal bh7_w93_0_c0, bh7_w93_0_c1 :  std_logic;
signal bh7_w94_0_c0, bh7_w94_0_c1 :  std_logic;
signal bh7_w95_0_c0, bh7_w95_0_c1 :  std_logic;
signal bh7_w96_0_c0, bh7_w96_0_c1 :  std_logic;
signal bh7_w97_0_c0, bh7_w97_0_c1 :  std_logic;
signal bh7_w98_0_c0, bh7_w98_0_c1 :  std_logic;
signal tile_14_X_c0 :  std_logic_vector(1 downto 0);
signal tile_14_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_14_output_c0 :  std_logic_vector(4 downto 0);
signal tile_14_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_1_c0 :  std_logic;
signal bh7_w97_1_c0 :  std_logic;
signal bh7_w98_1_c0 :  std_logic;
signal bh7_w99_0_c0 :  std_logic;
signal bh7_w100_0_c0 :  std_logic;
signal tile_15_X_c0 :  std_logic_vector(1 downto 0);
signal tile_15_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_15_output_c0 :  std_logic_vector(4 downto 0);
signal tile_15_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_1_c0 :  std_logic;
signal bh7_w94_1_c0 :  std_logic;
signal bh7_w95_1_c0 :  std_logic;
signal bh7_w96_2_c0 :  std_logic;
signal bh7_w97_2_c0 :  std_logic;
signal tile_16_X_c0 :  std_logic_vector(1 downto 0);
signal tile_16_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_16_output_c0 :  std_logic_vector(4 downto 0);
signal tile_16_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_1_c0 :  std_logic;
signal bh7_w91_1_c0 :  std_logic;
signal bh7_w92_1_c0 :  std_logic;
signal bh7_w93_2_c0 :  std_logic;
signal bh7_w94_2_c0 :  std_logic;
signal tile_17_X_c0 :  std_logic_vector(1 downto 0);
signal tile_17_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_17_output_c0 :  std_logic_vector(4 downto 0);
signal tile_17_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_1_c0 :  std_logic;
signal bh7_w88_1_c0 :  std_logic;
signal bh7_w89_1_c0 :  std_logic;
signal bh7_w90_2_c0 :  std_logic;
signal bh7_w91_2_c0 :  std_logic;
signal tile_18_X_c0 :  std_logic_vector(1 downto 0);
signal tile_18_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_18_output_c0 :  std_logic_vector(4 downto 0);
signal tile_18_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_1_c0 :  std_logic;
signal bh7_w85_1_c0 :  std_logic;
signal bh7_w86_1_c0 :  std_logic;
signal bh7_w87_2_c0 :  std_logic;
signal bh7_w88_2_c0 :  std_logic;
signal tile_19_X_c0 :  std_logic_vector(1 downto 0);
signal tile_19_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_19_output_c0 :  std_logic_vector(4 downto 0);
signal tile_19_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w81_2_c0 :  std_logic;
signal bh7_w82_1_c0 :  std_logic;
signal bh7_w83_1_c0 :  std_logic;
signal bh7_w84_2_c0 :  std_logic;
signal bh7_w85_2_c0 :  std_logic;
signal tile_20_X_c0 :  std_logic_vector(1 downto 0);
signal tile_20_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_20_output_c0 :  std_logic_vector(4 downto 0);
signal tile_20_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w78_2_c0 :  std_logic;
signal bh7_w79_2_c0 :  std_logic;
signal bh7_w80_2_c0 :  std_logic;
signal bh7_w81_3_c0 :  std_logic;
signal bh7_w82_2_c0 :  std_logic;
signal tile_21_X_c0 :  std_logic_vector(1 downto 0);
signal tile_21_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_21_output_c0 :  std_logic_vector(4 downto 0);
signal tile_21_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w75_3_c0 :  std_logic;
signal bh7_w76_3_c0 :  std_logic;
signal bh7_w77_2_c0 :  std_logic;
signal bh7_w78_3_c0 :  std_logic;
signal bh7_w79_3_c0 :  std_logic;
signal tile_22_X_c0 :  std_logic_vector(0 downto 0);
signal tile_22_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_22_output_c0 :  std_logic_vector(0 downto 0);
signal tile_22_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w68_4_c0 :  std_logic;
signal tile_23_X_c0 :  std_logic_vector(3 downto 0);
signal tile_23_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_23_output_c0 :  std_logic_vector(3 downto 0);
signal tile_23_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w64_6_c0 :  std_logic;
signal bh7_w65_4_c0 :  std_logic;
signal bh7_w66_5_c0 :  std_logic;
signal bh7_w67_5_c0 :  std_logic;
signal tile_24_X_c0 :  std_logic_vector(3 downto 0);
signal tile_24_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_24_output_c0 :  std_logic_vector(3 downto 0);
signal tile_24_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w60_6_c0 :  std_logic;
signal bh7_w61_6_c0 :  std_logic;
signal bh7_w62_5_c0 :  std_logic;
signal bh7_w63_6_c0 :  std_logic;
signal tile_25_X_c0 :  std_logic_vector(3 downto 0);
signal tile_25_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_25_output_c0 :  std_logic_vector(3 downto 0);
signal tile_25_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w56_5_c0 :  std_logic;
signal bh7_w57_6_c0 :  std_logic;
signal bh7_w58_6_c0 :  std_logic;
signal bh7_w59_5_c0 :  std_logic;
signal tile_26_X_c0 :  std_logic_vector(3 downto 0);
signal tile_26_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_26_output_c0 :  std_logic_vector(3 downto 0);
signal tile_26_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w52_5_c0 :  std_logic;
signal bh7_w53_5_c0 :  std_logic;
signal bh7_w54_6_c0 :  std_logic;
signal bh7_w55_6_c0 :  std_logic;
signal tile_27_X_c0 :  std_logic_vector(1 downto 0);
signal tile_27_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_27_output_c0 :  std_logic_vector(3 downto 0);
signal tile_27_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w65_5_c0 :  std_logic;
signal bh7_w66_6_c0 :  std_logic;
signal bh7_w67_6_c0 :  std_logic;
signal bh7_w68_5_c0 :  std_logic;
signal tile_28_X_c0 :  std_logic_vector(2 downto 0);
signal tile_28_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_28_output_c0 :  std_logic_vector(4 downto 0);
signal tile_28_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w62_6_c0 :  std_logic;
signal bh7_w63_7_c0 :  std_logic;
signal bh7_w64_7_c0 :  std_logic;
signal bh7_w65_6_c0 :  std_logic;
signal bh7_w66_7_c0 :  std_logic;
signal tile_29_X_c0 :  std_logic_vector(2 downto 0);
signal tile_29_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_29_output_c0 :  std_logic_vector(4 downto 0);
signal tile_29_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w59_6_c0 :  std_logic;
signal bh7_w60_7_c0 :  std_logic;
signal bh7_w61_7_c0 :  std_logic;
signal bh7_w62_7_c0 :  std_logic;
signal bh7_w63_8_c0 :  std_logic;
signal tile_30_X_c0 :  std_logic_vector(2 downto 0);
signal tile_30_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_30_output_c0 :  std_logic_vector(4 downto 0);
signal tile_30_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w56_6_c0 :  std_logic;
signal bh7_w57_7_c0 :  std_logic;
signal bh7_w58_7_c0 :  std_logic;
signal bh7_w59_7_c0 :  std_logic;
signal bh7_w60_8_c0 :  std_logic;
signal tile_31_X_c0 :  std_logic_vector(2 downto 0);
signal tile_31_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_31_output_c0 :  std_logic_vector(4 downto 0);
signal tile_31_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w53_6_c0 :  std_logic;
signal bh7_w54_7_c0 :  std_logic;
signal bh7_w55_7_c0 :  std_logic;
signal bh7_w56_7_c0 :  std_logic;
signal bh7_w57_8_c0 :  std_logic;
signal tile_32_X_c0 :  std_logic_vector(2 downto 0);
signal tile_32_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_32_output_c0 :  std_logic_vector(4 downto 0);
signal tile_32_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w50_4_c0 :  std_logic;
signal bh7_w51_5_c0 :  std_logic;
signal bh7_w52_6_c0 :  std_logic;
signal bh7_w53_7_c0 :  std_logic;
signal bh7_w54_8_c0 :  std_logic;
signal tile_33_X_c0 :  std_logic_vector(1 downto 0);
signal tile_33_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_33_output_c0 :  std_logic_vector(3 downto 0);
signal tile_33_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w63_9_c0 :  std_logic;
signal bh7_w64_8_c0 :  std_logic;
signal bh7_w65_7_c0 :  std_logic;
signal bh7_w66_8_c0 :  std_logic;
signal tile_34_X_c0 :  std_logic_vector(2 downto 0);
signal tile_34_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_34_output_c0 :  std_logic_vector(4 downto 0);
signal tile_34_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w60_9_c0 :  std_logic;
signal bh7_w61_8_c0 :  std_logic;
signal bh7_w62_8_c0 :  std_logic;
signal bh7_w63_10_c0 :  std_logic;
signal bh7_w64_9_c0 :  std_logic;
signal tile_35_X_c0 :  std_logic_vector(2 downto 0);
signal tile_35_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_35_output_c0 :  std_logic_vector(4 downto 0);
signal tile_35_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w57_9_c0 :  std_logic;
signal bh7_w58_8_c0 :  std_logic;
signal bh7_w59_8_c0 :  std_logic;
signal bh7_w60_10_c0 :  std_logic;
signal bh7_w61_9_c0 :  std_logic;
signal tile_36_X_c0 :  std_logic_vector(2 downto 0);
signal tile_36_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_36_output_c0 :  std_logic_vector(4 downto 0);
signal tile_36_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w54_9_c0 :  std_logic;
signal bh7_w55_8_c0 :  std_logic;
signal bh7_w56_8_c0 :  std_logic;
signal bh7_w57_10_c0 :  std_logic;
signal bh7_w58_9_c0 :  std_logic;
signal tile_37_X_c0 :  std_logic_vector(2 downto 0);
signal tile_37_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_37_output_c0 :  std_logic_vector(4 downto 0);
signal tile_37_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w51_6_c0 :  std_logic;
signal bh7_w52_7_c0 :  std_logic;
signal bh7_w53_8_c0 :  std_logic;
signal bh7_w54_10_c0 :  std_logic;
signal bh7_w55_9_c0 :  std_logic;
signal tile_38_X_c0 :  std_logic_vector(2 downto 0);
signal tile_38_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_38_output_c0 :  std_logic_vector(4 downto 0);
signal tile_38_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w48_4_c0 :  std_logic;
signal bh7_w49_4_c0 :  std_logic;
signal bh7_w50_5_c0 :  std_logic;
signal bh7_w51_7_c0 :  std_logic;
signal bh7_w52_8_c0 :  std_logic;
signal tile_39_X_c0 :  std_logic_vector(0 downto 0);
signal tile_39_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_39_output_c0 :  std_logic_vector(0 downto 0);
signal tile_39_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w85_3_c0 :  std_logic;
signal tile_40_X_c0 :  std_logic_vector(3 downto 0);
signal tile_40_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_40_output_c0 :  std_logic_vector(3 downto 0);
signal tile_40_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w81_4_c0 :  std_logic;
signal bh7_w82_3_c0 :  std_logic;
signal bh7_w83_2_c0 :  std_logic;
signal bh7_w84_3_c0 :  std_logic;
signal tile_41_X_c0 :  std_logic_vector(3 downto 0);
signal tile_41_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_41_output_c0 :  std_logic_vector(3 downto 0);
signal tile_41_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w77_3_c0 :  std_logic;
signal bh7_w78_4_c0 :  std_logic;
signal bh7_w79_4_c0 :  std_logic;
signal bh7_w80_3_c0 :  std_logic;
signal tile_42_X_c0 :  std_logic_vector(3 downto 0);
signal tile_42_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_42_output_c0 :  std_logic_vector(3 downto 0);
signal tile_42_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w73_5_c0 :  std_logic;
signal bh7_w74_4_c0 :  std_logic;
signal bh7_w75_4_c0 :  std_logic;
signal bh7_w76_4_c0 :  std_logic;
signal tile_43_X_c0 :  std_logic_vector(3 downto 0);
signal tile_43_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_43_output_c0 :  std_logic_vector(3 downto 0);
signal tile_43_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w69_5_c0 :  std_logic;
signal bh7_w70_5_c0 :  std_logic;
signal bh7_w71_4_c0 :  std_logic;
signal bh7_w72_5_c0 :  std_logic;
signal tile_44_X_c0 :  std_logic_vector(1 downto 0);
signal tile_44_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_44_output_c0 :  std_logic_vector(3 downto 0);
signal tile_44_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w82_4_c0 :  std_logic;
signal bh7_w83_3_c0 :  std_logic;
signal bh7_w84_4_c0 :  std_logic;
signal bh7_w85_4_c0 :  std_logic;
signal tile_45_X_c0 :  std_logic_vector(2 downto 0);
signal tile_45_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_45_output_c0 :  std_logic_vector(4 downto 0);
signal tile_45_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w79_5_c0 :  std_logic;
signal bh7_w80_4_c0 :  std_logic;
signal bh7_w81_5_c0 :  std_logic;
signal bh7_w82_5_c0 :  std_logic;
signal bh7_w83_4_c0 :  std_logic;
signal tile_46_X_c0 :  std_logic_vector(2 downto 0);
signal tile_46_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_46_output_c0 :  std_logic_vector(4 downto 0);
signal tile_46_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w76_5_c0 :  std_logic;
signal bh7_w77_4_c0 :  std_logic;
signal bh7_w78_5_c0 :  std_logic;
signal bh7_w79_6_c0 :  std_logic;
signal bh7_w80_5_c0 :  std_logic;
signal tile_47_X_c0 :  std_logic_vector(2 downto 0);
signal tile_47_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_47_output_c0 :  std_logic_vector(4 downto 0);
signal tile_47_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w73_6_c0 :  std_logic;
signal bh7_w74_5_c0 :  std_logic;
signal bh7_w75_5_c0 :  std_logic;
signal bh7_w76_6_c0 :  std_logic;
signal bh7_w77_5_c0 :  std_logic;
signal tile_48_X_c0 :  std_logic_vector(2 downto 0);
signal tile_48_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_48_output_c0 :  std_logic_vector(4 downto 0);
signal tile_48_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w70_6_c0 :  std_logic;
signal bh7_w71_5_c0 :  std_logic;
signal bh7_w72_6_c0 :  std_logic;
signal bh7_w73_7_c0 :  std_logic;
signal bh7_w74_6_c0 :  std_logic;
signal tile_49_X_c0 :  std_logic_vector(2 downto 0);
signal tile_49_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_49_output_c0 :  std_logic_vector(4 downto 0);
signal tile_49_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w67_7_c0 :  std_logic;
signal bh7_w68_6_c0 :  std_logic;
signal bh7_w69_6_c0 :  std_logic;
signal bh7_w70_7_c0 :  std_logic;
signal bh7_w71_6_c0 :  std_logic;
signal tile_50_X_c0 :  std_logic_vector(1 downto 0);
signal tile_50_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_50_output_c0 :  std_logic_vector(3 downto 0);
signal tile_50_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w80_6_c0 :  std_logic;
signal bh7_w81_6_c0 :  std_logic;
signal bh7_w82_6_c0 :  std_logic;
signal bh7_w83_5_c0 :  std_logic;
signal tile_51_X_c0 :  std_logic_vector(2 downto 0);
signal tile_51_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_51_output_c0 :  std_logic_vector(4 downto 0);
signal tile_51_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w77_6_c0 :  std_logic;
signal bh7_w78_6_c0 :  std_logic;
signal bh7_w79_7_c0 :  std_logic;
signal bh7_w80_7_c0 :  std_logic;
signal bh7_w81_7_c0 :  std_logic;
signal tile_52_X_c0 :  std_logic_vector(2 downto 0);
signal tile_52_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_52_output_c0 :  std_logic_vector(4 downto 0);
signal tile_52_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w74_7_c0 :  std_logic;
signal bh7_w75_6_c0 :  std_logic;
signal bh7_w76_7_c0 :  std_logic;
signal bh7_w77_7_c0 :  std_logic;
signal bh7_w78_7_c0 :  std_logic;
signal tile_53_X_c0 :  std_logic_vector(2 downto 0);
signal tile_53_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_53_output_c0 :  std_logic_vector(4 downto 0);
signal tile_53_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w71_7_c0 :  std_logic;
signal bh7_w72_7_c0 :  std_logic;
signal bh7_w73_8_c0 :  std_logic;
signal bh7_w74_8_c0 :  std_logic;
signal bh7_w75_7_c0 :  std_logic;
signal tile_54_X_c0 :  std_logic_vector(2 downto 0);
signal tile_54_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_54_output_c0 :  std_logic_vector(4 downto 0);
signal tile_54_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w68_7_c0 :  std_logic;
signal bh7_w69_7_c0 :  std_logic;
signal bh7_w70_8_c0 :  std_logic;
signal bh7_w71_8_c0 :  std_logic;
signal bh7_w72_8_c0 :  std_logic;
signal tile_55_X_c0 :  std_logic_vector(2 downto 0);
signal tile_55_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_55_output_c0 :  std_logic_vector(4 downto 0);
signal tile_55_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w65_8_c0 :  std_logic;
signal bh7_w66_9_c0 :  std_logic;
signal bh7_w67_8_c0 :  std_logic;
signal bh7_w68_8_c0 :  std_logic;
signal bh7_w69_8_c0 :  std_logic;
signal tile_56_X_c0 :  std_logic_vector(0 downto 0);
signal tile_56_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_56_output_c0 :  std_logic_vector(0 downto 0);
signal tile_56_filtered_output_c0 :  unsigned(0-0 downto 0);
signal bh7_w102_0_c0 :  std_logic;
signal tile_57_X_c0 :  std_logic_vector(3 downto 0);
signal tile_57_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_57_output_c0 :  std_logic_vector(3 downto 0);
signal tile_57_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w98_2_c0 :  std_logic;
signal bh7_w99_1_c0 :  std_logic;
signal bh7_w100_1_c0 :  std_logic;
signal bh7_w101_0_c0 :  std_logic;
signal tile_58_X_c0 :  std_logic_vector(3 downto 0);
signal tile_58_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_58_output_c0 :  std_logic_vector(3 downto 0);
signal tile_58_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w94_3_c0 :  std_logic;
signal bh7_w95_2_c0 :  std_logic;
signal bh7_w96_3_c0 :  std_logic;
signal bh7_w97_3_c0 :  std_logic;
signal tile_59_X_c0 :  std_logic_vector(3 downto 0);
signal tile_59_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_59_output_c0 :  std_logic_vector(3 downto 0);
signal tile_59_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w90_3_c0 :  std_logic;
signal bh7_w91_3_c0 :  std_logic;
signal bh7_w92_2_c0 :  std_logic;
signal bh7_w93_3_c0 :  std_logic;
signal tile_60_X_c0 :  std_logic_vector(3 downto 0);
signal tile_60_Y_c0 :  std_logic_vector(0 downto 0);
signal tile_60_output_c0 :  std_logic_vector(3 downto 0);
signal tile_60_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w86_2_c0 :  std_logic;
signal bh7_w87_3_c0 :  std_logic;
signal bh7_w88_3_c0 :  std_logic;
signal bh7_w89_2_c0 :  std_logic;
signal tile_61_X_c0 :  std_logic_vector(1 downto 0);
signal tile_61_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_61_output_c0 :  std_logic_vector(3 downto 0);
signal tile_61_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w99_2_c0 :  std_logic;
signal bh7_w100_2_c0 :  std_logic;
signal bh7_w101_1_c0 :  std_logic;
signal bh7_w102_1_c0 :  std_logic;
signal tile_62_X_c0 :  std_logic_vector(2 downto 0);
signal tile_62_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_62_output_c0 :  std_logic_vector(4 downto 0);
signal tile_62_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w96_4_c0 :  std_logic;
signal bh7_w97_4_c0 :  std_logic;
signal bh7_w98_3_c0 :  std_logic;
signal bh7_w99_3_c0 :  std_logic;
signal bh7_w100_3_c0 :  std_logic;
signal tile_63_X_c0 :  std_logic_vector(2 downto 0);
signal tile_63_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_63_output_c0 :  std_logic_vector(4 downto 0);
signal tile_63_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w93_4_c0 :  std_logic;
signal bh7_w94_4_c0 :  std_logic;
signal bh7_w95_3_c0 :  std_logic;
signal bh7_w96_5_c0 :  std_logic;
signal bh7_w97_5_c0 :  std_logic;
signal tile_64_X_c0 :  std_logic_vector(2 downto 0);
signal tile_64_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_64_output_c0 :  std_logic_vector(4 downto 0);
signal tile_64_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w90_4_c0 :  std_logic;
signal bh7_w91_4_c0 :  std_logic;
signal bh7_w92_3_c0 :  std_logic;
signal bh7_w93_5_c0 :  std_logic;
signal bh7_w94_5_c0 :  std_logic;
signal tile_65_X_c0 :  std_logic_vector(2 downto 0);
signal tile_65_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_65_output_c0 :  std_logic_vector(4 downto 0);
signal tile_65_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w87_4_c0 :  std_logic;
signal bh7_w88_4_c0 :  std_logic;
signal bh7_w89_3_c0 :  std_logic;
signal bh7_w90_5_c0 :  std_logic;
signal bh7_w91_5_c0 :  std_logic;
signal tile_66_X_c0 :  std_logic_vector(2 downto 0);
signal tile_66_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_66_output_c0 :  std_logic_vector(4 downto 0);
signal tile_66_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w84_5_c0 :  std_logic;
signal bh7_w85_5_c0 :  std_logic;
signal bh7_w86_3_c0 :  std_logic;
signal bh7_w87_5_c0 :  std_logic;
signal bh7_w88_5_c0 :  std_logic;
signal tile_67_X_c0 :  std_logic_vector(1 downto 0);
signal tile_67_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_67_output_c0 :  std_logic_vector(3 downto 0);
signal tile_67_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w97_6_c0 :  std_logic;
signal bh7_w98_4_c0 :  std_logic;
signal bh7_w99_4_c0 :  std_logic;
signal bh7_w100_4_c0 :  std_logic;
signal tile_68_X_c0 :  std_logic_vector(2 downto 0);
signal tile_68_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_68_output_c0 :  std_logic_vector(4 downto 0);
signal tile_68_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w94_6_c0 :  std_logic;
signal bh7_w95_4_c0 :  std_logic;
signal bh7_w96_6_c0 :  std_logic;
signal bh7_w97_7_c0 :  std_logic;
signal bh7_w98_5_c0 :  std_logic;
signal tile_69_X_c0 :  std_logic_vector(2 downto 0);
signal tile_69_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_69_output_c0 :  std_logic_vector(4 downto 0);
signal tile_69_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w91_6_c0 :  std_logic;
signal bh7_w92_4_c0 :  std_logic;
signal bh7_w93_6_c0 :  std_logic;
signal bh7_w94_7_c0 :  std_logic;
signal bh7_w95_5_c0 :  std_logic;
signal tile_70_X_c0 :  std_logic_vector(2 downto 0);
signal tile_70_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_70_output_c0 :  std_logic_vector(4 downto 0);
signal tile_70_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w88_6_c0 :  std_logic;
signal bh7_w89_4_c0 :  std_logic;
signal bh7_w90_6_c0 :  std_logic;
signal bh7_w91_7_c0 :  std_logic;
signal bh7_w92_5_c0 :  std_logic;
signal tile_71_X_c0 :  std_logic_vector(2 downto 0);
signal tile_71_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_71_output_c0 :  std_logic_vector(4 downto 0);
signal tile_71_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w85_6_c0 :  std_logic;
signal bh7_w86_4_c0 :  std_logic;
signal bh7_w87_6_c0 :  std_logic;
signal bh7_w88_7_c0 :  std_logic;
signal bh7_w89_5_c0 :  std_logic;
signal tile_72_X_c0 :  std_logic_vector(2 downto 0);
signal tile_72_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_72_output_c0 :  std_logic_vector(4 downto 0);
signal tile_72_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w82_7_c0 :  std_logic;
signal bh7_w83_6_c0 :  std_logic;
signal bh7_w84_6_c0 :  std_logic;
signal bh7_w85_7_c0 :  std_logic;
signal bh7_w86_5_c0 :  std_logic;
signal tile_73_X_c0 :  std_logic_vector(1 downto 0);
signal tile_73_Y_c0 :  std_logic_vector(1 downto 0);
signal tile_73_output_c0 :  std_logic_vector(3 downto 0);
signal tile_73_filtered_output_c0 :  unsigned(3-0 downto 0);
signal bh7_w102_2_c0 :  std_logic;
signal bh7_w103_0_c0 :  std_logic;
signal bh7_w104_0_c0 :  std_logic;
signal bh7_w105_0_c0 :  std_logic;
signal tile_74_X_c0 :  std_logic_vector(1 downto 0);
signal tile_74_Y_c0 :  std_logic_vector(2 downto 0);
signal tile_74_output_c0 :  std_logic_vector(4 downto 0);
signal tile_74_filtered_output_c0 :  unsigned(4-0 downto 0);
signal bh7_w99_5_c0 :  std_logic;
signal bh7_w100_5_c0 :  std_logic;
signal bh7_w101_2_c0 :  std_logic;
signal bh7_w102_3_c0 :  std_logic;
signal bh7_w103_1_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid323_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid323_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w49_5_c0 :  std_logic;
signal bh7_w50_6_c0 :  std_logic;
signal bh7_w51_8_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_copy324_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid327_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid327_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w51_9_c0 :  std_logic;
signal bh7_w52_9_c0 :  std_logic;
signal bh7_w53_9_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_copy328_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid329_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid329_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w52_10_c0 :  std_logic;
signal bh7_w53_10_c0 :  std_logic;
signal bh7_w54_11_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_copy330_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid331_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid331_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w53_11_c0 :  std_logic;
signal bh7_w54_12_c0 :  std_logic;
signal bh7_w55_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_copy332_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid335_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w54_13_c0 :  std_logic;
signal bh7_w55_11_c0 :  std_logic;
signal bh7_w56_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_copy336_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid337_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w55_12_c0 :  std_logic;
signal bh7_w56_10_c0 :  std_logic;
signal bh7_w57_11_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_copy338_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid339_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid339_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w56_11_c0 :  std_logic;
signal bh7_w57_12_c0 :  std_logic;
signal bh7_w58_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_copy340_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid341_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w57_13_c0 :  std_logic;
signal bh7_w58_11_c0 :  std_logic;
signal bh7_w59_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_copy342_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid343_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w58_12_c0 :  std_logic;
signal bh7_w59_10_c0 :  std_logic;
signal bh7_w60_11_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_copy344_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid345_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid345_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w59_11_c0 :  std_logic;
signal bh7_w60_12_c0 :  std_logic;
signal bh7_w61_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_copy346_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid347_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w60_13_c0 :  std_logic;
signal bh7_w61_11_c0 :  std_logic;
signal bh7_w62_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_copy348_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid349_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w61_12_c0 :  std_logic;
signal bh7_w62_10_c0 :  std_logic;
signal bh7_w63_11_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_copy350_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid351_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid351_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w62_11_c0 :  std_logic;
signal bh7_w63_12_c0 :  std_logic;
signal bh7_w64_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_copy352_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid353_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w63_13_c0 :  std_logic;
signal bh7_w64_11_c0 :  std_logic;
signal bh7_w65_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_copy354_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid355_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w64_12_c0 :  std_logic;
signal bh7_w65_10_c0 :  std_logic;
signal bh7_w66_10_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_copy356_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid357_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w65_11_c0 :  std_logic;
signal bh7_w66_11_c0 :  std_logic;
signal bh7_w67_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_copy358_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid359_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_12_c0 :  std_logic;
signal bh7_w67_10_c0 :  std_logic;
signal bh7_w68_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_copy360_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid361_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w67_11_c0 :  std_logic;
signal bh7_w68_10_c0 :  std_logic;
signal bh7_w69_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_copy362_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid363_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_11_c0 :  std_logic;
signal bh7_w69_10_c0 :  std_logic;
signal bh7_w70_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_copy364_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid365_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w69_11_c0 :  std_logic;
signal bh7_w70_10_c0 :  std_logic;
signal bh7_w71_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_copy366_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid367_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_11_c0 :  std_logic;
signal bh7_w71_10_c0 :  std_logic;
signal bh7_w72_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_copy368_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid369_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w71_11_c0 :  std_logic;
signal bh7_w72_10_c0 :  std_logic;
signal bh7_w73_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_copy370_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid371_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_11_c0 :  std_logic;
signal bh7_w73_10_c0 :  std_logic;
signal bh7_w74_9_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_copy372_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid373_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w73_11_c0 :  std_logic;
signal bh7_w74_10_c0 :  std_logic;
signal bh7_w75_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_copy374_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid375_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_11_c0 :  std_logic;
signal bh7_w75_9_c0 :  std_logic;
signal bh7_w76_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_copy376_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid377_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w75_10_c0 :  std_logic;
signal bh7_w76_9_c0 :  std_logic;
signal bh7_w77_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_copy378_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid379_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_10_c0 :  std_logic;
signal bh7_w77_9_c0 :  std_logic;
signal bh7_w78_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_copy380_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid381_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w77_10_c0 :  std_logic;
signal bh7_w78_9_c0 :  std_logic;
signal bh7_w79_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_copy382_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid383_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_10_c0 :  std_logic;
signal bh7_w79_9_c0 :  std_logic;
signal bh7_w80_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_copy384_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid385_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w79_10_c0 :  std_logic;
signal bh7_w80_9_c0 :  std_logic;
signal bh7_w81_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_copy386_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid387_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_10_c0 :  std_logic;
signal bh7_w81_9_c0 :  std_logic;
signal bh7_w82_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_copy388_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid389_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w81_10_c0 :  std_logic;
signal bh7_w82_9_c0 :  std_logic;
signal bh7_w83_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_copy390_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid391_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_10_c0 :  std_logic;
signal bh7_w83_8_c0 :  std_logic;
signal bh7_w84_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_copy392_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid393_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w83_9_c0 :  std_logic;
signal bh7_w84_8_c0 :  std_logic;
signal bh7_w85_8_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_copy394_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid395_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w84_9_c0 :  std_logic;
signal bh7_w85_9_c0 :  std_logic;
signal bh7_w86_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_copy396_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid397_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w85_10_c0 :  std_logic;
signal bh7_w86_7_c0 :  std_logic;
signal bh7_w87_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_copy398_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid401_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w86_8_c0 :  std_logic;
signal bh7_w87_8_c0 :  std_logic;
signal bh7_w88_8_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_copy402_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid403_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w87_9_c0 :  std_logic;
signal bh7_w88_9_c0 :  std_logic;
signal bh7_w89_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_copy404_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid405_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w88_10_c0 :  std_logic;
signal bh7_w89_7_c0 :  std_logic;
signal bh7_w90_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_copy406_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid407_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w89_8_c0 :  std_logic;
signal bh7_w90_8_c0 :  std_logic;
signal bh7_w91_8_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_copy408_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid409_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w90_9_c0 :  std_logic;
signal bh7_w91_9_c0 :  std_logic;
signal bh7_w92_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_copy410_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid411_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w91_10_c0 :  std_logic;
signal bh7_w92_7_c0 :  std_logic;
signal bh7_w93_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_copy412_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid413_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w92_8_c0 :  std_logic;
signal bh7_w93_8_c0 :  std_logic;
signal bh7_w94_8_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_copy414_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid415_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w93_9_c0 :  std_logic;
signal bh7_w94_9_c0 :  std_logic;
signal bh7_w95_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_copy416_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid417_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w94_10_c0 :  std_logic;
signal bh7_w95_7_c0 :  std_logic;
signal bh7_w96_7_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_copy418_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid419_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w95_8_c0 :  std_logic;
signal bh7_w96_8_c0 :  std_logic;
signal bh7_w97_8_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_copy420_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid421_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w96_9_c0 :  std_logic;
signal bh7_w97_9_c0 :  std_logic;
signal bh7_w98_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_copy422_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid423_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w97_10_c0 :  std_logic;
signal bh7_w98_7_c0 :  std_logic;
signal bh7_w99_6_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_copy424_c0 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid425_In0_c0 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w98_8_c0 :  std_logic;
signal bh7_w99_7_c0 :  std_logic;
signal bh7_w100_6_c0 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_copy426_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid427_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w99_8_c0 :  std_logic;
signal bh7_w100_7_c0 :  std_logic;
signal bh7_w101_3_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_copy428_c0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid429_In0_c0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w100_8_c0 :  std_logic;
signal bh7_w101_4_c0 :  std_logic;
signal bh7_w102_4_c0 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_copy430_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid433_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w101_5_c0 :  std_logic;
signal bh7_w102_5_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_copy434_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid435_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid435_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w102_6_c0 :  std_logic;
signal bh7_w103_2_c0 :  std_logic;
signal bh7_w104_1_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_copy436_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid437_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid437_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w51_10_c0 :  std_logic;
signal bh7_w52_11_c0 :  std_logic;
signal bh7_w53_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_copy438_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid439_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid439_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w53_13_c0 :  std_logic;
signal bh7_w54_14_c0 :  std_logic;
signal bh7_w55_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_copy440_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid441_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w55_14_c0 :  std_logic;
signal bh7_w56_12_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_copy442_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid443_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid443_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w56_13_c0 :  std_logic;
signal bh7_w57_14_c0 :  std_logic;
signal bh7_w58_13_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_copy444_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid445_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w57_15_c0 :  std_logic;
signal bh7_w58_14_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_copy446_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid447_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w58_15_c0 :  std_logic;
signal bh7_w59_12_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_copy448_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid449_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid449_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w59_13_c0 :  std_logic;
signal bh7_w60_14_c0 :  std_logic;
signal bh7_w61_13_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_copy450_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid451_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w60_15_c0 :  std_logic;
signal bh7_w61_14_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_copy452_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid453_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w61_15_c0 :  std_logic;
signal bh7_w62_12_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_copy454_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid455_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid455_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w62_13_c0 :  std_logic;
signal bh7_w63_14_c0 :  std_logic;
signal bh7_w64_13_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_copy456_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid457_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w63_15_c0 :  std_logic;
signal bh7_w64_14_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_copy458_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid459_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid459_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w64_15_c0 :  std_logic;
signal bh7_w65_12_c0 :  std_logic;
signal bh7_w66_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_copy460_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid461_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid461_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_14_c0 :  std_logic;
signal bh7_w67_12_c0 :  std_logic;
signal bh7_w68_12_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_copy462_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid463_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w67_13_c0 :  std_logic;
signal bh7_w68_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_copy464_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid465_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid465_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_14_c0 :  std_logic;
signal bh7_w69_12_c0 :  std_logic;
signal bh7_w70_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_copy466_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid467_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid467_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_13_c0 :  std_logic;
signal bh7_w71_12_c0 :  std_logic;
signal bh7_w72_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_copy468_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid469_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid469_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_13_c0 :  std_logic;
signal bh7_w73_12_c0 :  std_logic;
signal bh7_w74_12_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_copy470_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid471_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid471_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_13_c0 :  std_logic;
signal bh7_w75_11_c0 :  std_logic;
signal bh7_w76_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_copy472_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid473_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid473_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_12_c0 :  std_logic;
signal bh7_w77_11_c0 :  std_logic;
signal bh7_w78_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_copy474_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid475_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid475_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_12_c0 :  std_logic;
signal bh7_w79_11_c0 :  std_logic;
signal bh7_w80_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_copy476_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid477_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid477_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_12_c0 :  std_logic;
signal bh7_w81_11_c0 :  std_logic;
signal bh7_w82_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_copy478_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid479_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid479_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_12_c0 :  std_logic;
signal bh7_w83_10_c0 :  std_logic;
signal bh7_w84_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_copy480_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid481_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w83_11_c0 :  std_logic;
signal bh7_w84_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_copy482_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid483_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w84_12_c0 :  std_logic;
signal bh7_w85_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_copy484_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid485_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid485_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w85_12_c0 :  std_logic;
signal bh7_w86_9_c0 :  std_logic;
signal bh7_w87_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_copy486_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid487_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w86_10_c0 :  std_logic;
signal bh7_w87_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_copy488_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid489_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w87_12_c0 :  std_logic;
signal bh7_w88_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_copy490_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid491_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid491_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w88_12_c0 :  std_logic;
signal bh7_w89_9_c0 :  std_logic;
signal bh7_w90_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_copy492_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid493_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w89_10_c0 :  std_logic;
signal bh7_w90_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_copy494_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid495_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w90_12_c0 :  std_logic;
signal bh7_w91_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_copy496_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid497_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid497_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w91_12_c0 :  std_logic;
signal bh7_w92_9_c0 :  std_logic;
signal bh7_w93_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_copy498_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid499_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w92_10_c0 :  std_logic;
signal bh7_w93_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_copy500_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid501_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w93_12_c0 :  std_logic;
signal bh7_w94_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_copy502_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid503_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid503_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w94_12_c0 :  std_logic;
signal bh7_w95_9_c0 :  std_logic;
signal bh7_w96_10_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_copy504_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid505_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w95_10_c0 :  std_logic;
signal bh7_w96_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_copy506_c0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid507_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w96_12_c0 :  std_logic;
signal bh7_w97_11_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_copy508_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid509_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid509_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w97_12_c0 :  std_logic;
signal bh7_w98_9_c0 :  std_logic;
signal bh7_w99_9_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_copy510_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid511_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w98_10_c0 :  std_logic;
signal bh7_w99_10_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_copy512_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid513_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid513_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w99_11_c0 :  std_logic;
signal bh7_w100_9_c0 :  std_logic;
signal bh7_w101_6_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_copy514_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid515_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid515_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w101_7_c0 :  std_logic;
signal bh7_w102_7_c0 :  std_logic;
signal bh7_w103_3_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_copy516_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid517_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid517_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w103_4_c0 :  std_logic;
signal bh7_w104_2_c0 :  std_logic;
signal bh7_w105_1_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_copy518_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid519_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid519_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w53_14_c0 :  std_logic;
signal bh7_w54_15_c0 :  std_logic;
signal bh7_w55_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_copy520_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid521_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid521_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w55_16_c0 :  std_logic;
signal bh7_w56_14_c0 :  std_logic;
signal bh7_w57_16_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_copy522_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid523_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w57_17_c0 :  std_logic;
signal bh7_w58_16_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_copy524_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid525_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid525_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w58_17_c0 :  std_logic;
signal bh7_w59_14_c0 :  std_logic;
signal bh7_w60_16_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_copy526_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid527_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w60_17_c0 :  std_logic;
signal bh7_w61_16_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_copy528_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid529_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid529_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w61_17_c0 :  std_logic;
signal bh7_w62_14_c0 :  std_logic;
signal bh7_w63_16_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_copy530_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid531_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w63_17_c0 :  std_logic;
signal bh7_w64_16_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_copy532_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid533_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid533_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w64_17_c0 :  std_logic;
signal bh7_w65_13_c0 :  std_logic;
signal bh7_w66_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_copy534_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid535_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid535_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_16_c0 :  std_logic;
signal bh7_w67_14_c0 :  std_logic;
signal bh7_w68_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_copy536_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid537_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid537_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_16_c0 :  std_logic;
signal bh7_w69_13_c0 :  std_logic;
signal bh7_w70_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_copy538_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid539_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid539_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_15_c0 :  std_logic;
signal bh7_w71_13_c0 :  std_logic;
signal bh7_w72_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_copy540_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid541_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid541_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_15_c0 :  std_logic;
signal bh7_w73_13_c0 :  std_logic;
signal bh7_w74_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_copy542_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid543_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid543_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_15_c0 :  std_logic;
signal bh7_w75_12_c0 :  std_logic;
signal bh7_w76_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_copy544_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid545_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid545_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_14_c0 :  std_logic;
signal bh7_w77_12_c0 :  std_logic;
signal bh7_w78_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_copy546_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid547_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid547_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_14_c0 :  std_logic;
signal bh7_w79_12_c0 :  std_logic;
signal bh7_w80_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_copy548_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid549_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid549_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_14_c0 :  std_logic;
signal bh7_w81_12_c0 :  std_logic;
signal bh7_w82_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_copy550_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid551_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid551_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_14_c0 :  std_logic;
signal bh7_w83_12_c0 :  std_logic;
signal bh7_w84_13_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_copy552_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid553_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid553_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w84_14_c0 :  std_logic;
signal bh7_w85_13_c0 :  std_logic;
signal bh7_w86_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_copy554_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid555_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w86_12_c0 :  std_logic;
signal bh7_w87_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_copy556_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid557_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid557_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w87_14_c0 :  std_logic;
signal bh7_w88_13_c0 :  std_logic;
signal bh7_w89_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_copy558_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid559_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w89_12_c0 :  std_logic;
signal bh7_w90_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_copy560_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid561_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid561_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w90_14_c0 :  std_logic;
signal bh7_w91_13_c0 :  std_logic;
signal bh7_w92_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_copy562_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid563_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w92_12_c0 :  std_logic;
signal bh7_w93_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_copy564_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid565_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid565_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w93_14_c0 :  std_logic;
signal bh7_w94_13_c0 :  std_logic;
signal bh7_w95_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_copy566_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid567_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w95_12_c0 :  std_logic;
signal bh7_w96_13_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_copy568_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid569_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid569_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w96_14_c0 :  std_logic;
signal bh7_w97_13_c0 :  std_logic;
signal bh7_w98_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_copy570_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid571_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w98_12_c0 :  std_logic;
signal bh7_w99_12_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_copy572_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid573_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid573_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w99_13_c0 :  std_logic;
signal bh7_w100_10_c0 :  std_logic;
signal bh7_w101_8_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_copy574_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid575_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid575_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w101_9_c0 :  std_logic;
signal bh7_w102_8_c0 :  std_logic;
signal bh7_w103_5_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_copy576_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid577_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid577_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w103_6_c0 :  std_logic;
signal bh7_w104_3_c0 :  std_logic;
signal bh7_w105_2_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_copy578_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid579_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_c0 :  std_logic_vector(1 downto 0);
signal bh7_w105_3_c0 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_copy580_c0 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid581_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid581_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w55_17_c0 :  std_logic;
signal bh7_w56_15_c0 :  std_logic;
signal bh7_w57_18_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_copy582_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid583_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid583_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w57_19_c0 :  std_logic;
signal bh7_w58_18_c0 :  std_logic;
signal bh7_w59_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_copy584_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid585_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid585_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w60_18_c0 :  std_logic;
signal bh7_w61_18_c0, bh7_w61_18_c1 :  std_logic;
signal bh7_w62_15_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_copy586_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid587_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid587_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w63_18_c0 :  std_logic;
signal bh7_w64_18_c0, bh7_w64_18_c1 :  std_logic;
signal bh7_w65_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_copy588_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid589_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid589_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w66_17_c0 :  std_logic;
signal bh7_w67_15_c0, bh7_w67_15_c1 :  std_logic;
signal bh7_w68_17_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_copy590_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid591_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid591_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w68_18_c0 :  std_logic;
signal bh7_w69_14_c0 :  std_logic;
signal bh7_w70_16_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_copy592_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid593_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid593_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w70_17_c0 :  std_logic;
signal bh7_w71_14_c0 :  std_logic;
signal bh7_w72_16_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_copy594_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid595_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid595_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w72_17_c0 :  std_logic;
signal bh7_w73_14_c0 :  std_logic;
signal bh7_w74_16_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_copy596_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid597_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid597_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w74_17_c0 :  std_logic;
signal bh7_w75_13_c0 :  std_logic;
signal bh7_w76_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_copy598_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid599_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid599_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w76_16_c0 :  std_logic;
signal bh7_w77_13_c0 :  std_logic;
signal bh7_w78_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_copy600_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid601_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid601_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w78_16_c0 :  std_logic;
signal bh7_w79_13_c0 :  std_logic;
signal bh7_w80_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_copy602_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid603_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid603_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w80_16_c0 :  std_logic;
signal bh7_w81_13_c0 :  std_logic;
signal bh7_w82_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_copy604_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid605_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid605_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w82_16_c0 :  std_logic;
signal bh7_w83_13_c0 :  std_logic;
signal bh7_w84_15_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_copy606_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid607_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid607_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w84_16_c0 :  std_logic;
signal bh7_w85_14_c0 :  std_logic;
signal bh7_w86_13_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_copy608_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid609_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid609_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w86_14_c0 :  std_logic;
signal bh7_w87_15_c0 :  std_logic;
signal bh7_w88_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_copy610_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid611_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid611_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w89_13_c0 :  std_logic;
signal bh7_w90_15_c0, bh7_w90_15_c1 :  std_logic;
signal bh7_w91_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_copy612_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid613_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid613_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w92_13_c0 :  std_logic;
signal bh7_w93_15_c0, bh7_w93_15_c1 :  std_logic;
signal bh7_w94_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_copy614_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid615_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid615_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w95_13_c0 :  std_logic;
signal bh7_w96_15_c0, bh7_w96_15_c1 :  std_logic;
signal bh7_w97_14_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_copy616_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid617_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid617_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w98_13_c0 :  std_logic;
signal bh7_w99_14_c0, bh7_w99_14_c1 :  std_logic;
signal bh7_w100_11_c0 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_copy618_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid619_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid619_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w101_10_c0 :  std_logic;
signal bh7_w102_9_c0, bh7_w102_9_c1 :  std_logic;
signal bh7_w103_7_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_copy620_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid621_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid621_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w103_8_c0 :  std_logic;
signal bh7_w104_4_c0 :  std_logic;
signal bh7_w105_4_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_copy622_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid623_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid623_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_c0 :  std_logic_vector(2 downto 0);
signal bh7_w105_5_c0 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_copy624_c0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid625_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid625_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w57_20_c1 :  std_logic;
signal bh7_w58_19_c1 :  std_logic;
signal bh7_w59_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c0, Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid627_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid627_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_17_c1 :  std_logic;
signal bh7_w60_19_c1 :  std_logic;
signal bh7_w61_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c0, Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid629_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid629_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_16_c1 :  std_logic;
signal bh7_w63_19_c1 :  std_logic;
signal bh7_w64_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c0, Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid631_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid631_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w65_15_c1 :  std_logic;
signal bh7_w66_18_c1 :  std_logic;
signal bh7_w67_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c0, Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid633_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid633_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_19_c1 :  std_logic;
signal bh7_w69_15_c1 :  std_logic;
signal bh7_w70_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c0, Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid635_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid635_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_19_c1 :  std_logic;
signal bh7_w71_15_c1 :  std_logic;
signal bh7_w72_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c0, Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid637_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid637_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_19_c1 :  std_logic;
signal bh7_w73_15_c1 :  std_logic;
signal bh7_w74_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c0, Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid639_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid639_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_19_c1 :  std_logic;
signal bh7_w75_14_c1 :  std_logic;
signal bh7_w76_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c0, Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid641_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid641_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_18_c1 :  std_logic;
signal bh7_w77_14_c1 :  std_logic;
signal bh7_w78_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c0, Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid643_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid643_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_18_c1 :  std_logic;
signal bh7_w79_14_c1 :  std_logic;
signal bh7_w80_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c0, Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid645_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid645_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_18_c1 :  std_logic;
signal bh7_w81_14_c1 :  std_logic;
signal bh7_w82_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c0, Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid647_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid647_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_18_c1 :  std_logic;
signal bh7_w83_14_c1 :  std_logic;
signal bh7_w84_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c0, Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid649_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid649_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_18_c1 :  std_logic;
signal bh7_w85_15_c1 :  std_logic;
signal bh7_w86_15_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c0, Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid651_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid651_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_16_c1 :  std_logic;
signal bh7_w87_16_c1 :  std_logic;
signal bh7_w88_15_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c0, Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid653_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid653_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_16_c1 :  std_logic;
signal bh7_w89_14_c1 :  std_logic;
signal bh7_w90_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c0, Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid655_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid655_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w91_15_c1 :  std_logic;
signal bh7_w92_14_c1 :  std_logic;
signal bh7_w93_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c0, Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid657_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid657_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w94_15_c1 :  std_logic;
signal bh7_w95_14_c1 :  std_logic;
signal bh7_w96_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c0, Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid659_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid659_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w97_15_c1 :  std_logic;
signal bh7_w98_14_c1 :  std_logic;
signal bh7_w99_15_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c0, Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid661_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid661_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w100_12_c1 :  std_logic;
signal bh7_w101_11_c1 :  std_logic;
signal bh7_w102_10_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c0, Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid663_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid663_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w103_9_c1 :  std_logic;
signal bh7_w104_5_c1 :  std_logic;
signal bh7_w105_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c0, Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid665_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid665_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w105_7_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c0, Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid667_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid667_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w17_2_c1 :  std_logic;
signal bh7_w18_2_c1 :  std_logic;
signal bh7_w19_2_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c0, Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid669_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid669_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w19_3_c1 :  std_logic;
signal bh7_w20_2_c1 :  std_logic;
signal bh7_w21_2_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c0, Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid671_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid671_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_3_c1 :  std_logic;
signal bh7_w22_2_c1 :  std_logic;
signal bh7_w23_2_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c0, Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid673_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w23_3_c1 :  std_logic;
signal bh7_w24_3_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c0, Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid675_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid675_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w24_4_c1 :  std_logic;
signal bh7_w25_3_c1 :  std_logic;
signal bh7_w26_3_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c0, Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid677_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid677_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w26_4_c1 :  std_logic;
signal bh7_w27_3_c1 :  std_logic;
signal bh7_w28_3_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c0, Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid679_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid679_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w28_4_c1 :  std_logic;
signal bh7_w29_3_c1 :  std_logic;
signal bh7_w30_3_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c0, Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid681_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid681_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w30_4_c1 :  std_logic;
signal bh7_w31_3_c1 :  std_logic;
signal bh7_w32_3_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c0, Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid683_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid683_In1_c0 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w32_4_c1 :  std_logic;
signal bh7_w33_3_c1 :  std_logic;
signal bh7_w34_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c0, Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid685_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid685_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w34_5_c1 :  std_logic;
signal bh7_w35_4_c1 :  std_logic;
signal bh7_w36_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c0, Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid687_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w35_5_c1 :  std_logic;
signal bh7_w36_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c0, Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid689_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid689_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w36_6_c1 :  std_logic;
signal bh7_w37_4_c1 :  std_logic;
signal bh7_w38_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c0, Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid691_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w37_5_c1 :  std_logic;
signal bh7_w38_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c0, Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid693_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid693_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w38_6_c1 :  std_logic;
signal bh7_w39_4_c1 :  std_logic;
signal bh7_w40_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c0, Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid695_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w39_5_c1 :  std_logic;
signal bh7_w40_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c0, Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid697_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid697_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w40_6_c1 :  std_logic;
signal bh7_w41_4_c1 :  std_logic;
signal bh7_w42_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c0, Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid699_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w41_5_c1 :  std_logic;
signal bh7_w42_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c0, Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid701_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid701_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w42_6_c1 :  std_logic;
signal bh7_w43_4_c1 :  std_logic;
signal bh7_w44_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c0, Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid703_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w43_5_c1 :  std_logic;
signal bh7_w44_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c0, Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid705_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid705_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w44_6_c1 :  std_logic;
signal bh7_w45_4_c1 :  std_logic;
signal bh7_w46_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c0, Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid707_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w45_5_c1 :  std_logic;
signal bh7_w46_5_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c0, Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid709_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid709_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w46_6_c1 :  std_logic;
signal bh7_w47_4_c1 :  std_logic;
signal bh7_w48_5_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c0, Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid711_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w47_5_c1 :  std_logic;
signal bh7_w48_6_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c0, Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid713_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid713_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w48_7_c1 :  std_logic;
signal bh7_w49_6_c1 :  std_logic;
signal bh7_w50_7_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c0, Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid715_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid715_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w49_7_c1 :  std_logic;
signal bh7_w50_8_c1 :  std_logic;
signal bh7_w51_11_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c0, Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid717_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid717_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w50_9_c1 :  std_logic;
signal bh7_w51_12_c1 :  std_logic;
signal bh7_w52_12_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c0, Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid719_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid719_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w51_13_c1 :  std_logic;
signal bh7_w52_13_c1 :  std_logic;
signal bh7_w53_15_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c0, Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid721_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid721_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w52_14_c1 :  std_logic;
signal bh7_w53_16_c1 :  std_logic;
signal bh7_w54_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c0, Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid723_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid723_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w53_17_c1 :  std_logic;
signal bh7_w54_17_c1 :  std_logic;
signal bh7_w55_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c0, Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid725_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid725_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w54_18_c1 :  std_logic;
signal bh7_w55_19_c1 :  std_logic;
signal bh7_w56_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c0, Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid727_In0_c0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid727_In1_c0 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w55_20_c1 :  std_logic;
signal bh7_w56_17_c1 :  std_logic;
signal bh7_w57_21_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c0, Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c0, Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid729_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_18_c1 :  std_logic;
signal bh7_w57_22_c1 :  std_logic;
signal bh7_w58_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_copy730_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c0, Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid731_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w57_23_c1 :  std_logic;
signal bh7_w58_21_c1 :  std_logic;
signal bh7_w59_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_copy732_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid733_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w58_22_c1 :  std_logic;
signal bh7_w59_19_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c0, Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c1 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid735_In0_c1 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_20_c1 :  std_logic;
signal bh7_w60_20_c1 :  std_logic;
signal bh7_w61_20_c1 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_copy736_c1 :  std_logic_vector(2 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid737_In0_c1 :  std_logic_vector(4 downto 0);
signal Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w60_21_c1 :  std_logic;
signal bh7_w61_21_c1 :  std_logic;
signal bh7_w62_17_c1 :  std_logic;
signal Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_copy738_c1 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid739_In0_c1 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w61_22_c1 :  std_logic;
signal bh7_w62_18_c1 :  std_logic;
signal bh7_w63_20_c1 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_copy740_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid741_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid741_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_19_c1 :  std_logic;
signal bh7_w63_21_c1 :  std_logic;
signal bh7_w64_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_copy742_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid743_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w63_22_c1 :  std_logic;
signal bh7_w64_21_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c0, Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c1 :  std_logic_vector(1 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid745_In0_c1 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_22_c1 :  std_logic;
signal bh7_w65_16_c1 :  std_logic;
signal bh7_w66_19_c1 :  std_logic;
signal Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_copy746_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid747_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid747_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w65_17_c1 :  std_logic;
signal bh7_w66_20_c1 :  std_logic;
signal bh7_w67_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_copy748_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid749_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w66_21_c1 :  std_logic;
signal bh7_w67_18_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c0, Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid751_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid751_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w67_19_c1 :  std_logic;
signal bh7_w68_20_c1 :  std_logic;
signal bh7_w69_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_copy752_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid753_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w68_21_c1 :  std_logic;
signal bh7_w69_17_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c0, Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid755_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid755_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w69_18_c1 :  std_logic;
signal bh7_w70_20_c1 :  std_logic;
signal bh7_w71_16_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_copy756_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid757_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid757_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w70_21_c1 :  std_logic;
signal bh7_w71_17_c1 :  std_logic;
signal bh7_w72_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_copy758_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid759_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w71_18_c1 :  std_logic;
signal bh7_w72_21_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c0, Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid761_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid761_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_22_c1 :  std_logic;
signal bh7_w73_16_c1 :  std_logic;
signal bh7_w74_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_copy762_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid763_In0_c0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w73_17_c1 :  std_logic;
signal bh7_w74_21_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c0, Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid765_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_22_c1 :  std_logic;
signal bh7_w75_15_c1 :  std_logic;
signal bh7_w76_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_copy766_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid767_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid767_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_23_c1 :  std_logic;
signal bh7_w75_16_c1 :  std_logic;
signal bh7_w76_20_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_copy768_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid769_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_21_c1 :  std_logic;
signal bh7_w77_15_c1 :  std_logic;
signal bh7_w78_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_copy770_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid771_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w77_16_c1 :  std_logic;
signal bh7_w78_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_copy772_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid773_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_21_c1 :  std_logic;
signal bh7_w79_15_c1 :  std_logic;
signal bh7_w80_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_copy774_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid775_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w79_16_c1 :  std_logic;
signal bh7_w80_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_copy776_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid777_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_21_c1 :  std_logic;
signal bh7_w81_15_c1 :  std_logic;
signal bh7_w82_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_copy778_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid779_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w81_16_c1 :  std_logic;
signal bh7_w82_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_copy780_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid781_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid781_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_21_c1 :  std_logic;
signal bh7_w83_15_c1 :  std_logic;
signal bh7_w84_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_copy782_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid783_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid783_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_20_c1 :  std_logic;
signal bh7_w85_16_c1 :  std_logic;
signal bh7_w86_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_copy784_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid785_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid785_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_18_c1 :  std_logic;
signal bh7_w87_17_c1 :  std_logic;
signal bh7_w88_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_copy786_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid787_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid787_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_18_c1 :  std_logic;
signal bh7_w89_15_c1 :  std_logic;
signal bh7_w90_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_copy788_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid789_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid789_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w90_18_c1 :  std_logic;
signal bh7_w91_16_c1 :  std_logic;
signal bh7_w92_15_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_copy790_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid791_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w92_16_c1 :  std_logic;
signal bh7_w93_17_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_copy792_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid793_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid793_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w93_18_c1 :  std_logic;
signal bh7_w94_16_c1 :  std_logic;
signal bh7_w95_15_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_copy794_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid795_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w95_16_c1 :  std_logic;
signal bh7_w96_17_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_copy796_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid797_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid797_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w96_18_c1 :  std_logic;
signal bh7_w97_16_c1 :  std_logic;
signal bh7_w98_15_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_copy798_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid799_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid799_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w98_16_c1 :  std_logic;
signal bh7_w99_16_c1 :  std_logic;
signal bh7_w100_13_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_copy800_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid801_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid801_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w102_11_c1 :  std_logic;
signal bh7_w103_10_c1 :  std_logic;
signal bh7_w104_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_copy802_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid803_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w105_8_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_copy804_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid805_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid805_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w19_4_c1 :  std_logic;
signal bh7_w20_3_c1 :  std_logic;
signal bh7_w21_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_copy806_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid807_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid807_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_5_c1 :  std_logic;
signal bh7_w22_3_c1 :  std_logic;
signal bh7_w23_4_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_copy808_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid809_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid809_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w23_5_c1 :  std_logic;
signal bh7_w24_5_c1 :  std_logic;
signal bh7_w25_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_copy810_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid811_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid811_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w25_5_c1 :  std_logic;
signal bh7_w26_5_c1 :  std_logic;
signal bh7_w27_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_copy812_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid813_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid813_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w27_5_c1 :  std_logic;
signal bh7_w28_5_c1 :  std_logic;
signal bh7_w29_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_copy814_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid815_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid815_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_5_c1 :  std_logic;
signal bh7_w30_5_c1 :  std_logic;
signal bh7_w31_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_copy816_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid817_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid817_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_5_c1 :  std_logic;
signal bh7_w32_5_c1 :  std_logic;
signal bh7_w33_4_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_copy818_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid819_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid819_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_5_c1 :  std_logic;
signal bh7_w34_6_c1 :  std_logic;
signal bh7_w35_6_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_copy820_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid821_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w35_7_c1 :  std_logic;
signal bh7_w36_7_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_copy822_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid823_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid823_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w36_8_c1 :  std_logic;
signal bh7_w37_6_c1 :  std_logic;
signal bh7_w38_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_copy824_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid825_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid825_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w38_8_c1 :  std_logic;
signal bh7_w39_6_c1 :  std_logic;
signal bh7_w40_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_copy826_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid827_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid827_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w40_8_c1 :  std_logic;
signal bh7_w41_6_c1 :  std_logic;
signal bh7_w42_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_copy828_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid829_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid829_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w42_8_c1 :  std_logic;
signal bh7_w43_6_c1 :  std_logic;
signal bh7_w44_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_copy830_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid831_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid831_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w44_8_c1 :  std_logic;
signal bh7_w45_6_c1 :  std_logic;
signal bh7_w46_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_copy832_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid833_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid833_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w46_8_c1 :  std_logic;
signal bh7_w47_6_c1 :  std_logic;
signal bh7_w48_8_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_copy834_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid835_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid835_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w48_9_c1 :  std_logic;
signal bh7_w49_8_c1 :  std_logic;
signal bh7_w50_10_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_copy836_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid837_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid837_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w50_11_c1 :  std_logic;
signal bh7_w51_14_c1 :  std_logic;
signal bh7_w52_15_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_copy838_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid839_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid839_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w52_16_c1 :  std_logic;
signal bh7_w53_18_c1 :  std_logic;
signal bh7_w54_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_copy840_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid841_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid841_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w54_20_c1 :  std_logic;
signal bh7_w55_21_c1 :  std_logic;
signal bh7_w56_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_copy842_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid843_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid843_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_20_c1 :  std_logic;
signal bh7_w57_24_c1 :  std_logic;
signal bh7_w58_23_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_copy844_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid845_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c0, Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w58_24_c1 :  std_logic;
signal bh7_w59_21_c1 :  std_logic;
signal bh7_w60_22_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_copy846_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid847_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid847_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w59_22_c1 :  std_logic;
signal bh7_w60_23_c1 :  std_logic;
signal bh7_w61_23_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_copy848_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid849_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w61_24_c1 :  std_logic;
signal bh7_w62_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_copy850_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid851_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid851_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_21_c1 :  std_logic;
signal bh7_w63_23_c1 :  std_logic;
signal bh7_w64_23_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_copy852_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid853_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c0, Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w63_24_c1 :  std_logic;
signal bh7_w64_24_c1 :  std_logic;
signal bh7_w65_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_copy854_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid855_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid855_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_25_c1 :  std_logic;
signal bh7_w65_19_c1 :  std_logic;
signal bh7_w66_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_copy856_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid857_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w66_23_c1 :  std_logic;
signal bh7_w67_20_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_copy858_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid859_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid859_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w67_21_c1 :  std_logic;
signal bh7_w68_22_c1 :  std_logic;
signal bh7_w69_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_copy860_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid861_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid861_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w69_20_c1 :  std_logic;
signal bh7_w70_22_c1 :  std_logic;
signal bh7_w71_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_copy862_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid863_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w71_20_c1 :  std_logic;
signal bh7_w72_23_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_copy864_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid865_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid865_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w72_24_c1 :  std_logic;
signal bh7_w73_18_c1 :  std_logic;
signal bh7_w74_24_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_copy866_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid867_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid867_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w74_25_c1 :  std_logic;
signal bh7_w75_17_c1 :  std_logic;
signal bh7_w76_22_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_copy868_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid869_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid869_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w76_23_c1 :  std_logic;
signal bh7_w77_17_c1 :  std_logic;
signal bh7_w78_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_copy870_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid871_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid871_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_23_c1 :  std_logic;
signal bh7_w79_17_c1 :  std_logic;
signal bh7_w80_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_copy872_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid873_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid873_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_23_c1 :  std_logic;
signal bh7_w81_17_c1 :  std_logic;
signal bh7_w82_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_copy874_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid875_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_c1 :  std_logic_vector(1 downto 0);
signal bh7_w82_23_c1 :  std_logic;
signal bh7_w83_16_c1 :  std_logic;
signal Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_copy876_c1 :  std_logic_vector(1 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid877_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid877_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w84_21_c1 :  std_logic;
signal bh7_w85_17_c1 :  std_logic;
signal bh7_w86_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_copy878_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid879_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid879_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_20_c1 :  std_logic;
signal bh7_w87_18_c1 :  std_logic;
signal bh7_w88_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_copy880_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid881_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid881_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_20_c1 :  std_logic;
signal bh7_w89_16_c1 :  std_logic;
signal bh7_w90_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_copy882_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid883_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid883_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w90_20_c1 :  std_logic;
signal bh7_w91_17_c1 :  std_logic;
signal bh7_w92_17_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_copy884_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid885_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid885_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w92_18_c1 :  std_logic;
signal bh7_w93_19_c1 :  std_logic;
signal bh7_w94_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_copy886_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid887_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid887_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w95_17_c1 :  std_logic;
signal bh7_w96_19_c1 :  std_logic;
signal bh7_w97_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_copy888_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid889_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid889_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w98_17_c1 :  std_logic;
signal bh7_w99_17_c1 :  std_logic;
signal bh7_w100_14_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_copy890_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid891_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid891_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w100_15_c1 :  std_logic;
signal bh7_w101_12_c1 :  std_logic;
signal bh7_w102_12_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_copy892_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid893_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid893_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w104_7_c1 :  std_logic;
signal bh7_w105_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_copy894_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid895_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid895_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w21_6_c1 :  std_logic;
signal bh7_w22_4_c1 :  std_logic;
signal bh7_w23_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_copy896_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid897_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid897_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w23_7_c1 :  std_logic;
signal bh7_w24_6_c1 :  std_logic;
signal bh7_w25_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_copy898_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid899_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid899_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w25_7_c1 :  std_logic;
signal bh7_w26_6_c1 :  std_logic;
signal bh7_w27_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_copy900_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid901_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid901_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w27_7_c1 :  std_logic;
signal bh7_w28_6_c1 :  std_logic;
signal bh7_w29_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_copy902_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid903_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid903_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w29_7_c1 :  std_logic;
signal bh7_w30_6_c1 :  std_logic;
signal bh7_w31_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_copy904_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid905_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid905_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w31_7_c1 :  std_logic;
signal bh7_w32_6_c1 :  std_logic;
signal bh7_w33_6_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_copy906_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid907_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid907_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w33_7_c1 :  std_logic;
signal bh7_w34_7_c1 :  std_logic;
signal bh7_w35_8_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_copy908_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid909_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid909_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w35_9_c1 :  std_logic;
signal bh7_w36_9_c1 :  std_logic;
signal bh7_w37_7_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_copy910_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid911_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid911_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w38_9_c1 :  std_logic;
signal bh7_w39_7_c1 :  std_logic;
signal bh7_w40_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_copy912_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid913_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid913_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w40_10_c1 :  std_logic;
signal bh7_w41_7_c1 :  std_logic;
signal bh7_w42_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_copy914_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid915_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid915_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w42_10_c1 :  std_logic;
signal bh7_w43_7_c1 :  std_logic;
signal bh7_w44_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_copy916_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid917_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid917_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w44_10_c1 :  std_logic;
signal bh7_w45_7_c1 :  std_logic;
signal bh7_w46_9_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_copy918_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid919_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid919_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w46_10_c1 :  std_logic;
signal bh7_w47_7_c1 :  std_logic;
signal bh7_w48_10_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_copy920_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid921_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid921_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w48_11_c1 :  std_logic;
signal bh7_w49_9_c1 :  std_logic;
signal bh7_w50_12_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_copy922_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid923_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid923_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w50_13_c1 :  std_logic;
signal bh7_w51_15_c1 :  std_logic;
signal bh7_w52_17_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_copy924_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid925_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid925_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w52_18_c1 :  std_logic;
signal bh7_w53_19_c1 :  std_logic;
signal bh7_w54_21_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_copy926_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid927_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid927_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w54_22_c1 :  std_logic;
signal bh7_w55_22_c1 :  std_logic;
signal bh7_w56_21_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_copy928_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid929_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid929_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w56_22_c1 :  std_logic;
signal bh7_w57_25_c1 :  std_logic;
signal bh7_w58_25_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_copy930_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid931_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid931_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w58_26_c1 :  std_logic;
signal bh7_w59_23_c1 :  std_logic;
signal bh7_w60_24_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_copy932_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid933_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid933_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w60_25_c1 :  std_logic;
signal bh7_w61_25_c1 :  std_logic;
signal bh7_w62_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_copy934_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid935_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid935_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w62_23_c1 :  std_logic;
signal bh7_w63_25_c1 :  std_logic;
signal bh7_w64_26_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_copy936_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid937_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid937_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w64_27_c1 :  std_logic;
signal bh7_w65_20_c1 :  std_logic;
signal bh7_w66_24_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_copy938_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid939_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid939_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w66_25_c1 :  std_logic;
signal bh7_w67_22_c1 :  std_logic;
signal bh7_w68_23_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_copy940_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid941_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid941_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w68_24_c1 :  std_logic;
signal bh7_w69_21_c1 :  std_logic;
signal bh7_w70_23_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_copy942_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid943_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid943_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w71_21_c1 :  std_logic;
signal bh7_w72_25_c1 :  std_logic;
signal bh7_w73_19_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_copy944_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid945_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid945_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w73_20_c1 :  std_logic;
signal bh7_w74_26_c1 :  std_logic;
signal bh7_w75_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_copy946_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid947_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid947_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w75_19_c1 :  std_logic;
signal bh7_w76_24_c1 :  std_logic;
signal bh7_w77_18_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_copy948_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid949_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid949_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w78_24_c1 :  std_logic;
signal bh7_w79_18_c1 :  std_logic;
signal bh7_w80_24_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_copy950_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid951_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid951_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w80_25_c1 :  std_logic;
signal bh7_w81_18_c1 :  std_logic;
signal bh7_w82_24_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_copy952_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid953_In0_c1 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid953_In1_c1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w82_25_c1 :  std_logic;
signal bh7_w83_17_c1 :  std_logic;
signal bh7_w84_22_c1 :  std_logic;
signal Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_copy954_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid955_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid955_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w86_21_c1 :  std_logic;
signal bh7_w87_19_c1 :  std_logic;
signal bh7_w88_21_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_copy956_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid957_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid957_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w88_22_c1 :  std_logic;
signal bh7_w89_17_c1 :  std_logic;
signal bh7_w90_21_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_copy958_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid959_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid959_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w90_22_c1 :  std_logic;
signal bh7_w91_18_c1 :  std_logic;
signal bh7_w92_19_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_copy960_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid961_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid961_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w92_20_c1 :  std_logic;
signal bh7_w93_20_c1 :  std_logic;
signal bh7_w94_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_copy962_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid963_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid963_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w94_19_c1 :  std_logic;
signal bh7_w95_18_c1 :  std_logic;
signal bh7_w96_20_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_copy964_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid965_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid965_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w97_18_c1 :  std_logic;
signal bh7_w98_18_c1 :  std_logic;
signal bh7_w99_18_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_copy966_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid967_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid967_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w100_16_c1 :  std_logic;
signal bh7_w101_13_c1 :  std_logic;
signal bh7_w102_13_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_copy968_c1 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid969_In0_c1 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid969_In1_c1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1 :  std_logic_vector(2 downto 0);
signal bh7_w102_14_c1 :  std_logic;
signal bh7_w103_11_c1 :  std_logic;
signal bh7_w104_8_c1 :  std_logic;
signal Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_copy970_c1 :  std_logic_vector(2 downto 0);
signal tmp_bitheapResult_bh7_22_c1, tmp_bitheapResult_bh7_22_c2 :  std_logic_vector(22 downto 0);
signal bitheapFinalAdd_bh7_In0_c1 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_In1_c1 :  std_logic_vector(83 downto 0);
signal bitheapFinalAdd_bh7_Cin_c0 :  std_logic;
signal bitheapFinalAdd_bh7_Out_c2 :  std_logic_vector(83 downto 0);
signal bitheapResult_bh7_c2 :  std_logic_vector(105 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               bh7_w0_0_c1 <= bh7_w0_0_c0;
               bh7_w1_0_c1 <= bh7_w1_0_c0;
               bh7_w2_0_c1 <= bh7_w2_0_c0;
               bh7_w3_0_c1 <= bh7_w3_0_c0;
               bh7_w4_0_c1 <= bh7_w4_0_c0;
               bh7_w5_0_c1 <= bh7_w5_0_c0;
               bh7_w6_0_c1 <= bh7_w6_0_c0;
               bh7_w7_0_c1 <= bh7_w7_0_c0;
               bh7_w8_0_c1 <= bh7_w8_0_c0;
               bh7_w9_0_c1 <= bh7_w9_0_c0;
               bh7_w10_0_c1 <= bh7_w10_0_c0;
               bh7_w11_0_c1 <= bh7_w11_0_c0;
               bh7_w12_0_c1 <= bh7_w12_0_c0;
               bh7_w13_0_c1 <= bh7_w13_0_c0;
               bh7_w14_0_c1 <= bh7_w14_0_c0;
               bh7_w15_0_c1 <= bh7_w15_0_c0;
               bh7_w16_0_c1 <= bh7_w16_0_c0;
               bh7_w59_0_c1 <= bh7_w59_0_c0;
               bh7_w60_0_c1 <= bh7_w60_0_c0;
               bh7_w61_0_c1 <= bh7_w61_0_c0;
               bh7_w62_0_c1 <= bh7_w62_0_c0;
               bh7_w64_0_c1 <= bh7_w64_0_c0;
               bh7_w65_0_c1 <= bh7_w65_0_c0;
               bh7_w67_0_c1 <= bh7_w67_0_c0;
               bh7_w69_0_c1 <= bh7_w69_0_c0;
               bh7_w70_0_c1 <= bh7_w70_0_c0;
               bh7_w72_0_c1 <= bh7_w72_0_c0;
               bh7_w74_0_c1 <= bh7_w74_0_c0;
               bh7_w25_2_c1 <= bh7_w25_2_c0;
               bh7_w27_2_c1 <= bh7_w27_2_c0;
               bh7_w29_2_c1 <= bh7_w29_2_c0;
               bh7_w31_2_c1 <= bh7_w31_2_c0;
               bh7_w33_2_c1 <= bh7_w33_2_c0;
               bh7_w59_2_c1 <= bh7_w59_2_c0;
               bh7_w60_3_c1 <= bh7_w60_3_c0;
               bh7_w61_3_c1 <= bh7_w61_3_c0;
               bh7_w62_2_c1 <= bh7_w62_2_c0;
               bh7_w64_3_c1 <= bh7_w64_3_c0;
               bh7_w48_3_c1 <= bh7_w48_3_c0;
               bh7_w59_3_c1 <= bh7_w59_3_c0;
               bh7_w60_4_c1 <= bh7_w60_4_c0;
               bh7_w61_4_c1 <= bh7_w61_4_c0;
               bh7_w62_3_c1 <= bh7_w62_3_c0;
               bh7_w64_4_c1 <= bh7_w64_4_c0;
               bh7_w65_2_c1 <= bh7_w65_2_c0;
               bh7_w67_3_c1 <= bh7_w67_3_c0;
               bh7_w69_3_c1 <= bh7_w69_3_c0;
               bh7_w70_3_c1 <= bh7_w70_3_c0;
               bh7_w72_3_c1 <= bh7_w72_3_c0;
               bh7_w74_2_c1 <= bh7_w74_2_c0;
               bh7_w76_1_c1 <= bh7_w76_1_c0;
               bh7_w77_0_c1 <= bh7_w77_0_c0;
               bh7_w78_0_c1 <= bh7_w78_0_c0;
               bh7_w79_0_c1 <= bh7_w79_0_c0;
               bh7_w80_0_c1 <= bh7_w80_0_c0;
               bh7_w81_0_c1 <= bh7_w81_0_c0;
               bh7_w58_5_c1 <= bh7_w58_5_c0;
               bh7_w59_4_c1 <= bh7_w59_4_c0;
               bh7_w60_5_c1 <= bh7_w60_5_c0;
               bh7_w61_5_c1 <= bh7_w61_5_c0;
               bh7_w62_4_c1 <= bh7_w62_4_c0;
               bh7_w63_5_c1 <= bh7_w63_5_c0;
               bh7_w64_5_c1 <= bh7_w64_5_c0;
               bh7_w65_3_c1 <= bh7_w65_3_c0;
               bh7_w67_4_c1 <= bh7_w67_4_c0;
               bh7_w69_4_c1 <= bh7_w69_4_c0;
               bh7_w70_4_c1 <= bh7_w70_4_c0;
               bh7_w72_4_c1 <= bh7_w72_4_c0;
               bh7_w74_3_c1 <= bh7_w74_3_c0;
               bh7_w75_2_c1 <= bh7_w75_2_c0;
               bh7_w76_2_c1 <= bh7_w76_2_c0;
               bh7_w77_1_c1 <= bh7_w77_1_c0;
               bh7_w78_1_c1 <= bh7_w78_1_c0;
               bh7_w79_1_c1 <= bh7_w79_1_c0;
               bh7_w80_1_c1 <= bh7_w80_1_c0;
               bh7_w81_1_c1 <= bh7_w81_1_c0;
               bh7_w82_0_c1 <= bh7_w82_0_c0;
               bh7_w83_0_c1 <= bh7_w83_0_c0;
               bh7_w84_0_c1 <= bh7_w84_0_c0;
               bh7_w85_0_c1 <= bh7_w85_0_c0;
               bh7_w86_0_c1 <= bh7_w86_0_c0;
               bh7_w87_0_c1 <= bh7_w87_0_c0;
               bh7_w88_0_c1 <= bh7_w88_0_c0;
               bh7_w89_0_c1 <= bh7_w89_0_c0;
               bh7_w90_0_c1 <= bh7_w90_0_c0;
               bh7_w91_0_c1 <= bh7_w91_0_c0;
               bh7_w92_0_c1 <= bh7_w92_0_c0;
               bh7_w93_0_c1 <= bh7_w93_0_c0;
               bh7_w94_0_c1 <= bh7_w94_0_c0;
               bh7_w95_0_c1 <= bh7_w95_0_c0;
               bh7_w96_0_c1 <= bh7_w96_0_c0;
               bh7_w97_0_c1 <= bh7_w97_0_c0;
               bh7_w98_0_c1 <= bh7_w98_0_c0;
               bh7_w61_18_c1 <= bh7_w61_18_c0;
               bh7_w64_18_c1 <= bh7_w64_18_c0;
               bh7_w67_15_c1 <= bh7_w67_15_c0;
               bh7_w90_15_c1 <= bh7_w90_15_c0;
               bh7_w93_15_c1 <= bh7_w93_15_c0;
               bh7_w96_15_c1 <= bh7_w96_15_c0;
               bh7_w99_14_c1 <= bh7_w99_14_c0;
               bh7_w102_9_c1 <= bh7_w102_9_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c0;
               Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c0;
               Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c0;
               Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c0;
            end if;
            if ce_2 = '1' then
               tmp_bitheapResult_bh7_22_c2 <= tmp_bitheapResult_bh7_22_c1;
            end if;
         end if;
      end process;
   XX_m6_c0 <= X ;
   YY_m6_c0 <= Y ;
   tile_0_X_c0 <= X(16 downto 0);
   tile_0_Y_c0 <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_Freq300_uid9
      port map ( clk  => clk,
                 X => tile_0_X_c0,
                 Y => tile_0_Y_c0,
                 R => tile_0_output_c0);

   tile_0_filtered_output_c0 <= unsigned(tile_0_output_c0(40 downto 0));
   bh7_w0_0_c0 <= tile_0_filtered_output_c0(0);
   bh7_w1_0_c0 <= tile_0_filtered_output_c0(1);
   bh7_w2_0_c0 <= tile_0_filtered_output_c0(2);
   bh7_w3_0_c0 <= tile_0_filtered_output_c0(3);
   bh7_w4_0_c0 <= tile_0_filtered_output_c0(4);
   bh7_w5_0_c0 <= tile_0_filtered_output_c0(5);
   bh7_w6_0_c0 <= tile_0_filtered_output_c0(6);
   bh7_w7_0_c0 <= tile_0_filtered_output_c0(7);
   bh7_w8_0_c0 <= tile_0_filtered_output_c0(8);
   bh7_w9_0_c0 <= tile_0_filtered_output_c0(9);
   bh7_w10_0_c0 <= tile_0_filtered_output_c0(10);
   bh7_w11_0_c0 <= tile_0_filtered_output_c0(11);
   bh7_w12_0_c0 <= tile_0_filtered_output_c0(12);
   bh7_w13_0_c0 <= tile_0_filtered_output_c0(13);
   bh7_w14_0_c0 <= tile_0_filtered_output_c0(14);
   bh7_w15_0_c0 <= tile_0_filtered_output_c0(15);
   bh7_w16_0_c0 <= tile_0_filtered_output_c0(16);
   bh7_w17_0_c0 <= tile_0_filtered_output_c0(17);
   bh7_w18_0_c0 <= tile_0_filtered_output_c0(18);
   bh7_w19_0_c0 <= tile_0_filtered_output_c0(19);
   bh7_w20_0_c0 <= tile_0_filtered_output_c0(20);
   bh7_w21_0_c0 <= tile_0_filtered_output_c0(21);
   bh7_w22_0_c0 <= tile_0_filtered_output_c0(22);
   bh7_w23_0_c0 <= tile_0_filtered_output_c0(23);
   bh7_w24_0_c0 <= tile_0_filtered_output_c0(24);
   bh7_w25_0_c0 <= tile_0_filtered_output_c0(25);
   bh7_w26_0_c0 <= tile_0_filtered_output_c0(26);
   bh7_w27_0_c0 <= tile_0_filtered_output_c0(27);
   bh7_w28_0_c0 <= tile_0_filtered_output_c0(28);
   bh7_w29_0_c0 <= tile_0_filtered_output_c0(29);
   bh7_w30_0_c0 <= tile_0_filtered_output_c0(30);
   bh7_w31_0_c0 <= tile_0_filtered_output_c0(31);
   bh7_w32_0_c0 <= tile_0_filtered_output_c0(32);
   bh7_w33_0_c0 <= tile_0_filtered_output_c0(33);
   bh7_w34_0_c0 <= tile_0_filtered_output_c0(34);
   bh7_w35_0_c0 <= tile_0_filtered_output_c0(35);
   bh7_w36_0_c0 <= tile_0_filtered_output_c0(36);
   bh7_w37_0_c0 <= tile_0_filtered_output_c0(37);
   bh7_w38_0_c0 <= tile_0_filtered_output_c0(38);
   bh7_w39_0_c0 <= tile_0_filtered_output_c0(39);
   bh7_w40_0_c0 <= tile_0_filtered_output_c0(40);
   tile_1_X_c0 <= X(33 downto 17);
   tile_1_Y_c0 <= Y(23 downto 0);
   tile_1_mult: DSPBlock_17x24_Freq300_uid11
      port map ( clk  => clk,
                 X => tile_1_X_c0,
                 Y => tile_1_Y_c0,
                 R => tile_1_output_c0);

   tile_1_filtered_output_c0 <= unsigned(tile_1_output_c0(40 downto 0));
   bh7_w17_1_c0 <= tile_1_filtered_output_c0(0);
   bh7_w18_1_c0 <= tile_1_filtered_output_c0(1);
   bh7_w19_1_c0 <= tile_1_filtered_output_c0(2);
   bh7_w20_1_c0 <= tile_1_filtered_output_c0(3);
   bh7_w21_1_c0 <= tile_1_filtered_output_c0(4);
   bh7_w22_1_c0 <= tile_1_filtered_output_c0(5);
   bh7_w23_1_c0 <= tile_1_filtered_output_c0(6);
   bh7_w24_1_c0 <= tile_1_filtered_output_c0(7);
   bh7_w25_1_c0 <= tile_1_filtered_output_c0(8);
   bh7_w26_1_c0 <= tile_1_filtered_output_c0(9);
   bh7_w27_1_c0 <= tile_1_filtered_output_c0(10);
   bh7_w28_1_c0 <= tile_1_filtered_output_c0(11);
   bh7_w29_1_c0 <= tile_1_filtered_output_c0(12);
   bh7_w30_1_c0 <= tile_1_filtered_output_c0(13);
   bh7_w31_1_c0 <= tile_1_filtered_output_c0(14);
   bh7_w32_1_c0 <= tile_1_filtered_output_c0(15);
   bh7_w33_1_c0 <= tile_1_filtered_output_c0(16);
   bh7_w34_1_c0 <= tile_1_filtered_output_c0(17);
   bh7_w35_1_c0 <= tile_1_filtered_output_c0(18);
   bh7_w36_1_c0 <= tile_1_filtered_output_c0(19);
   bh7_w37_1_c0 <= tile_1_filtered_output_c0(20);
   bh7_w38_1_c0 <= tile_1_filtered_output_c0(21);
   bh7_w39_1_c0 <= tile_1_filtered_output_c0(22);
   bh7_w40_1_c0 <= tile_1_filtered_output_c0(23);
   bh7_w41_0_c0 <= tile_1_filtered_output_c0(24);
   bh7_w42_0_c0 <= tile_1_filtered_output_c0(25);
   bh7_w43_0_c0 <= tile_1_filtered_output_c0(26);
   bh7_w44_0_c0 <= tile_1_filtered_output_c0(27);
   bh7_w45_0_c0 <= tile_1_filtered_output_c0(28);
   bh7_w46_0_c0 <= tile_1_filtered_output_c0(29);
   bh7_w47_0_c0 <= tile_1_filtered_output_c0(30);
   bh7_w48_0_c0 <= tile_1_filtered_output_c0(31);
   bh7_w49_0_c0 <= tile_1_filtered_output_c0(32);
   bh7_w50_0_c0 <= tile_1_filtered_output_c0(33);
   bh7_w51_0_c0 <= tile_1_filtered_output_c0(34);
   bh7_w52_0_c0 <= tile_1_filtered_output_c0(35);
   bh7_w53_0_c0 <= tile_1_filtered_output_c0(36);
   bh7_w54_0_c0 <= tile_1_filtered_output_c0(37);
   bh7_w55_0_c0 <= tile_1_filtered_output_c0(38);
   bh7_w56_0_c0 <= tile_1_filtered_output_c0(39);
   bh7_w57_0_c0 <= tile_1_filtered_output_c0(40);
   tile_2_X_c0 <= X(50 downto 34);
   tile_2_Y_c0 <= Y(23 downto 0);
   tile_2_mult: DSPBlock_17x24_Freq300_uid13
      port map ( clk  => clk,
                 X => tile_2_X_c0,
                 Y => tile_2_Y_c0,
                 R => tile_2_output_c0);

   tile_2_filtered_output_c0 <= unsigned(tile_2_output_c0(40 downto 0));
   bh7_w34_2_c0 <= tile_2_filtered_output_c0(0);
   bh7_w35_2_c0 <= tile_2_filtered_output_c0(1);
   bh7_w36_2_c0 <= tile_2_filtered_output_c0(2);
   bh7_w37_2_c0 <= tile_2_filtered_output_c0(3);
   bh7_w38_2_c0 <= tile_2_filtered_output_c0(4);
   bh7_w39_2_c0 <= tile_2_filtered_output_c0(5);
   bh7_w40_2_c0 <= tile_2_filtered_output_c0(6);
   bh7_w41_1_c0 <= tile_2_filtered_output_c0(7);
   bh7_w42_1_c0 <= tile_2_filtered_output_c0(8);
   bh7_w43_1_c0 <= tile_2_filtered_output_c0(9);
   bh7_w44_1_c0 <= tile_2_filtered_output_c0(10);
   bh7_w45_1_c0 <= tile_2_filtered_output_c0(11);
   bh7_w46_1_c0 <= tile_2_filtered_output_c0(12);
   bh7_w47_1_c0 <= tile_2_filtered_output_c0(13);
   bh7_w48_1_c0 <= tile_2_filtered_output_c0(14);
   bh7_w49_1_c0 <= tile_2_filtered_output_c0(15);
   bh7_w50_1_c0 <= tile_2_filtered_output_c0(16);
   bh7_w51_1_c0 <= tile_2_filtered_output_c0(17);
   bh7_w52_1_c0 <= tile_2_filtered_output_c0(18);
   bh7_w53_1_c0 <= tile_2_filtered_output_c0(19);
   bh7_w54_1_c0 <= tile_2_filtered_output_c0(20);
   bh7_w55_1_c0 <= tile_2_filtered_output_c0(21);
   bh7_w56_1_c0 <= tile_2_filtered_output_c0(22);
   bh7_w57_1_c0 <= tile_2_filtered_output_c0(23);
   bh7_w58_0_c0 <= tile_2_filtered_output_c0(24);
   bh7_w59_0_c0 <= tile_2_filtered_output_c0(25);
   bh7_w60_0_c0 <= tile_2_filtered_output_c0(26);
   bh7_w61_0_c0 <= tile_2_filtered_output_c0(27);
   bh7_w62_0_c0 <= tile_2_filtered_output_c0(28);
   bh7_w63_0_c0 <= tile_2_filtered_output_c0(29);
   bh7_w64_0_c0 <= tile_2_filtered_output_c0(30);
   bh7_w65_0_c0 <= tile_2_filtered_output_c0(31);
   bh7_w66_0_c0 <= tile_2_filtered_output_c0(32);
   bh7_w67_0_c0 <= tile_2_filtered_output_c0(33);
   bh7_w68_0_c0 <= tile_2_filtered_output_c0(34);
   bh7_w69_0_c0 <= tile_2_filtered_output_c0(35);
   bh7_w70_0_c0 <= tile_2_filtered_output_c0(36);
   bh7_w71_0_c0 <= tile_2_filtered_output_c0(37);
   bh7_w72_0_c0 <= tile_2_filtered_output_c0(38);
   bh7_w73_0_c0 <= tile_2_filtered_output_c0(39);
   bh7_w74_0_c0 <= tile_2_filtered_output_c0(40);
   tile_3_X_c0 <= X(52 downto 51);
   tile_3_Y_c0 <= Y(23 downto 21);
   tile_3_mult: IntMultiplierLUT_2x3_Freq300_uid15
      port map ( clk  => clk,
                 X => tile_3_X_c0,
                 Y => tile_3_Y_c0,
                 R => tile_3_output_c0);

   tile_3_filtered_output_c0 <= unsigned(tile_3_output_c0(4 downto 0));
   bh7_w72_1_c0 <= tile_3_filtered_output_c0(0);
   bh7_w73_1_c0 <= tile_3_filtered_output_c0(1);
   bh7_w74_1_c0 <= tile_3_filtered_output_c0(2);
   bh7_w75_0_c0 <= tile_3_filtered_output_c0(3);
   bh7_w76_0_c0 <= tile_3_filtered_output_c0(4);
   tile_4_X_c0 <= X(52 downto 51);
   tile_4_Y_c0 <= Y(20 downto 18);
   tile_4_mult: IntMultiplierLUT_2x3_Freq300_uid20
      port map ( clk  => clk,
                 X => tile_4_X_c0,
                 Y => tile_4_Y_c0,
                 R => tile_4_output_c0);

   tile_4_filtered_output_c0 <= unsigned(tile_4_output_c0(4 downto 0));
   bh7_w69_1_c0 <= tile_4_filtered_output_c0(0);
   bh7_w70_1_c0 <= tile_4_filtered_output_c0(1);
   bh7_w71_1_c0 <= tile_4_filtered_output_c0(2);
   bh7_w72_2_c0 <= tile_4_filtered_output_c0(3);
   bh7_w73_2_c0 <= tile_4_filtered_output_c0(4);
   tile_5_X_c0 <= X(52 downto 51);
   tile_5_Y_c0 <= Y(17 downto 15);
   tile_5_mult: IntMultiplierLUT_2x3_Freq300_uid25
      port map ( clk  => clk,
                 X => tile_5_X_c0,
                 Y => tile_5_Y_c0,
                 R => tile_5_output_c0);

   tile_5_filtered_output_c0 <= unsigned(tile_5_output_c0(4 downto 0));
   bh7_w66_1_c0 <= tile_5_filtered_output_c0(0);
   bh7_w67_1_c0 <= tile_5_filtered_output_c0(1);
   bh7_w68_1_c0 <= tile_5_filtered_output_c0(2);
   bh7_w69_2_c0 <= tile_5_filtered_output_c0(3);
   bh7_w70_2_c0 <= tile_5_filtered_output_c0(4);
   tile_6_X_c0 <= X(52 downto 51);
   tile_6_Y_c0 <= Y(14 downto 12);
   tile_6_mult: IntMultiplierLUT_2x3_Freq300_uid30
      port map ( clk  => clk,
                 X => tile_6_X_c0,
                 Y => tile_6_Y_c0,
                 R => tile_6_output_c0);

   tile_6_filtered_output_c0 <= unsigned(tile_6_output_c0(4 downto 0));
   bh7_w63_1_c0 <= tile_6_filtered_output_c0(0);
   bh7_w64_1_c0 <= tile_6_filtered_output_c0(1);
   bh7_w65_1_c0 <= tile_6_filtered_output_c0(2);
   bh7_w66_2_c0 <= tile_6_filtered_output_c0(3);
   bh7_w67_2_c0 <= tile_6_filtered_output_c0(4);
   tile_7_X_c0 <= X(52 downto 51);
   tile_7_Y_c0 <= Y(11 downto 9);
   tile_7_mult: IntMultiplierLUT_2x3_Freq300_uid35
      port map ( clk  => clk,
                 X => tile_7_X_c0,
                 Y => tile_7_Y_c0,
                 R => tile_7_output_c0);

   tile_7_filtered_output_c0 <= unsigned(tile_7_output_c0(4 downto 0));
   bh7_w60_1_c0 <= tile_7_filtered_output_c0(0);
   bh7_w61_1_c0 <= tile_7_filtered_output_c0(1);
   bh7_w62_1_c0 <= tile_7_filtered_output_c0(2);
   bh7_w63_2_c0 <= tile_7_filtered_output_c0(3);
   bh7_w64_2_c0 <= tile_7_filtered_output_c0(4);
   tile_8_X_c0 <= X(52 downto 51);
   tile_8_Y_c0 <= Y(8 downto 6);
   tile_8_mult: IntMultiplierLUT_2x3_Freq300_uid40
      port map ( clk  => clk,
                 X => tile_8_X_c0,
                 Y => tile_8_Y_c0,
                 R => tile_8_output_c0);

   tile_8_filtered_output_c0 <= unsigned(tile_8_output_c0(4 downto 0));
   bh7_w57_2_c0 <= tile_8_filtered_output_c0(0);
   bh7_w58_1_c0 <= tile_8_filtered_output_c0(1);
   bh7_w59_1_c0 <= tile_8_filtered_output_c0(2);
   bh7_w60_2_c0 <= tile_8_filtered_output_c0(3);
   bh7_w61_2_c0 <= tile_8_filtered_output_c0(4);
   tile_9_X_c0 <= X(52 downto 51);
   tile_9_Y_c0 <= Y(5 downto 3);
   tile_9_mult: IntMultiplierLUT_2x3_Freq300_uid45
      port map ( clk  => clk,
                 X => tile_9_X_c0,
                 Y => tile_9_Y_c0,
                 R => tile_9_output_c0);

   tile_9_filtered_output_c0 <= unsigned(tile_9_output_c0(4 downto 0));
   bh7_w54_2_c0 <= tile_9_filtered_output_c0(0);
   bh7_w55_2_c0 <= tile_9_filtered_output_c0(1);
   bh7_w56_2_c0 <= tile_9_filtered_output_c0(2);
   bh7_w57_3_c0 <= tile_9_filtered_output_c0(3);
   bh7_w58_2_c0 <= tile_9_filtered_output_c0(4);
   tile_10_X_c0 <= X(52 downto 51);
   tile_10_Y_c0 <= Y(2 downto 0);
   tile_10_mult: IntMultiplierLUT_2x3_Freq300_uid50
      port map ( clk  => clk,
                 X => tile_10_X_c0,
                 Y => tile_10_Y_c0,
                 R => tile_10_output_c0);

   tile_10_filtered_output_c0 <= unsigned(tile_10_output_c0(4 downto 0));
   bh7_w51_2_c0 <= tile_10_filtered_output_c0(0);
   bh7_w52_2_c0 <= tile_10_filtered_output_c0(1);
   bh7_w53_2_c0 <= tile_10_filtered_output_c0(2);
   bh7_w54_3_c0 <= tile_10_filtered_output_c0(3);
   bh7_w55_3_c0 <= tile_10_filtered_output_c0(4);
   tile_11_X_c0 <= X(16 downto 0);
   tile_11_Y_c0 <= Y(47 downto 24);
   tile_11_mult: DSPBlock_17x24_Freq300_uid55
      port map ( clk  => clk,
                 X => tile_11_X_c0,
                 Y => tile_11_Y_c0,
                 R => tile_11_output_c0);

   tile_11_filtered_output_c0 <= unsigned(tile_11_output_c0(40 downto 0));
   bh7_w24_2_c0 <= tile_11_filtered_output_c0(0);
   bh7_w25_2_c0 <= tile_11_filtered_output_c0(1);
   bh7_w26_2_c0 <= tile_11_filtered_output_c0(2);
   bh7_w27_2_c0 <= tile_11_filtered_output_c0(3);
   bh7_w28_2_c0 <= tile_11_filtered_output_c0(4);
   bh7_w29_2_c0 <= tile_11_filtered_output_c0(5);
   bh7_w30_2_c0 <= tile_11_filtered_output_c0(6);
   bh7_w31_2_c0 <= tile_11_filtered_output_c0(7);
   bh7_w32_2_c0 <= tile_11_filtered_output_c0(8);
   bh7_w33_2_c0 <= tile_11_filtered_output_c0(9);
   bh7_w34_3_c0 <= tile_11_filtered_output_c0(10);
   bh7_w35_3_c0 <= tile_11_filtered_output_c0(11);
   bh7_w36_3_c0 <= tile_11_filtered_output_c0(12);
   bh7_w37_3_c0 <= tile_11_filtered_output_c0(13);
   bh7_w38_3_c0 <= tile_11_filtered_output_c0(14);
   bh7_w39_3_c0 <= tile_11_filtered_output_c0(15);
   bh7_w40_3_c0 <= tile_11_filtered_output_c0(16);
   bh7_w41_2_c0 <= tile_11_filtered_output_c0(17);
   bh7_w42_2_c0 <= tile_11_filtered_output_c0(18);
   bh7_w43_2_c0 <= tile_11_filtered_output_c0(19);
   bh7_w44_2_c0 <= tile_11_filtered_output_c0(20);
   bh7_w45_2_c0 <= tile_11_filtered_output_c0(21);
   bh7_w46_2_c0 <= tile_11_filtered_output_c0(22);
   bh7_w47_2_c0 <= tile_11_filtered_output_c0(23);
   bh7_w48_2_c0 <= tile_11_filtered_output_c0(24);
   bh7_w49_2_c0 <= tile_11_filtered_output_c0(25);
   bh7_w50_2_c0 <= tile_11_filtered_output_c0(26);
   bh7_w51_3_c0 <= tile_11_filtered_output_c0(27);
   bh7_w52_3_c0 <= tile_11_filtered_output_c0(28);
   bh7_w53_3_c0 <= tile_11_filtered_output_c0(29);
   bh7_w54_4_c0 <= tile_11_filtered_output_c0(30);
   bh7_w55_4_c0 <= tile_11_filtered_output_c0(31);
   bh7_w56_3_c0 <= tile_11_filtered_output_c0(32);
   bh7_w57_4_c0 <= tile_11_filtered_output_c0(33);
   bh7_w58_3_c0 <= tile_11_filtered_output_c0(34);
   bh7_w59_2_c0 <= tile_11_filtered_output_c0(35);
   bh7_w60_3_c0 <= tile_11_filtered_output_c0(36);
   bh7_w61_3_c0 <= tile_11_filtered_output_c0(37);
   bh7_w62_2_c0 <= tile_11_filtered_output_c0(38);
   bh7_w63_3_c0 <= tile_11_filtered_output_c0(39);
   bh7_w64_3_c0 <= tile_11_filtered_output_c0(40);
   tile_12_X_c0 <= X(33 downto 17);
   tile_12_Y_c0 <= Y(47 downto 24);
   tile_12_mult: DSPBlock_17x24_Freq300_uid57
      port map ( clk  => clk,
                 X => tile_12_X_c0,
                 Y => tile_12_Y_c0,
                 R => tile_12_output_c0);

   tile_12_filtered_output_c0 <= unsigned(tile_12_output_c0(40 downto 0));
   bh7_w41_3_c0 <= tile_12_filtered_output_c0(0);
   bh7_w42_3_c0 <= tile_12_filtered_output_c0(1);
   bh7_w43_3_c0 <= tile_12_filtered_output_c0(2);
   bh7_w44_3_c0 <= tile_12_filtered_output_c0(3);
   bh7_w45_3_c0 <= tile_12_filtered_output_c0(4);
   bh7_w46_3_c0 <= tile_12_filtered_output_c0(5);
   bh7_w47_3_c0 <= tile_12_filtered_output_c0(6);
   bh7_w48_3_c0 <= tile_12_filtered_output_c0(7);
   bh7_w49_3_c0 <= tile_12_filtered_output_c0(8);
   bh7_w50_3_c0 <= tile_12_filtered_output_c0(9);
   bh7_w51_4_c0 <= tile_12_filtered_output_c0(10);
   bh7_w52_4_c0 <= tile_12_filtered_output_c0(11);
   bh7_w53_4_c0 <= tile_12_filtered_output_c0(12);
   bh7_w54_5_c0 <= tile_12_filtered_output_c0(13);
   bh7_w55_5_c0 <= tile_12_filtered_output_c0(14);
   bh7_w56_4_c0 <= tile_12_filtered_output_c0(15);
   bh7_w57_5_c0 <= tile_12_filtered_output_c0(16);
   bh7_w58_4_c0 <= tile_12_filtered_output_c0(17);
   bh7_w59_3_c0 <= tile_12_filtered_output_c0(18);
   bh7_w60_4_c0 <= tile_12_filtered_output_c0(19);
   bh7_w61_4_c0 <= tile_12_filtered_output_c0(20);
   bh7_w62_3_c0 <= tile_12_filtered_output_c0(21);
   bh7_w63_4_c0 <= tile_12_filtered_output_c0(22);
   bh7_w64_4_c0 <= tile_12_filtered_output_c0(23);
   bh7_w65_2_c0 <= tile_12_filtered_output_c0(24);
   bh7_w66_3_c0 <= tile_12_filtered_output_c0(25);
   bh7_w67_3_c0 <= tile_12_filtered_output_c0(26);
   bh7_w68_2_c0 <= tile_12_filtered_output_c0(27);
   bh7_w69_3_c0 <= tile_12_filtered_output_c0(28);
   bh7_w70_3_c0 <= tile_12_filtered_output_c0(29);
   bh7_w71_2_c0 <= tile_12_filtered_output_c0(30);
   bh7_w72_3_c0 <= tile_12_filtered_output_c0(31);
   bh7_w73_3_c0 <= tile_12_filtered_output_c0(32);
   bh7_w74_2_c0 <= tile_12_filtered_output_c0(33);
   bh7_w75_1_c0 <= tile_12_filtered_output_c0(34);
   bh7_w76_1_c0 <= tile_12_filtered_output_c0(35);
   bh7_w77_0_c0 <= tile_12_filtered_output_c0(36);
   bh7_w78_0_c0 <= tile_12_filtered_output_c0(37);
   bh7_w79_0_c0 <= tile_12_filtered_output_c0(38);
   bh7_w80_0_c0 <= tile_12_filtered_output_c0(39);
   bh7_w81_0_c0 <= tile_12_filtered_output_c0(40);
   tile_13_X_c0 <= X(50 downto 34);
   tile_13_Y_c0 <= Y(47 downto 24);
   tile_13_mult: DSPBlock_17x24_Freq300_uid59
      port map ( clk  => clk,
                 X => tile_13_X_c0,
                 Y => tile_13_Y_c0,
                 R => tile_13_output_c0);

   tile_13_filtered_output_c0 <= unsigned(tile_13_output_c0(40 downto 0));
   bh7_w58_5_c0 <= tile_13_filtered_output_c0(0);
   bh7_w59_4_c0 <= tile_13_filtered_output_c0(1);
   bh7_w60_5_c0 <= tile_13_filtered_output_c0(2);
   bh7_w61_5_c0 <= tile_13_filtered_output_c0(3);
   bh7_w62_4_c0 <= tile_13_filtered_output_c0(4);
   bh7_w63_5_c0 <= tile_13_filtered_output_c0(5);
   bh7_w64_5_c0 <= tile_13_filtered_output_c0(6);
   bh7_w65_3_c0 <= tile_13_filtered_output_c0(7);
   bh7_w66_4_c0 <= tile_13_filtered_output_c0(8);
   bh7_w67_4_c0 <= tile_13_filtered_output_c0(9);
   bh7_w68_3_c0 <= tile_13_filtered_output_c0(10);
   bh7_w69_4_c0 <= tile_13_filtered_output_c0(11);
   bh7_w70_4_c0 <= tile_13_filtered_output_c0(12);
   bh7_w71_3_c0 <= tile_13_filtered_output_c0(13);
   bh7_w72_4_c0 <= tile_13_filtered_output_c0(14);
   bh7_w73_4_c0 <= tile_13_filtered_output_c0(15);
   bh7_w74_3_c0 <= tile_13_filtered_output_c0(16);
   bh7_w75_2_c0 <= tile_13_filtered_output_c0(17);
   bh7_w76_2_c0 <= tile_13_filtered_output_c0(18);
   bh7_w77_1_c0 <= tile_13_filtered_output_c0(19);
   bh7_w78_1_c0 <= tile_13_filtered_output_c0(20);
   bh7_w79_1_c0 <= tile_13_filtered_output_c0(21);
   bh7_w80_1_c0 <= tile_13_filtered_output_c0(22);
   bh7_w81_1_c0 <= tile_13_filtered_output_c0(23);
   bh7_w82_0_c0 <= tile_13_filtered_output_c0(24);
   bh7_w83_0_c0 <= tile_13_filtered_output_c0(25);
   bh7_w84_0_c0 <= tile_13_filtered_output_c0(26);
   bh7_w85_0_c0 <= tile_13_filtered_output_c0(27);
   bh7_w86_0_c0 <= tile_13_filtered_output_c0(28);
   bh7_w87_0_c0 <= tile_13_filtered_output_c0(29);
   bh7_w88_0_c0 <= tile_13_filtered_output_c0(30);
   bh7_w89_0_c0 <= tile_13_filtered_output_c0(31);
   bh7_w90_0_c0 <= tile_13_filtered_output_c0(32);
   bh7_w91_0_c0 <= tile_13_filtered_output_c0(33);
   bh7_w92_0_c0 <= tile_13_filtered_output_c0(34);
   bh7_w93_0_c0 <= tile_13_filtered_output_c0(35);
   bh7_w94_0_c0 <= tile_13_filtered_output_c0(36);
   bh7_w95_0_c0 <= tile_13_filtered_output_c0(37);
   bh7_w96_0_c0 <= tile_13_filtered_output_c0(38);
   bh7_w97_0_c0 <= tile_13_filtered_output_c0(39);
   bh7_w98_0_c0 <= tile_13_filtered_output_c0(40);
   tile_14_X_c0 <= X(52 downto 51);
   tile_14_Y_c0 <= Y(47 downto 45);
   tile_14_mult: IntMultiplierLUT_2x3_Freq300_uid61
      port map ( clk  => clk,
                 X => tile_14_X_c0,
                 Y => tile_14_Y_c0,
                 R => tile_14_output_c0);

   tile_14_filtered_output_c0 <= unsigned(tile_14_output_c0(4 downto 0));
   bh7_w96_1_c0 <= tile_14_filtered_output_c0(0);
   bh7_w97_1_c0 <= tile_14_filtered_output_c0(1);
   bh7_w98_1_c0 <= tile_14_filtered_output_c0(2);
   bh7_w99_0_c0 <= tile_14_filtered_output_c0(3);
   bh7_w100_0_c0 <= tile_14_filtered_output_c0(4);
   tile_15_X_c0 <= X(52 downto 51);
   tile_15_Y_c0 <= Y(44 downto 42);
   tile_15_mult: IntMultiplierLUT_2x3_Freq300_uid66
      port map ( clk  => clk,
                 X => tile_15_X_c0,
                 Y => tile_15_Y_c0,
                 R => tile_15_output_c0);

   tile_15_filtered_output_c0 <= unsigned(tile_15_output_c0(4 downto 0));
   bh7_w93_1_c0 <= tile_15_filtered_output_c0(0);
   bh7_w94_1_c0 <= tile_15_filtered_output_c0(1);
   bh7_w95_1_c0 <= tile_15_filtered_output_c0(2);
   bh7_w96_2_c0 <= tile_15_filtered_output_c0(3);
   bh7_w97_2_c0 <= tile_15_filtered_output_c0(4);
   tile_16_X_c0 <= X(52 downto 51);
   tile_16_Y_c0 <= Y(41 downto 39);
   tile_16_mult: IntMultiplierLUT_2x3_Freq300_uid71
      port map ( clk  => clk,
                 X => tile_16_X_c0,
                 Y => tile_16_Y_c0,
                 R => tile_16_output_c0);

   tile_16_filtered_output_c0 <= unsigned(tile_16_output_c0(4 downto 0));
   bh7_w90_1_c0 <= tile_16_filtered_output_c0(0);
   bh7_w91_1_c0 <= tile_16_filtered_output_c0(1);
   bh7_w92_1_c0 <= tile_16_filtered_output_c0(2);
   bh7_w93_2_c0 <= tile_16_filtered_output_c0(3);
   bh7_w94_2_c0 <= tile_16_filtered_output_c0(4);
   tile_17_X_c0 <= X(52 downto 51);
   tile_17_Y_c0 <= Y(38 downto 36);
   tile_17_mult: IntMultiplierLUT_2x3_Freq300_uid76
      port map ( clk  => clk,
                 X => tile_17_X_c0,
                 Y => tile_17_Y_c0,
                 R => tile_17_output_c0);

   tile_17_filtered_output_c0 <= unsigned(tile_17_output_c0(4 downto 0));
   bh7_w87_1_c0 <= tile_17_filtered_output_c0(0);
   bh7_w88_1_c0 <= tile_17_filtered_output_c0(1);
   bh7_w89_1_c0 <= tile_17_filtered_output_c0(2);
   bh7_w90_2_c0 <= tile_17_filtered_output_c0(3);
   bh7_w91_2_c0 <= tile_17_filtered_output_c0(4);
   tile_18_X_c0 <= X(52 downto 51);
   tile_18_Y_c0 <= Y(35 downto 33);
   tile_18_mult: IntMultiplierLUT_2x3_Freq300_uid81
      port map ( clk  => clk,
                 X => tile_18_X_c0,
                 Y => tile_18_Y_c0,
                 R => tile_18_output_c0);

   tile_18_filtered_output_c0 <= unsigned(tile_18_output_c0(4 downto 0));
   bh7_w84_1_c0 <= tile_18_filtered_output_c0(0);
   bh7_w85_1_c0 <= tile_18_filtered_output_c0(1);
   bh7_w86_1_c0 <= tile_18_filtered_output_c0(2);
   bh7_w87_2_c0 <= tile_18_filtered_output_c0(3);
   bh7_w88_2_c0 <= tile_18_filtered_output_c0(4);
   tile_19_X_c0 <= X(52 downto 51);
   tile_19_Y_c0 <= Y(32 downto 30);
   tile_19_mult: IntMultiplierLUT_2x3_Freq300_uid86
      port map ( clk  => clk,
                 X => tile_19_X_c0,
                 Y => tile_19_Y_c0,
                 R => tile_19_output_c0);

   tile_19_filtered_output_c0 <= unsigned(tile_19_output_c0(4 downto 0));
   bh7_w81_2_c0 <= tile_19_filtered_output_c0(0);
   bh7_w82_1_c0 <= tile_19_filtered_output_c0(1);
   bh7_w83_1_c0 <= tile_19_filtered_output_c0(2);
   bh7_w84_2_c0 <= tile_19_filtered_output_c0(3);
   bh7_w85_2_c0 <= tile_19_filtered_output_c0(4);
   tile_20_X_c0 <= X(52 downto 51);
   tile_20_Y_c0 <= Y(29 downto 27);
   tile_20_mult: IntMultiplierLUT_2x3_Freq300_uid91
      port map ( clk  => clk,
                 X => tile_20_X_c0,
                 Y => tile_20_Y_c0,
                 R => tile_20_output_c0);

   tile_20_filtered_output_c0 <= unsigned(tile_20_output_c0(4 downto 0));
   bh7_w78_2_c0 <= tile_20_filtered_output_c0(0);
   bh7_w79_2_c0 <= tile_20_filtered_output_c0(1);
   bh7_w80_2_c0 <= tile_20_filtered_output_c0(2);
   bh7_w81_3_c0 <= tile_20_filtered_output_c0(3);
   bh7_w82_2_c0 <= tile_20_filtered_output_c0(4);
   tile_21_X_c0 <= X(52 downto 51);
   tile_21_Y_c0 <= Y(26 downto 24);
   tile_21_mult: IntMultiplierLUT_2x3_Freq300_uid96
      port map ( clk  => clk,
                 X => tile_21_X_c0,
                 Y => tile_21_Y_c0,
                 R => tile_21_output_c0);

   tile_21_filtered_output_c0 <= unsigned(tile_21_output_c0(4 downto 0));
   bh7_w75_3_c0 <= tile_21_filtered_output_c0(0);
   bh7_w76_3_c0 <= tile_21_filtered_output_c0(1);
   bh7_w77_2_c0 <= tile_21_filtered_output_c0(2);
   bh7_w78_3_c0 <= tile_21_filtered_output_c0(3);
   bh7_w79_3_c0 <= tile_21_filtered_output_c0(4);
   tile_22_X_c0 <= X(16 downto 16);
   tile_22_Y_c0 <= Y(52 downto 52);
   tile_22_mult: IntMultiplierLUT_1x1_Freq300_uid101
      port map ( clk  => clk,
                 X => tile_22_X_c0,
                 Y => tile_22_Y_c0,
                 R => tile_22_output_c0);

   tile_22_filtered_output_c0 <= unsigned(tile_22_output_c0(0 downto 0));
   bh7_w68_4_c0 <= tile_22_filtered_output_c0(0);
   tile_23_X_c0 <= X(15 downto 12);
   tile_23_Y_c0 <= Y(52 downto 52);
   tile_23_mult: IntMultiplierLUT_4x1_Freq300_uid103
      port map ( clk  => clk,
                 X => tile_23_X_c0,
                 Y => tile_23_Y_c0,
                 R => tile_23_output_c0);

   tile_23_filtered_output_c0 <= unsigned(tile_23_output_c0(3 downto 0));
   bh7_w64_6_c0 <= tile_23_filtered_output_c0(0);
   bh7_w65_4_c0 <= tile_23_filtered_output_c0(1);
   bh7_w66_5_c0 <= tile_23_filtered_output_c0(2);
   bh7_w67_5_c0 <= tile_23_filtered_output_c0(3);
   tile_24_X_c0 <= X(11 downto 8);
   tile_24_Y_c0 <= Y(52 downto 52);
   tile_24_mult: IntMultiplierLUT_4x1_Freq300_uid105
      port map ( clk  => clk,
                 X => tile_24_X_c0,
                 Y => tile_24_Y_c0,
                 R => tile_24_output_c0);

   tile_24_filtered_output_c0 <= unsigned(tile_24_output_c0(3 downto 0));
   bh7_w60_6_c0 <= tile_24_filtered_output_c0(0);
   bh7_w61_6_c0 <= tile_24_filtered_output_c0(1);
   bh7_w62_5_c0 <= tile_24_filtered_output_c0(2);
   bh7_w63_6_c0 <= tile_24_filtered_output_c0(3);
   tile_25_X_c0 <= X(7 downto 4);
   tile_25_Y_c0 <= Y(52 downto 52);
   tile_25_mult: IntMultiplierLUT_4x1_Freq300_uid107
      port map ( clk  => clk,
                 X => tile_25_X_c0,
                 Y => tile_25_Y_c0,
                 R => tile_25_output_c0);

   tile_25_filtered_output_c0 <= unsigned(tile_25_output_c0(3 downto 0));
   bh7_w56_5_c0 <= tile_25_filtered_output_c0(0);
   bh7_w57_6_c0 <= tile_25_filtered_output_c0(1);
   bh7_w58_6_c0 <= tile_25_filtered_output_c0(2);
   bh7_w59_5_c0 <= tile_25_filtered_output_c0(3);
   tile_26_X_c0 <= X(3 downto 0);
   tile_26_Y_c0 <= Y(52 downto 52);
   tile_26_mult: IntMultiplierLUT_4x1_Freq300_uid109
      port map ( clk  => clk,
                 X => tile_26_X_c0,
                 Y => tile_26_Y_c0,
                 R => tile_26_output_c0);

   tile_26_filtered_output_c0 <= unsigned(tile_26_output_c0(3 downto 0));
   bh7_w52_5_c0 <= tile_26_filtered_output_c0(0);
   bh7_w53_5_c0 <= tile_26_filtered_output_c0(1);
   bh7_w54_6_c0 <= tile_26_filtered_output_c0(2);
   bh7_w55_6_c0 <= tile_26_filtered_output_c0(3);
   tile_27_X_c0 <= X(16 downto 15);
   tile_27_Y_c0 <= Y(51 downto 50);
   tile_27_mult: IntMultiplierLUT_2x2_Freq300_uid111
      port map ( clk  => clk,
                 X => tile_27_X_c0,
                 Y => tile_27_Y_c0,
                 R => tile_27_output_c0);

   tile_27_filtered_output_c0 <= unsigned(tile_27_output_c0(3 downto 0));
   bh7_w65_5_c0 <= tile_27_filtered_output_c0(0);
   bh7_w66_6_c0 <= tile_27_filtered_output_c0(1);
   bh7_w67_6_c0 <= tile_27_filtered_output_c0(2);
   bh7_w68_5_c0 <= tile_27_filtered_output_c0(3);
   tile_28_X_c0 <= X(14 downto 12);
   tile_28_Y_c0 <= Y(51 downto 50);
   tile_28_mult: IntMultiplierLUT_3x2_Freq300_uid116
      port map ( clk  => clk,
                 X => tile_28_X_c0,
                 Y => tile_28_Y_c0,
                 R => tile_28_output_c0);

   tile_28_filtered_output_c0 <= unsigned(tile_28_output_c0(4 downto 0));
   bh7_w62_6_c0 <= tile_28_filtered_output_c0(0);
   bh7_w63_7_c0 <= tile_28_filtered_output_c0(1);
   bh7_w64_7_c0 <= tile_28_filtered_output_c0(2);
   bh7_w65_6_c0 <= tile_28_filtered_output_c0(3);
   bh7_w66_7_c0 <= tile_28_filtered_output_c0(4);
   tile_29_X_c0 <= X(11 downto 9);
   tile_29_Y_c0 <= Y(51 downto 50);
   tile_29_mult: IntMultiplierLUT_3x2_Freq300_uid121
      port map ( clk  => clk,
                 X => tile_29_X_c0,
                 Y => tile_29_Y_c0,
                 R => tile_29_output_c0);

   tile_29_filtered_output_c0 <= unsigned(tile_29_output_c0(4 downto 0));
   bh7_w59_6_c0 <= tile_29_filtered_output_c0(0);
   bh7_w60_7_c0 <= tile_29_filtered_output_c0(1);
   bh7_w61_7_c0 <= tile_29_filtered_output_c0(2);
   bh7_w62_7_c0 <= tile_29_filtered_output_c0(3);
   bh7_w63_8_c0 <= tile_29_filtered_output_c0(4);
   tile_30_X_c0 <= X(8 downto 6);
   tile_30_Y_c0 <= Y(51 downto 50);
   tile_30_mult: IntMultiplierLUT_3x2_Freq300_uid126
      port map ( clk  => clk,
                 X => tile_30_X_c0,
                 Y => tile_30_Y_c0,
                 R => tile_30_output_c0);

   tile_30_filtered_output_c0 <= unsigned(tile_30_output_c0(4 downto 0));
   bh7_w56_6_c0 <= tile_30_filtered_output_c0(0);
   bh7_w57_7_c0 <= tile_30_filtered_output_c0(1);
   bh7_w58_7_c0 <= tile_30_filtered_output_c0(2);
   bh7_w59_7_c0 <= tile_30_filtered_output_c0(3);
   bh7_w60_8_c0 <= tile_30_filtered_output_c0(4);
   tile_31_X_c0 <= X(5 downto 3);
   tile_31_Y_c0 <= Y(51 downto 50);
   tile_31_mult: IntMultiplierLUT_3x2_Freq300_uid131
      port map ( clk  => clk,
                 X => tile_31_X_c0,
                 Y => tile_31_Y_c0,
                 R => tile_31_output_c0);

   tile_31_filtered_output_c0 <= unsigned(tile_31_output_c0(4 downto 0));
   bh7_w53_6_c0 <= tile_31_filtered_output_c0(0);
   bh7_w54_7_c0 <= tile_31_filtered_output_c0(1);
   bh7_w55_7_c0 <= tile_31_filtered_output_c0(2);
   bh7_w56_7_c0 <= tile_31_filtered_output_c0(3);
   bh7_w57_8_c0 <= tile_31_filtered_output_c0(4);
   tile_32_X_c0 <= X(2 downto 0);
   tile_32_Y_c0 <= Y(51 downto 50);
   tile_32_mult: IntMultiplierLUT_3x2_Freq300_uid136
      port map ( clk  => clk,
                 X => tile_32_X_c0,
                 Y => tile_32_Y_c0,
                 R => tile_32_output_c0);

   tile_32_filtered_output_c0 <= unsigned(tile_32_output_c0(4 downto 0));
   bh7_w50_4_c0 <= tile_32_filtered_output_c0(0);
   bh7_w51_5_c0 <= tile_32_filtered_output_c0(1);
   bh7_w52_6_c0 <= tile_32_filtered_output_c0(2);
   bh7_w53_7_c0 <= tile_32_filtered_output_c0(3);
   bh7_w54_8_c0 <= tile_32_filtered_output_c0(4);
   tile_33_X_c0 <= X(16 downto 15);
   tile_33_Y_c0 <= Y(49 downto 48);
   tile_33_mult: IntMultiplierLUT_2x2_Freq300_uid141
      port map ( clk  => clk,
                 X => tile_33_X_c0,
                 Y => tile_33_Y_c0,
                 R => tile_33_output_c0);

   tile_33_filtered_output_c0 <= unsigned(tile_33_output_c0(3 downto 0));
   bh7_w63_9_c0 <= tile_33_filtered_output_c0(0);
   bh7_w64_8_c0 <= tile_33_filtered_output_c0(1);
   bh7_w65_7_c0 <= tile_33_filtered_output_c0(2);
   bh7_w66_8_c0 <= tile_33_filtered_output_c0(3);
   tile_34_X_c0 <= X(14 downto 12);
   tile_34_Y_c0 <= Y(49 downto 48);
   tile_34_mult: IntMultiplierLUT_3x2_Freq300_uid146
      port map ( clk  => clk,
                 X => tile_34_X_c0,
                 Y => tile_34_Y_c0,
                 R => tile_34_output_c0);

   tile_34_filtered_output_c0 <= unsigned(tile_34_output_c0(4 downto 0));
   bh7_w60_9_c0 <= tile_34_filtered_output_c0(0);
   bh7_w61_8_c0 <= tile_34_filtered_output_c0(1);
   bh7_w62_8_c0 <= tile_34_filtered_output_c0(2);
   bh7_w63_10_c0 <= tile_34_filtered_output_c0(3);
   bh7_w64_9_c0 <= tile_34_filtered_output_c0(4);
   tile_35_X_c0 <= X(11 downto 9);
   tile_35_Y_c0 <= Y(49 downto 48);
   tile_35_mult: IntMultiplierLUT_3x2_Freq300_uid151
      port map ( clk  => clk,
                 X => tile_35_X_c0,
                 Y => tile_35_Y_c0,
                 R => tile_35_output_c0);

   tile_35_filtered_output_c0 <= unsigned(tile_35_output_c0(4 downto 0));
   bh7_w57_9_c0 <= tile_35_filtered_output_c0(0);
   bh7_w58_8_c0 <= tile_35_filtered_output_c0(1);
   bh7_w59_8_c0 <= tile_35_filtered_output_c0(2);
   bh7_w60_10_c0 <= tile_35_filtered_output_c0(3);
   bh7_w61_9_c0 <= tile_35_filtered_output_c0(4);
   tile_36_X_c0 <= X(8 downto 6);
   tile_36_Y_c0 <= Y(49 downto 48);
   tile_36_mult: IntMultiplierLUT_3x2_Freq300_uid156
      port map ( clk  => clk,
                 X => tile_36_X_c0,
                 Y => tile_36_Y_c0,
                 R => tile_36_output_c0);

   tile_36_filtered_output_c0 <= unsigned(tile_36_output_c0(4 downto 0));
   bh7_w54_9_c0 <= tile_36_filtered_output_c0(0);
   bh7_w55_8_c0 <= tile_36_filtered_output_c0(1);
   bh7_w56_8_c0 <= tile_36_filtered_output_c0(2);
   bh7_w57_10_c0 <= tile_36_filtered_output_c0(3);
   bh7_w58_9_c0 <= tile_36_filtered_output_c0(4);
   tile_37_X_c0 <= X(5 downto 3);
   tile_37_Y_c0 <= Y(49 downto 48);
   tile_37_mult: IntMultiplierLUT_3x2_Freq300_uid161
      port map ( clk  => clk,
                 X => tile_37_X_c0,
                 Y => tile_37_Y_c0,
                 R => tile_37_output_c0);

   tile_37_filtered_output_c0 <= unsigned(tile_37_output_c0(4 downto 0));
   bh7_w51_6_c0 <= tile_37_filtered_output_c0(0);
   bh7_w52_7_c0 <= tile_37_filtered_output_c0(1);
   bh7_w53_8_c0 <= tile_37_filtered_output_c0(2);
   bh7_w54_10_c0 <= tile_37_filtered_output_c0(3);
   bh7_w55_9_c0 <= tile_37_filtered_output_c0(4);
   tile_38_X_c0 <= X(2 downto 0);
   tile_38_Y_c0 <= Y(49 downto 48);
   tile_38_mult: IntMultiplierLUT_3x2_Freq300_uid166
      port map ( clk  => clk,
                 X => tile_38_X_c0,
                 Y => tile_38_Y_c0,
                 R => tile_38_output_c0);

   tile_38_filtered_output_c0 <= unsigned(tile_38_output_c0(4 downto 0));
   bh7_w48_4_c0 <= tile_38_filtered_output_c0(0);
   bh7_w49_4_c0 <= tile_38_filtered_output_c0(1);
   bh7_w50_5_c0 <= tile_38_filtered_output_c0(2);
   bh7_w51_7_c0 <= tile_38_filtered_output_c0(3);
   bh7_w52_8_c0 <= tile_38_filtered_output_c0(4);
   tile_39_X_c0 <= X(33 downto 33);
   tile_39_Y_c0 <= Y(52 downto 52);
   tile_39_mult: IntMultiplierLUT_1x1_Freq300_uid171
      port map ( clk  => clk,
                 X => tile_39_X_c0,
                 Y => tile_39_Y_c0,
                 R => tile_39_output_c0);

   tile_39_filtered_output_c0 <= unsigned(tile_39_output_c0(0 downto 0));
   bh7_w85_3_c0 <= tile_39_filtered_output_c0(0);
   tile_40_X_c0 <= X(32 downto 29);
   tile_40_Y_c0 <= Y(52 downto 52);
   tile_40_mult: IntMultiplierLUT_4x1_Freq300_uid173
      port map ( clk  => clk,
                 X => tile_40_X_c0,
                 Y => tile_40_Y_c0,
                 R => tile_40_output_c0);

   tile_40_filtered_output_c0 <= unsigned(tile_40_output_c0(3 downto 0));
   bh7_w81_4_c0 <= tile_40_filtered_output_c0(0);
   bh7_w82_3_c0 <= tile_40_filtered_output_c0(1);
   bh7_w83_2_c0 <= tile_40_filtered_output_c0(2);
   bh7_w84_3_c0 <= tile_40_filtered_output_c0(3);
   tile_41_X_c0 <= X(28 downto 25);
   tile_41_Y_c0 <= Y(52 downto 52);
   tile_41_mult: IntMultiplierLUT_4x1_Freq300_uid175
      port map ( clk  => clk,
                 X => tile_41_X_c0,
                 Y => tile_41_Y_c0,
                 R => tile_41_output_c0);

   tile_41_filtered_output_c0 <= unsigned(tile_41_output_c0(3 downto 0));
   bh7_w77_3_c0 <= tile_41_filtered_output_c0(0);
   bh7_w78_4_c0 <= tile_41_filtered_output_c0(1);
   bh7_w79_4_c0 <= tile_41_filtered_output_c0(2);
   bh7_w80_3_c0 <= tile_41_filtered_output_c0(3);
   tile_42_X_c0 <= X(24 downto 21);
   tile_42_Y_c0 <= Y(52 downto 52);
   tile_42_mult: IntMultiplierLUT_4x1_Freq300_uid177
      port map ( clk  => clk,
                 X => tile_42_X_c0,
                 Y => tile_42_Y_c0,
                 R => tile_42_output_c0);

   tile_42_filtered_output_c0 <= unsigned(tile_42_output_c0(3 downto 0));
   bh7_w73_5_c0 <= tile_42_filtered_output_c0(0);
   bh7_w74_4_c0 <= tile_42_filtered_output_c0(1);
   bh7_w75_4_c0 <= tile_42_filtered_output_c0(2);
   bh7_w76_4_c0 <= tile_42_filtered_output_c0(3);
   tile_43_X_c0 <= X(20 downto 17);
   tile_43_Y_c0 <= Y(52 downto 52);
   tile_43_mult: IntMultiplierLUT_4x1_Freq300_uid179
      port map ( clk  => clk,
                 X => tile_43_X_c0,
                 Y => tile_43_Y_c0,
                 R => tile_43_output_c0);

   tile_43_filtered_output_c0 <= unsigned(tile_43_output_c0(3 downto 0));
   bh7_w69_5_c0 <= tile_43_filtered_output_c0(0);
   bh7_w70_5_c0 <= tile_43_filtered_output_c0(1);
   bh7_w71_4_c0 <= tile_43_filtered_output_c0(2);
   bh7_w72_5_c0 <= tile_43_filtered_output_c0(3);
   tile_44_X_c0 <= X(33 downto 32);
   tile_44_Y_c0 <= Y(51 downto 50);
   tile_44_mult: IntMultiplierLUT_2x2_Freq300_uid181
      port map ( clk  => clk,
                 X => tile_44_X_c0,
                 Y => tile_44_Y_c0,
                 R => tile_44_output_c0);

   tile_44_filtered_output_c0 <= unsigned(tile_44_output_c0(3 downto 0));
   bh7_w82_4_c0 <= tile_44_filtered_output_c0(0);
   bh7_w83_3_c0 <= tile_44_filtered_output_c0(1);
   bh7_w84_4_c0 <= tile_44_filtered_output_c0(2);
   bh7_w85_4_c0 <= tile_44_filtered_output_c0(3);
   tile_45_X_c0 <= X(31 downto 29);
   tile_45_Y_c0 <= Y(51 downto 50);
   tile_45_mult: IntMultiplierLUT_3x2_Freq300_uid186
      port map ( clk  => clk,
                 X => tile_45_X_c0,
                 Y => tile_45_Y_c0,
                 R => tile_45_output_c0);

   tile_45_filtered_output_c0 <= unsigned(tile_45_output_c0(4 downto 0));
   bh7_w79_5_c0 <= tile_45_filtered_output_c0(0);
   bh7_w80_4_c0 <= tile_45_filtered_output_c0(1);
   bh7_w81_5_c0 <= tile_45_filtered_output_c0(2);
   bh7_w82_5_c0 <= tile_45_filtered_output_c0(3);
   bh7_w83_4_c0 <= tile_45_filtered_output_c0(4);
   tile_46_X_c0 <= X(28 downto 26);
   tile_46_Y_c0 <= Y(51 downto 50);
   tile_46_mult: IntMultiplierLUT_3x2_Freq300_uid191
      port map ( clk  => clk,
                 X => tile_46_X_c0,
                 Y => tile_46_Y_c0,
                 R => tile_46_output_c0);

   tile_46_filtered_output_c0 <= unsigned(tile_46_output_c0(4 downto 0));
   bh7_w76_5_c0 <= tile_46_filtered_output_c0(0);
   bh7_w77_4_c0 <= tile_46_filtered_output_c0(1);
   bh7_w78_5_c0 <= tile_46_filtered_output_c0(2);
   bh7_w79_6_c0 <= tile_46_filtered_output_c0(3);
   bh7_w80_5_c0 <= tile_46_filtered_output_c0(4);
   tile_47_X_c0 <= X(25 downto 23);
   tile_47_Y_c0 <= Y(51 downto 50);
   tile_47_mult: IntMultiplierLUT_3x2_Freq300_uid196
      port map ( clk  => clk,
                 X => tile_47_X_c0,
                 Y => tile_47_Y_c0,
                 R => tile_47_output_c0);

   tile_47_filtered_output_c0 <= unsigned(tile_47_output_c0(4 downto 0));
   bh7_w73_6_c0 <= tile_47_filtered_output_c0(0);
   bh7_w74_5_c0 <= tile_47_filtered_output_c0(1);
   bh7_w75_5_c0 <= tile_47_filtered_output_c0(2);
   bh7_w76_6_c0 <= tile_47_filtered_output_c0(3);
   bh7_w77_5_c0 <= tile_47_filtered_output_c0(4);
   tile_48_X_c0 <= X(22 downto 20);
   tile_48_Y_c0 <= Y(51 downto 50);
   tile_48_mult: IntMultiplierLUT_3x2_Freq300_uid201
      port map ( clk  => clk,
                 X => tile_48_X_c0,
                 Y => tile_48_Y_c0,
                 R => tile_48_output_c0);

   tile_48_filtered_output_c0 <= unsigned(tile_48_output_c0(4 downto 0));
   bh7_w70_6_c0 <= tile_48_filtered_output_c0(0);
   bh7_w71_5_c0 <= tile_48_filtered_output_c0(1);
   bh7_w72_6_c0 <= tile_48_filtered_output_c0(2);
   bh7_w73_7_c0 <= tile_48_filtered_output_c0(3);
   bh7_w74_6_c0 <= tile_48_filtered_output_c0(4);
   tile_49_X_c0 <= X(19 downto 17);
   tile_49_Y_c0 <= Y(51 downto 50);
   tile_49_mult: IntMultiplierLUT_3x2_Freq300_uid206
      port map ( clk  => clk,
                 X => tile_49_X_c0,
                 Y => tile_49_Y_c0,
                 R => tile_49_output_c0);

   tile_49_filtered_output_c0 <= unsigned(tile_49_output_c0(4 downto 0));
   bh7_w67_7_c0 <= tile_49_filtered_output_c0(0);
   bh7_w68_6_c0 <= tile_49_filtered_output_c0(1);
   bh7_w69_6_c0 <= tile_49_filtered_output_c0(2);
   bh7_w70_7_c0 <= tile_49_filtered_output_c0(3);
   bh7_w71_6_c0 <= tile_49_filtered_output_c0(4);
   tile_50_X_c0 <= X(33 downto 32);
   tile_50_Y_c0 <= Y(49 downto 48);
   tile_50_mult: IntMultiplierLUT_2x2_Freq300_uid211
      port map ( clk  => clk,
                 X => tile_50_X_c0,
                 Y => tile_50_Y_c0,
                 R => tile_50_output_c0);

   tile_50_filtered_output_c0 <= unsigned(tile_50_output_c0(3 downto 0));
   bh7_w80_6_c0 <= tile_50_filtered_output_c0(0);
   bh7_w81_6_c0 <= tile_50_filtered_output_c0(1);
   bh7_w82_6_c0 <= tile_50_filtered_output_c0(2);
   bh7_w83_5_c0 <= tile_50_filtered_output_c0(3);
   tile_51_X_c0 <= X(31 downto 29);
   tile_51_Y_c0 <= Y(49 downto 48);
   tile_51_mult: IntMultiplierLUT_3x2_Freq300_uid216
      port map ( clk  => clk,
                 X => tile_51_X_c0,
                 Y => tile_51_Y_c0,
                 R => tile_51_output_c0);

   tile_51_filtered_output_c0 <= unsigned(tile_51_output_c0(4 downto 0));
   bh7_w77_6_c0 <= tile_51_filtered_output_c0(0);
   bh7_w78_6_c0 <= tile_51_filtered_output_c0(1);
   bh7_w79_7_c0 <= tile_51_filtered_output_c0(2);
   bh7_w80_7_c0 <= tile_51_filtered_output_c0(3);
   bh7_w81_7_c0 <= tile_51_filtered_output_c0(4);
   tile_52_X_c0 <= X(28 downto 26);
   tile_52_Y_c0 <= Y(49 downto 48);
   tile_52_mult: IntMultiplierLUT_3x2_Freq300_uid221
      port map ( clk  => clk,
                 X => tile_52_X_c0,
                 Y => tile_52_Y_c0,
                 R => tile_52_output_c0);

   tile_52_filtered_output_c0 <= unsigned(tile_52_output_c0(4 downto 0));
   bh7_w74_7_c0 <= tile_52_filtered_output_c0(0);
   bh7_w75_6_c0 <= tile_52_filtered_output_c0(1);
   bh7_w76_7_c0 <= tile_52_filtered_output_c0(2);
   bh7_w77_7_c0 <= tile_52_filtered_output_c0(3);
   bh7_w78_7_c0 <= tile_52_filtered_output_c0(4);
   tile_53_X_c0 <= X(25 downto 23);
   tile_53_Y_c0 <= Y(49 downto 48);
   tile_53_mult: IntMultiplierLUT_3x2_Freq300_uid226
      port map ( clk  => clk,
                 X => tile_53_X_c0,
                 Y => tile_53_Y_c0,
                 R => tile_53_output_c0);

   tile_53_filtered_output_c0 <= unsigned(tile_53_output_c0(4 downto 0));
   bh7_w71_7_c0 <= tile_53_filtered_output_c0(0);
   bh7_w72_7_c0 <= tile_53_filtered_output_c0(1);
   bh7_w73_8_c0 <= tile_53_filtered_output_c0(2);
   bh7_w74_8_c0 <= tile_53_filtered_output_c0(3);
   bh7_w75_7_c0 <= tile_53_filtered_output_c0(4);
   tile_54_X_c0 <= X(22 downto 20);
   tile_54_Y_c0 <= Y(49 downto 48);
   tile_54_mult: IntMultiplierLUT_3x2_Freq300_uid231
      port map ( clk  => clk,
                 X => tile_54_X_c0,
                 Y => tile_54_Y_c0,
                 R => tile_54_output_c0);

   tile_54_filtered_output_c0 <= unsigned(tile_54_output_c0(4 downto 0));
   bh7_w68_7_c0 <= tile_54_filtered_output_c0(0);
   bh7_w69_7_c0 <= tile_54_filtered_output_c0(1);
   bh7_w70_8_c0 <= tile_54_filtered_output_c0(2);
   bh7_w71_8_c0 <= tile_54_filtered_output_c0(3);
   bh7_w72_8_c0 <= tile_54_filtered_output_c0(4);
   tile_55_X_c0 <= X(19 downto 17);
   tile_55_Y_c0 <= Y(49 downto 48);
   tile_55_mult: IntMultiplierLUT_3x2_Freq300_uid236
      port map ( clk  => clk,
                 X => tile_55_X_c0,
                 Y => tile_55_Y_c0,
                 R => tile_55_output_c0);

   tile_55_filtered_output_c0 <= unsigned(tile_55_output_c0(4 downto 0));
   bh7_w65_8_c0 <= tile_55_filtered_output_c0(0);
   bh7_w66_9_c0 <= tile_55_filtered_output_c0(1);
   bh7_w67_8_c0 <= tile_55_filtered_output_c0(2);
   bh7_w68_8_c0 <= tile_55_filtered_output_c0(3);
   bh7_w69_8_c0 <= tile_55_filtered_output_c0(4);
   tile_56_X_c0 <= X(50 downto 50);
   tile_56_Y_c0 <= Y(52 downto 52);
   tile_56_mult: IntMultiplierLUT_1x1_Freq300_uid241
      port map ( clk  => clk,
                 X => tile_56_X_c0,
                 Y => tile_56_Y_c0,
                 R => tile_56_output_c0);

   tile_56_filtered_output_c0 <= unsigned(tile_56_output_c0(0 downto 0));
   bh7_w102_0_c0 <= tile_56_filtered_output_c0(0);
   tile_57_X_c0 <= X(49 downto 46);
   tile_57_Y_c0 <= Y(52 downto 52);
   tile_57_mult: IntMultiplierLUT_4x1_Freq300_uid243
      port map ( clk  => clk,
                 X => tile_57_X_c0,
                 Y => tile_57_Y_c0,
                 R => tile_57_output_c0);

   tile_57_filtered_output_c0 <= unsigned(tile_57_output_c0(3 downto 0));
   bh7_w98_2_c0 <= tile_57_filtered_output_c0(0);
   bh7_w99_1_c0 <= tile_57_filtered_output_c0(1);
   bh7_w100_1_c0 <= tile_57_filtered_output_c0(2);
   bh7_w101_0_c0 <= tile_57_filtered_output_c0(3);
   tile_58_X_c0 <= X(45 downto 42);
   tile_58_Y_c0 <= Y(52 downto 52);
   tile_58_mult: IntMultiplierLUT_4x1_Freq300_uid245
      port map ( clk  => clk,
                 X => tile_58_X_c0,
                 Y => tile_58_Y_c0,
                 R => tile_58_output_c0);

   tile_58_filtered_output_c0 <= unsigned(tile_58_output_c0(3 downto 0));
   bh7_w94_3_c0 <= tile_58_filtered_output_c0(0);
   bh7_w95_2_c0 <= tile_58_filtered_output_c0(1);
   bh7_w96_3_c0 <= tile_58_filtered_output_c0(2);
   bh7_w97_3_c0 <= tile_58_filtered_output_c0(3);
   tile_59_X_c0 <= X(41 downto 38);
   tile_59_Y_c0 <= Y(52 downto 52);
   tile_59_mult: IntMultiplierLUT_4x1_Freq300_uid247
      port map ( clk  => clk,
                 X => tile_59_X_c0,
                 Y => tile_59_Y_c0,
                 R => tile_59_output_c0);

   tile_59_filtered_output_c0 <= unsigned(tile_59_output_c0(3 downto 0));
   bh7_w90_3_c0 <= tile_59_filtered_output_c0(0);
   bh7_w91_3_c0 <= tile_59_filtered_output_c0(1);
   bh7_w92_2_c0 <= tile_59_filtered_output_c0(2);
   bh7_w93_3_c0 <= tile_59_filtered_output_c0(3);
   tile_60_X_c0 <= X(37 downto 34);
   tile_60_Y_c0 <= Y(52 downto 52);
   tile_60_mult: IntMultiplierLUT_4x1_Freq300_uid249
      port map ( clk  => clk,
                 X => tile_60_X_c0,
                 Y => tile_60_Y_c0,
                 R => tile_60_output_c0);

   tile_60_filtered_output_c0 <= unsigned(tile_60_output_c0(3 downto 0));
   bh7_w86_2_c0 <= tile_60_filtered_output_c0(0);
   bh7_w87_3_c0 <= tile_60_filtered_output_c0(1);
   bh7_w88_3_c0 <= tile_60_filtered_output_c0(2);
   bh7_w89_2_c0 <= tile_60_filtered_output_c0(3);
   tile_61_X_c0 <= X(50 downto 49);
   tile_61_Y_c0 <= Y(51 downto 50);
   tile_61_mult: IntMultiplierLUT_2x2_Freq300_uid251
      port map ( clk  => clk,
                 X => tile_61_X_c0,
                 Y => tile_61_Y_c0,
                 R => tile_61_output_c0);

   tile_61_filtered_output_c0 <= unsigned(tile_61_output_c0(3 downto 0));
   bh7_w99_2_c0 <= tile_61_filtered_output_c0(0);
   bh7_w100_2_c0 <= tile_61_filtered_output_c0(1);
   bh7_w101_1_c0 <= tile_61_filtered_output_c0(2);
   bh7_w102_1_c0 <= tile_61_filtered_output_c0(3);
   tile_62_X_c0 <= X(48 downto 46);
   tile_62_Y_c0 <= Y(51 downto 50);
   tile_62_mult: IntMultiplierLUT_3x2_Freq300_uid256
      port map ( clk  => clk,
                 X => tile_62_X_c0,
                 Y => tile_62_Y_c0,
                 R => tile_62_output_c0);

   tile_62_filtered_output_c0 <= unsigned(tile_62_output_c0(4 downto 0));
   bh7_w96_4_c0 <= tile_62_filtered_output_c0(0);
   bh7_w97_4_c0 <= tile_62_filtered_output_c0(1);
   bh7_w98_3_c0 <= tile_62_filtered_output_c0(2);
   bh7_w99_3_c0 <= tile_62_filtered_output_c0(3);
   bh7_w100_3_c0 <= tile_62_filtered_output_c0(4);
   tile_63_X_c0 <= X(45 downto 43);
   tile_63_Y_c0 <= Y(51 downto 50);
   tile_63_mult: IntMultiplierLUT_3x2_Freq300_uid261
      port map ( clk  => clk,
                 X => tile_63_X_c0,
                 Y => tile_63_Y_c0,
                 R => tile_63_output_c0);

   tile_63_filtered_output_c0 <= unsigned(tile_63_output_c0(4 downto 0));
   bh7_w93_4_c0 <= tile_63_filtered_output_c0(0);
   bh7_w94_4_c0 <= tile_63_filtered_output_c0(1);
   bh7_w95_3_c0 <= tile_63_filtered_output_c0(2);
   bh7_w96_5_c0 <= tile_63_filtered_output_c0(3);
   bh7_w97_5_c0 <= tile_63_filtered_output_c0(4);
   tile_64_X_c0 <= X(42 downto 40);
   tile_64_Y_c0 <= Y(51 downto 50);
   tile_64_mult: IntMultiplierLUT_3x2_Freq300_uid266
      port map ( clk  => clk,
                 X => tile_64_X_c0,
                 Y => tile_64_Y_c0,
                 R => tile_64_output_c0);

   tile_64_filtered_output_c0 <= unsigned(tile_64_output_c0(4 downto 0));
   bh7_w90_4_c0 <= tile_64_filtered_output_c0(0);
   bh7_w91_4_c0 <= tile_64_filtered_output_c0(1);
   bh7_w92_3_c0 <= tile_64_filtered_output_c0(2);
   bh7_w93_5_c0 <= tile_64_filtered_output_c0(3);
   bh7_w94_5_c0 <= tile_64_filtered_output_c0(4);
   tile_65_X_c0 <= X(39 downto 37);
   tile_65_Y_c0 <= Y(51 downto 50);
   tile_65_mult: IntMultiplierLUT_3x2_Freq300_uid271
      port map ( clk  => clk,
                 X => tile_65_X_c0,
                 Y => tile_65_Y_c0,
                 R => tile_65_output_c0);

   tile_65_filtered_output_c0 <= unsigned(tile_65_output_c0(4 downto 0));
   bh7_w87_4_c0 <= tile_65_filtered_output_c0(0);
   bh7_w88_4_c0 <= tile_65_filtered_output_c0(1);
   bh7_w89_3_c0 <= tile_65_filtered_output_c0(2);
   bh7_w90_5_c0 <= tile_65_filtered_output_c0(3);
   bh7_w91_5_c0 <= tile_65_filtered_output_c0(4);
   tile_66_X_c0 <= X(36 downto 34);
   tile_66_Y_c0 <= Y(51 downto 50);
   tile_66_mult: IntMultiplierLUT_3x2_Freq300_uid276
      port map ( clk  => clk,
                 X => tile_66_X_c0,
                 Y => tile_66_Y_c0,
                 R => tile_66_output_c0);

   tile_66_filtered_output_c0 <= unsigned(tile_66_output_c0(4 downto 0));
   bh7_w84_5_c0 <= tile_66_filtered_output_c0(0);
   bh7_w85_5_c0 <= tile_66_filtered_output_c0(1);
   bh7_w86_3_c0 <= tile_66_filtered_output_c0(2);
   bh7_w87_5_c0 <= tile_66_filtered_output_c0(3);
   bh7_w88_5_c0 <= tile_66_filtered_output_c0(4);
   tile_67_X_c0 <= X(50 downto 49);
   tile_67_Y_c0 <= Y(49 downto 48);
   tile_67_mult: IntMultiplierLUT_2x2_Freq300_uid281
      port map ( clk  => clk,
                 X => tile_67_X_c0,
                 Y => tile_67_Y_c0,
                 R => tile_67_output_c0);

   tile_67_filtered_output_c0 <= unsigned(tile_67_output_c0(3 downto 0));
   bh7_w97_6_c0 <= tile_67_filtered_output_c0(0);
   bh7_w98_4_c0 <= tile_67_filtered_output_c0(1);
   bh7_w99_4_c0 <= tile_67_filtered_output_c0(2);
   bh7_w100_4_c0 <= tile_67_filtered_output_c0(3);
   tile_68_X_c0 <= X(48 downto 46);
   tile_68_Y_c0 <= Y(49 downto 48);
   tile_68_mult: IntMultiplierLUT_3x2_Freq300_uid286
      port map ( clk  => clk,
                 X => tile_68_X_c0,
                 Y => tile_68_Y_c0,
                 R => tile_68_output_c0);

   tile_68_filtered_output_c0 <= unsigned(tile_68_output_c0(4 downto 0));
   bh7_w94_6_c0 <= tile_68_filtered_output_c0(0);
   bh7_w95_4_c0 <= tile_68_filtered_output_c0(1);
   bh7_w96_6_c0 <= tile_68_filtered_output_c0(2);
   bh7_w97_7_c0 <= tile_68_filtered_output_c0(3);
   bh7_w98_5_c0 <= tile_68_filtered_output_c0(4);
   tile_69_X_c0 <= X(45 downto 43);
   tile_69_Y_c0 <= Y(49 downto 48);
   tile_69_mult: IntMultiplierLUT_3x2_Freq300_uid291
      port map ( clk  => clk,
                 X => tile_69_X_c0,
                 Y => tile_69_Y_c0,
                 R => tile_69_output_c0);

   tile_69_filtered_output_c0 <= unsigned(tile_69_output_c0(4 downto 0));
   bh7_w91_6_c0 <= tile_69_filtered_output_c0(0);
   bh7_w92_4_c0 <= tile_69_filtered_output_c0(1);
   bh7_w93_6_c0 <= tile_69_filtered_output_c0(2);
   bh7_w94_7_c0 <= tile_69_filtered_output_c0(3);
   bh7_w95_5_c0 <= tile_69_filtered_output_c0(4);
   tile_70_X_c0 <= X(42 downto 40);
   tile_70_Y_c0 <= Y(49 downto 48);
   tile_70_mult: IntMultiplierLUT_3x2_Freq300_uid296
      port map ( clk  => clk,
                 X => tile_70_X_c0,
                 Y => tile_70_Y_c0,
                 R => tile_70_output_c0);

   tile_70_filtered_output_c0 <= unsigned(tile_70_output_c0(4 downto 0));
   bh7_w88_6_c0 <= tile_70_filtered_output_c0(0);
   bh7_w89_4_c0 <= tile_70_filtered_output_c0(1);
   bh7_w90_6_c0 <= tile_70_filtered_output_c0(2);
   bh7_w91_7_c0 <= tile_70_filtered_output_c0(3);
   bh7_w92_5_c0 <= tile_70_filtered_output_c0(4);
   tile_71_X_c0 <= X(39 downto 37);
   tile_71_Y_c0 <= Y(49 downto 48);
   tile_71_mult: IntMultiplierLUT_3x2_Freq300_uid301
      port map ( clk  => clk,
                 X => tile_71_X_c0,
                 Y => tile_71_Y_c0,
                 R => tile_71_output_c0);

   tile_71_filtered_output_c0 <= unsigned(tile_71_output_c0(4 downto 0));
   bh7_w85_6_c0 <= tile_71_filtered_output_c0(0);
   bh7_w86_4_c0 <= tile_71_filtered_output_c0(1);
   bh7_w87_6_c0 <= tile_71_filtered_output_c0(2);
   bh7_w88_7_c0 <= tile_71_filtered_output_c0(3);
   bh7_w89_5_c0 <= tile_71_filtered_output_c0(4);
   tile_72_X_c0 <= X(36 downto 34);
   tile_72_Y_c0 <= Y(49 downto 48);
   tile_72_mult: IntMultiplierLUT_3x2_Freq300_uid306
      port map ( clk  => clk,
                 X => tile_72_X_c0,
                 Y => tile_72_Y_c0,
                 R => tile_72_output_c0);

   tile_72_filtered_output_c0 <= unsigned(tile_72_output_c0(4 downto 0));
   bh7_w82_7_c0 <= tile_72_filtered_output_c0(0);
   bh7_w83_6_c0 <= tile_72_filtered_output_c0(1);
   bh7_w84_6_c0 <= tile_72_filtered_output_c0(2);
   bh7_w85_7_c0 <= tile_72_filtered_output_c0(3);
   bh7_w86_5_c0 <= tile_72_filtered_output_c0(4);
   tile_73_X_c0 <= X(52 downto 51);
   tile_73_Y_c0 <= Y(52 downto 51);
   tile_73_mult: IntMultiplierLUT_2x2_Freq300_uid311
      port map ( clk  => clk,
                 X => tile_73_X_c0,
                 Y => tile_73_Y_c0,
                 R => tile_73_output_c0);

   tile_73_filtered_output_c0 <= unsigned(tile_73_output_c0(3 downto 0));
   bh7_w102_2_c0 <= tile_73_filtered_output_c0(0);
   bh7_w103_0_c0 <= tile_73_filtered_output_c0(1);
   bh7_w104_0_c0 <= tile_73_filtered_output_c0(2);
   bh7_w105_0_c0 <= tile_73_filtered_output_c0(3);
   tile_74_X_c0 <= X(52 downto 51);
   tile_74_Y_c0 <= Y(50 downto 48);
   tile_74_mult: IntMultiplierLUT_2x3_Freq300_uid316
      port map ( clk  => clk,
                 X => tile_74_X_c0,
                 Y => tile_74_Y_c0,
                 R => tile_74_output_c0);

   tile_74_filtered_output_c0 <= unsigned(tile_74_output_c0(4 downto 0));
   bh7_w99_5_c0 <= tile_74_filtered_output_c0(0);
   bh7_w100_5_c0 <= tile_74_filtered_output_c0(1);
   bh7_w101_2_c0 <= tile_74_filtered_output_c0(2);
   bh7_w102_3_c0 <= tile_74_filtered_output_c0(3);
   bh7_w103_1_c0 <= tile_74_filtered_output_c0(4);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq300_uid322_bh7_uid323_In0_c0 <= "" & bh7_w49_4_c0 & "0" & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid323_In1_c0 <= "" & bh7_w50_4_c0 & bh7_w50_5_c0;
   bh7_w49_5_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0(0);
   bh7_w50_6_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0(1);
   bh7_w51_8_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid323: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid323_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid323_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_copy324_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid323_Out0_copy324_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid327_In0_c0 <= "" & bh7_w51_2_c0 & bh7_w51_5_c0 & bh7_w51_6_c0 & bh7_w51_7_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid327_In1_c0 <= "" & bh7_w52_2_c0;
   bh7_w51_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0(0);
   bh7_w52_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0(1);
   bh7_w53_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid327: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid327_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid327_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_copy328_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid327_Out0_copy328_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid329_In0_c0 <= "" & bh7_w52_5_c0 & bh7_w52_6_c0 & bh7_w52_7_c0 & bh7_w52_8_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid329_In1_c0 <= "" & bh7_w53_2_c0;
   bh7_w52_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0(0);
   bh7_w53_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0(1);
   bh7_w54_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid329: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid329_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid329_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_copy330_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid329_Out0_copy330_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid331_In0_c0 <= "" & bh7_w53_5_c0 & bh7_w53_6_c0 & bh7_w53_7_c0 & bh7_w53_8_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid331_In1_c0 <= "" & bh7_w54_2_c0;
   bh7_w53_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0(0);
   bh7_w54_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0(1);
   bh7_w55_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid331: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid331_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid331_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_copy332_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid331_Out0_copy332_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid335_In0_c0 <= "" & bh7_w54_3_c0 & bh7_w54_6_c0 & bh7_w54_7_c0 & bh7_w54_8_c0 & bh7_w54_9_c0 & bh7_w54_10_c0;
   bh7_w54_13_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0(0);
   bh7_w55_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0(1);
   bh7_w56_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid335: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid335_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_copy336_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid335_Out0_copy336_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid337_In0_c0 <= "" & bh7_w55_2_c0 & bh7_w55_3_c0 & bh7_w55_6_c0 & bh7_w55_7_c0 & bh7_w55_8_c0 & bh7_w55_9_c0;
   bh7_w55_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0(0);
   bh7_w56_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0(1);
   bh7_w57_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid337: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid337_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_copy338_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid337_Out0_copy338_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid339_In0_c0 <= "" & bh7_w56_2_c0 & bh7_w56_5_c0 & bh7_w56_6_c0 & bh7_w56_7_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid339_In1_c0 <= "" & bh7_w57_2_c0;
   bh7_w56_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0(0);
   bh7_w57_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0(1);
   bh7_w58_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid339: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid339_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid339_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_copy340_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid339_Out0_copy340_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid341_In0_c0 <= "" & bh7_w57_3_c0 & bh7_w57_6_c0 & bh7_w57_7_c0 & bh7_w57_8_c0 & bh7_w57_9_c0 & bh7_w57_10_c0;
   bh7_w57_13_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0(0);
   bh7_w58_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0(1);
   bh7_w59_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid341: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid341_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_copy342_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid341_Out0_copy342_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid343_In0_c0 <= "" & bh7_w58_1_c0 & bh7_w58_2_c0 & bh7_w58_6_c0 & bh7_w58_7_c0 & bh7_w58_8_c0 & bh7_w58_9_c0;
   bh7_w58_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0(0);
   bh7_w59_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0(1);
   bh7_w60_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid343: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid343_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_copy344_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid343_Out0_copy344_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid345_In0_c0 <= "" & bh7_w59_1_c0 & bh7_w59_5_c0 & bh7_w59_6_c0 & bh7_w59_7_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid345_In1_c0 <= "" & bh7_w60_1_c0;
   bh7_w59_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0(0);
   bh7_w60_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0(1);
   bh7_w61_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid345: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid345_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid345_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_copy346_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid345_Out0_copy346_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid347_In0_c0 <= "" & bh7_w60_2_c0 & bh7_w60_6_c0 & bh7_w60_7_c0 & bh7_w60_8_c0 & bh7_w60_9_c0 & bh7_w60_10_c0;
   bh7_w60_13_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0(0);
   bh7_w61_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0(1);
   bh7_w62_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid347: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid347_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_copy348_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid347_Out0_copy348_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid349_In0_c0 <= "" & bh7_w61_1_c0 & bh7_w61_2_c0 & bh7_w61_6_c0 & bh7_w61_7_c0 & bh7_w61_8_c0 & bh7_w61_9_c0;
   bh7_w61_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0(0);
   bh7_w62_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0(1);
   bh7_w63_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid349: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid349_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_copy350_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid349_Out0_copy350_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid351_In0_c0 <= "" & bh7_w62_1_c0 & bh7_w62_5_c0 & bh7_w62_6_c0 & bh7_w62_7_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid351_In1_c0 <= "" & bh7_w63_1_c0;
   bh7_w62_11_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0(0);
   bh7_w63_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0(1);
   bh7_w64_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid351: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid351_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid351_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_copy352_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid351_Out0_copy352_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid353_In0_c0 <= "" & bh7_w63_2_c0 & bh7_w63_6_c0 & bh7_w63_7_c0 & bh7_w63_8_c0 & bh7_w63_9_c0 & bh7_w63_10_c0;
   bh7_w63_13_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0(0);
   bh7_w64_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0(1);
   bh7_w65_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid353: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid353_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_copy354_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid353_Out0_copy354_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid355_In0_c0 <= "" & bh7_w64_1_c0 & bh7_w64_2_c0 & bh7_w64_6_c0 & bh7_w64_7_c0 & bh7_w64_8_c0 & bh7_w64_9_c0;
   bh7_w64_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0(0);
   bh7_w65_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0(1);
   bh7_w66_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid355: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid355_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_copy356_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid355_Out0_copy356_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid357_In0_c0 <= "" & bh7_w65_1_c0 & bh7_w65_4_c0 & bh7_w65_5_c0 & bh7_w65_6_c0 & bh7_w65_7_c0 & bh7_w65_8_c0;
   bh7_w65_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0(0);
   bh7_w66_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0(1);
   bh7_w67_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid357: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid357_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_copy358_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid357_Out0_copy358_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid359_In0_c0 <= "" & bh7_w66_1_c0 & bh7_w66_2_c0 & bh7_w66_5_c0 & bh7_w66_6_c0 & bh7_w66_7_c0 & bh7_w66_8_c0;
   bh7_w66_12_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0(0);
   bh7_w67_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0(1);
   bh7_w68_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid359: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid359_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_copy360_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid359_Out0_copy360_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid361_In0_c0 <= "" & bh7_w67_1_c0 & bh7_w67_2_c0 & bh7_w67_5_c0 & bh7_w67_6_c0 & bh7_w67_7_c0 & bh7_w67_8_c0;
   bh7_w67_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0(0);
   bh7_w68_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0(1);
   bh7_w69_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid361: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid361_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_copy362_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid361_Out0_copy362_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid363_In0_c0 <= "" & bh7_w68_1_c0 & bh7_w68_4_c0 & bh7_w68_5_c0 & bh7_w68_6_c0 & bh7_w68_7_c0 & bh7_w68_8_c0;
   bh7_w68_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0(0);
   bh7_w69_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0(1);
   bh7_w70_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid363: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid363_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_copy364_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid363_Out0_copy364_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid365_In0_c0 <= "" & bh7_w69_1_c0 & bh7_w69_2_c0 & bh7_w69_5_c0 & bh7_w69_6_c0 & bh7_w69_7_c0 & bh7_w69_8_c0;
   bh7_w69_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0(0);
   bh7_w70_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0(1);
   bh7_w71_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid365: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid365_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_copy366_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid365_Out0_copy366_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid367_In0_c0 <= "" & bh7_w70_1_c0 & bh7_w70_2_c0 & bh7_w70_5_c0 & bh7_w70_6_c0 & bh7_w70_7_c0 & bh7_w70_8_c0;
   bh7_w70_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0(0);
   bh7_w71_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0(1);
   bh7_w72_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid367: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid367_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_copy368_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid367_Out0_copy368_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid369_In0_c0 <= "" & bh7_w71_1_c0 & bh7_w71_4_c0 & bh7_w71_5_c0 & bh7_w71_6_c0 & bh7_w71_7_c0 & bh7_w71_8_c0;
   bh7_w71_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0(0);
   bh7_w72_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0(1);
   bh7_w73_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid369: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid369_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_copy370_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid369_Out0_copy370_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid371_In0_c0 <= "" & bh7_w72_1_c0 & bh7_w72_2_c0 & bh7_w72_5_c0 & bh7_w72_6_c0 & bh7_w72_7_c0 & bh7_w72_8_c0;
   bh7_w72_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0(0);
   bh7_w73_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0(1);
   bh7_w74_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid371: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid371_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_copy372_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid371_Out0_copy372_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid373_In0_c0 <= "" & bh7_w73_1_c0 & bh7_w73_2_c0 & bh7_w73_5_c0 & bh7_w73_6_c0 & bh7_w73_7_c0 & bh7_w73_8_c0;
   bh7_w73_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0(0);
   bh7_w74_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0(1);
   bh7_w75_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid373: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid373_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_copy374_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid373_Out0_copy374_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid375_In0_c0 <= "" & bh7_w74_1_c0 & bh7_w74_4_c0 & bh7_w74_5_c0 & bh7_w74_6_c0 & bh7_w74_7_c0 & bh7_w74_8_c0;
   bh7_w74_11_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0(0);
   bh7_w75_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0(1);
   bh7_w76_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid375: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid375_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_copy376_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid375_Out0_copy376_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid377_In0_c0 <= "" & bh7_w75_0_c0 & bh7_w75_3_c0 & bh7_w75_4_c0 & bh7_w75_5_c0 & bh7_w75_6_c0 & bh7_w75_7_c0;
   bh7_w75_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0(0);
   bh7_w76_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0(1);
   bh7_w77_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid377: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid377_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_copy378_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid377_Out0_copy378_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid379_In0_c0 <= "" & bh7_w76_0_c0 & bh7_w76_3_c0 & bh7_w76_4_c0 & bh7_w76_5_c0 & bh7_w76_6_c0 & bh7_w76_7_c0;
   bh7_w76_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0(0);
   bh7_w77_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0(1);
   bh7_w78_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid379: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid379_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_copy380_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid379_Out0_copy380_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid381_In0_c0 <= "" & bh7_w77_2_c0 & bh7_w77_3_c0 & bh7_w77_4_c0 & bh7_w77_5_c0 & bh7_w77_6_c0 & bh7_w77_7_c0;
   bh7_w77_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0(0);
   bh7_w78_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0(1);
   bh7_w79_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid381: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid381_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_copy382_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid381_Out0_copy382_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid383_In0_c0 <= "" & bh7_w78_2_c0 & bh7_w78_3_c0 & bh7_w78_4_c0 & bh7_w78_5_c0 & bh7_w78_6_c0 & bh7_w78_7_c0;
   bh7_w78_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0(0);
   bh7_w79_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0(1);
   bh7_w80_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid383: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid383_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_copy384_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid383_Out0_copy384_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid385_In0_c0 <= "" & bh7_w79_2_c0 & bh7_w79_3_c0 & bh7_w79_4_c0 & bh7_w79_5_c0 & bh7_w79_6_c0 & bh7_w79_7_c0;
   bh7_w79_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0(0);
   bh7_w80_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0(1);
   bh7_w81_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid385: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid385_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_copy386_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid385_Out0_copy386_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid387_In0_c0 <= "" & bh7_w80_2_c0 & bh7_w80_3_c0 & bh7_w80_4_c0 & bh7_w80_5_c0 & bh7_w80_6_c0 & bh7_w80_7_c0;
   bh7_w80_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0(0);
   bh7_w81_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0(1);
   bh7_w82_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid387: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid387_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_copy388_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid387_Out0_copy388_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid389_In0_c0 <= "" & bh7_w81_2_c0 & bh7_w81_3_c0 & bh7_w81_4_c0 & bh7_w81_5_c0 & bh7_w81_6_c0 & bh7_w81_7_c0;
   bh7_w81_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0(0);
   bh7_w82_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0(1);
   bh7_w83_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid389: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid389_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_copy390_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid389_Out0_copy390_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid391_In0_c0 <= "" & bh7_w82_1_c0 & bh7_w82_2_c0 & bh7_w82_3_c0 & bh7_w82_4_c0 & bh7_w82_5_c0 & bh7_w82_6_c0;
   bh7_w82_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0(0);
   bh7_w83_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0(1);
   bh7_w84_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid391: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid391_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_copy392_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid391_Out0_copy392_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid393_In0_c0 <= "" & bh7_w83_1_c0 & bh7_w83_2_c0 & bh7_w83_3_c0 & bh7_w83_4_c0 & bh7_w83_5_c0 & bh7_w83_6_c0;
   bh7_w83_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0(0);
   bh7_w84_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0(1);
   bh7_w85_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid393: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid393_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_copy394_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid393_Out0_copy394_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid395_In0_c0 <= "" & bh7_w84_1_c0 & bh7_w84_2_c0 & bh7_w84_3_c0 & bh7_w84_4_c0 & bh7_w84_5_c0 & bh7_w84_6_c0;
   bh7_w84_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0(0);
   bh7_w85_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0(1);
   bh7_w86_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid395: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid395_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_copy396_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid395_Out0_copy396_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid397_In0_c0 <= "" & bh7_w85_1_c0 & bh7_w85_2_c0 & bh7_w85_3_c0 & bh7_w85_4_c0 & bh7_w85_5_c0 & bh7_w85_6_c0;
   bh7_w85_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0(0);
   bh7_w86_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0(1);
   bh7_w87_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid397: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid397_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_copy398_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid397_Out0_copy398_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid401_In0_c0 <= "" & bh7_w86_1_c0 & bh7_w86_2_c0 & bh7_w86_3_c0 & bh7_w86_4_c0 & bh7_w86_5_c0;
   bh7_w86_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0(0);
   bh7_w87_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0(1);
   bh7_w88_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid401: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid401_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_copy402_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid401_Out0_copy402_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid403_In0_c0 <= "" & bh7_w87_1_c0 & bh7_w87_2_c0 & bh7_w87_3_c0 & bh7_w87_4_c0 & bh7_w87_5_c0 & bh7_w87_6_c0;
   bh7_w87_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0(0);
   bh7_w88_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0(1);
   bh7_w89_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid403: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid403_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_copy404_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid403_Out0_copy404_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid405_In0_c0 <= "" & bh7_w88_1_c0 & bh7_w88_2_c0 & bh7_w88_3_c0 & bh7_w88_4_c0 & bh7_w88_5_c0 & bh7_w88_6_c0;
   bh7_w88_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0(0);
   bh7_w89_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0(1);
   bh7_w90_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid405: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid405_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_copy406_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid405_Out0_copy406_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid407_In0_c0 <= "" & bh7_w89_1_c0 & bh7_w89_2_c0 & bh7_w89_3_c0 & bh7_w89_4_c0 & bh7_w89_5_c0;
   bh7_w89_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0(0);
   bh7_w90_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0(1);
   bh7_w91_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid407: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid407_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_copy408_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid407_Out0_copy408_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid409_In0_c0 <= "" & bh7_w90_1_c0 & bh7_w90_2_c0 & bh7_w90_3_c0 & bh7_w90_4_c0 & bh7_w90_5_c0 & bh7_w90_6_c0;
   bh7_w90_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0(0);
   bh7_w91_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0(1);
   bh7_w92_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid409: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid409_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_copy410_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid409_Out0_copy410_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid411_In0_c0 <= "" & bh7_w91_1_c0 & bh7_w91_2_c0 & bh7_w91_3_c0 & bh7_w91_4_c0 & bh7_w91_5_c0 & bh7_w91_6_c0;
   bh7_w91_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0(0);
   bh7_w92_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0(1);
   bh7_w93_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid411: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid411_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_copy412_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid411_Out0_copy412_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid413_In0_c0 <= "" & bh7_w92_1_c0 & bh7_w92_2_c0 & bh7_w92_3_c0 & bh7_w92_4_c0 & bh7_w92_5_c0;
   bh7_w92_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0(0);
   bh7_w93_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0(1);
   bh7_w94_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid413: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid413_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_copy414_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid413_Out0_copy414_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid415_In0_c0 <= "" & bh7_w93_1_c0 & bh7_w93_2_c0 & bh7_w93_3_c0 & bh7_w93_4_c0 & bh7_w93_5_c0 & bh7_w93_6_c0;
   bh7_w93_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0(0);
   bh7_w94_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0(1);
   bh7_w95_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid415: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid415_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_copy416_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid415_Out0_copy416_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid417_In0_c0 <= "" & bh7_w94_1_c0 & bh7_w94_2_c0 & bh7_w94_3_c0 & bh7_w94_4_c0 & bh7_w94_5_c0 & bh7_w94_6_c0;
   bh7_w94_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0(0);
   bh7_w95_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0(1);
   bh7_w96_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid417: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid417_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_copy418_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid417_Out0_copy418_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid419_In0_c0 <= "" & bh7_w95_1_c0 & bh7_w95_2_c0 & bh7_w95_3_c0 & bh7_w95_4_c0 & bh7_w95_5_c0;
   bh7_w95_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0(0);
   bh7_w96_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0(1);
   bh7_w97_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid419: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid419_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_copy420_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid419_Out0_copy420_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid421_In0_c0 <= "" & bh7_w96_1_c0 & bh7_w96_2_c0 & bh7_w96_3_c0 & bh7_w96_4_c0 & bh7_w96_5_c0 & bh7_w96_6_c0;
   bh7_w96_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0(0);
   bh7_w97_9_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0(1);
   bh7_w98_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid421: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid421_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_copy422_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid421_Out0_copy422_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid423_In0_c0 <= "" & bh7_w97_1_c0 & bh7_w97_2_c0 & bh7_w97_3_c0 & bh7_w97_4_c0 & bh7_w97_5_c0 & bh7_w97_6_c0;
   bh7_w97_10_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0(0);
   bh7_w98_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0(1);
   bh7_w99_6_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid423: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid423_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_copy424_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid423_Out0_copy424_c0; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid425_In0_c0 <= "" & bh7_w98_1_c0 & bh7_w98_2_c0 & bh7_w98_3_c0 & bh7_w98_4_c0 & bh7_w98_5_c0;
   bh7_w98_8_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0(0);
   bh7_w99_7_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0(1);
   bh7_w100_6_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0(2);
   Compressor_5_3_Freq300_uid400_uid425: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid425_In0_c0,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_copy426_c0);
   Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_c0 <= Compressor_5_3_Freq300_uid400_bh7_uid425_Out0_copy426_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid427_In0_c0 <= "" & bh7_w99_0_c0 & bh7_w99_1_c0 & bh7_w99_2_c0 & bh7_w99_3_c0 & bh7_w99_4_c0 & bh7_w99_5_c0;
   bh7_w99_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0(0);
   bh7_w100_7_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0(1);
   bh7_w101_3_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid427: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid427_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_copy428_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid427_Out0_copy428_c0; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid429_In0_c0 <= "" & bh7_w100_0_c0 & bh7_w100_1_c0 & bh7_w100_2_c0 & bh7_w100_3_c0 & bh7_w100_4_c0 & bh7_w100_5_c0;
   bh7_w100_8_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0(0);
   bh7_w101_4_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0(1);
   bh7_w102_4_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0(2);
   Compressor_6_3_Freq300_uid334_uid429: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid429_In0_c0,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_copy430_c0);
   Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_c0 <= Compressor_6_3_Freq300_uid334_bh7_uid429_Out0_copy430_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid433_In0_c0 <= "" & bh7_w101_0_c0 & bh7_w101_1_c0 & bh7_w101_2_c0;
   bh7_w101_5_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_c0(0);
   bh7_w102_5_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid433: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid433_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_copy434_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid433_Out0_copy434_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid435_In0_c0 <= "" & bh7_w102_0_c0 & bh7_w102_1_c0 & bh7_w102_2_c0 & bh7_w102_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid435_In1_c0 <= "" & bh7_w103_0_c0;
   bh7_w102_6_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0(0);
   bh7_w103_2_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0(1);
   bh7_w104_1_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid435: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid435_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid435_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_copy436_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid435_Out0_copy436_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid437_In0_c0 <= "" & bh7_w51_9_c0 & bh7_w51_8_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid437_In1_c0 <= "" & bh7_w52_10_c0 & bh7_w52_9_c0;
   bh7_w51_10_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0(0);
   bh7_w52_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0(1);
   bh7_w53_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid437: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid437_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid437_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_copy438_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid437_Out0_copy438_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid439_In0_c0 <= "" & bh7_w53_11_c0 & bh7_w53_10_c0 & bh7_w53_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid439_In1_c0 <= "" & bh7_w54_12_c0 & bh7_w54_11_c0;
   bh7_w53_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0(0);
   bh7_w54_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0(1);
   bh7_w55_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid439: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid439_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid439_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_copy440_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid439_Out0_copy440_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid441_In0_c0 <= "" & bh7_w55_10_c0 & bh7_w55_12_c0 & bh7_w55_11_c0;
   bh7_w55_14_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_c0(0);
   bh7_w56_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid441: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid441_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_copy442_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid441_Out0_copy442_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid443_In0_c0 <= "" & bh7_w56_8_c0 & bh7_w56_11_c0 & bh7_w56_10_c0 & bh7_w56_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid443_In1_c0 <= "" & "0";
   bh7_w56_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0(0);
   bh7_w57_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0(1);
   bh7_w58_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid443: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid443_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid443_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_copy444_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid443_Out0_copy444_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid445_In0_c0 <= "" & bh7_w57_12_c0 & bh7_w57_13_c0 & bh7_w57_11_c0;
   bh7_w57_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_c0(0);
   bh7_w58_14_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid445: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid445_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_copy446_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid445_Out0_copy446_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid447_In0_c0 <= "" & bh7_w58_10_c0 & bh7_w58_12_c0 & bh7_w58_11_c0;
   bh7_w58_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_c0(0);
   bh7_w59_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid447: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid447_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_copy448_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid447_Out0_copy448_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid449_In0_c0 <= "" & bh7_w59_8_c0 & bh7_w59_11_c0 & bh7_w59_10_c0 & bh7_w59_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid449_In1_c0 <= "" & "0";
   bh7_w59_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0(0);
   bh7_w60_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0(1);
   bh7_w61_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid449: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid449_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid449_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_copy450_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid449_Out0_copy450_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid451_In0_c0 <= "" & bh7_w60_12_c0 & bh7_w60_13_c0 & bh7_w60_11_c0;
   bh7_w60_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_c0(0);
   bh7_w61_14_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid451: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid451_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_copy452_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid451_Out0_copy452_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid453_In0_c0 <= "" & bh7_w61_10_c0 & bh7_w61_12_c0 & bh7_w61_11_c0;
   bh7_w61_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_c0(0);
   bh7_w62_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid453: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid453_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_copy454_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid453_Out0_copy454_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid455_In0_c0 <= "" & bh7_w62_8_c0 & bh7_w62_11_c0 & bh7_w62_10_c0 & bh7_w62_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid455_In1_c0 <= "" & "0";
   bh7_w62_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0(0);
   bh7_w63_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0(1);
   bh7_w64_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid455: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid455_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid455_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_copy456_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid455_Out0_copy456_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid457_In0_c0 <= "" & bh7_w63_12_c0 & bh7_w63_13_c0 & bh7_w63_11_c0;
   bh7_w63_15_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_c0(0);
   bh7_w64_14_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid457: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid457_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_copy458_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid457_Out0_copy458_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid459_In0_c0 <= "" & bh7_w64_10_c0 & bh7_w64_12_c0 & bh7_w64_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid459_In1_c0 <= "" & bh7_w65_11_c0 & bh7_w65_10_c0;
   bh7_w64_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0(0);
   bh7_w65_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0(1);
   bh7_w66_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid459: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid459_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid459_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_copy460_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid459_Out0_copy460_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid461_In0_c0 <= "" & bh7_w66_9_c0 & bh7_w66_12_c0 & bh7_w66_11_c0 & bh7_w66_10_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid461_In1_c0 <= "" & "0";
   bh7_w66_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0(0);
   bh7_w67_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0(1);
   bh7_w68_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid461: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid461_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid461_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_copy462_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid461_Out0_copy462_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid463_In0_c0 <= "" & bh7_w67_11_c0 & bh7_w67_10_c0 & bh7_w67_9_c0;
   bh7_w67_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_c0(0);
   bh7_w68_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid463: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid463_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_copy464_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid463_Out0_copy464_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid465_In0_c0 <= "" & bh7_w68_11_c0 & bh7_w68_10_c0 & bh7_w68_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid465_In1_c0 <= "" & bh7_w69_11_c0 & bh7_w69_10_c0;
   bh7_w68_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0(0);
   bh7_w69_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0(1);
   bh7_w70_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid465: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid465_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid465_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_copy466_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid465_Out0_copy466_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid467_In0_c0 <= "" & bh7_w70_11_c0 & bh7_w70_10_c0 & bh7_w70_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid467_In1_c0 <= "" & bh7_w71_11_c0 & bh7_w71_10_c0;
   bh7_w70_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0(0);
   bh7_w71_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0(1);
   bh7_w72_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid467: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid467_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid467_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_copy468_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid467_Out0_copy468_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid469_In0_c0 <= "" & bh7_w72_11_c0 & bh7_w72_10_c0 & bh7_w72_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid469_In1_c0 <= "" & bh7_w73_11_c0 & bh7_w73_10_c0;
   bh7_w72_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0(0);
   bh7_w73_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0(1);
   bh7_w74_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid469: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid469_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid469_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_copy470_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid469_Out0_copy470_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid471_In0_c0 <= "" & bh7_w74_11_c0 & bh7_w74_10_c0 & bh7_w74_9_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid471_In1_c0 <= "" & bh7_w75_10_c0 & bh7_w75_9_c0;
   bh7_w74_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0(0);
   bh7_w75_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0(1);
   bh7_w76_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid471: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid471_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid471_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_copy472_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid471_Out0_copy472_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid473_In0_c0 <= "" & bh7_w76_10_c0 & bh7_w76_9_c0 & bh7_w76_8_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid473_In1_c0 <= "" & bh7_w77_10_c0 & bh7_w77_9_c0;
   bh7_w76_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0(0);
   bh7_w77_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0(1);
   bh7_w78_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid473: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid473_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid473_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_copy474_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid473_Out0_copy474_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid475_In0_c0 <= "" & bh7_w78_10_c0 & bh7_w78_9_c0 & bh7_w78_8_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid475_In1_c0 <= "" & bh7_w79_10_c0 & bh7_w79_9_c0;
   bh7_w78_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0(0);
   bh7_w79_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0(1);
   bh7_w80_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid475: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid475_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid475_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_copy476_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid475_Out0_copy476_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid477_In0_c0 <= "" & bh7_w80_10_c0 & bh7_w80_9_c0 & bh7_w80_8_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid477_In1_c0 <= "" & bh7_w81_10_c0 & bh7_w81_9_c0;
   bh7_w80_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0(0);
   bh7_w81_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0(1);
   bh7_w82_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid477: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid477_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid477_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_copy478_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid477_Out0_copy478_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid479_In0_c0 <= "" & bh7_w82_7_c0 & bh7_w82_10_c0 & bh7_w82_9_c0 & bh7_w82_8_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid479_In1_c0 <= "" & "0";
   bh7_w82_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0(0);
   bh7_w83_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0(1);
   bh7_w84_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid479: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid479_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid479_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_copy480_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid479_Out0_copy480_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid481_In0_c0 <= "" & bh7_w83_9_c0 & bh7_w83_8_c0 & bh7_w83_7_c0;
   bh7_w83_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_c0(0);
   bh7_w84_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid481: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid481_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_copy482_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid481_Out0_copy482_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid483_In0_c0 <= "" & bh7_w84_9_c0 & bh7_w84_8_c0 & bh7_w84_7_c0;
   bh7_w84_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_c0(0);
   bh7_w85_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid483: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid483_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_copy484_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid483_Out0_copy484_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid485_In0_c0 <= "" & bh7_w85_7_c0 & bh7_w85_10_c0 & bh7_w85_9_c0 & bh7_w85_8_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid485_In1_c0 <= "" & "0";
   bh7_w85_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0(0);
   bh7_w86_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0(1);
   bh7_w87_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid485: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid485_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid485_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_copy486_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid485_Out0_copy486_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid487_In0_c0 <= "" & bh7_w86_8_c0 & bh7_w86_7_c0 & bh7_w86_6_c0;
   bh7_w86_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_c0(0);
   bh7_w87_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid487: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid487_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_copy488_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid487_Out0_copy488_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid489_In0_c0 <= "" & bh7_w87_8_c0 & bh7_w87_9_c0 & bh7_w87_7_c0;
   bh7_w87_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_c0(0);
   bh7_w88_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid489: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid489_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_copy490_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid489_Out0_copy490_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid491_In0_c0 <= "" & bh7_w88_7_c0 & bh7_w88_8_c0 & bh7_w88_10_c0 & bh7_w88_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid491_In1_c0 <= "" & "0";
   bh7_w88_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0(0);
   bh7_w89_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0(1);
   bh7_w90_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid491: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid491_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid491_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_copy492_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid491_Out0_copy492_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid493_In0_c0 <= "" & bh7_w89_8_c0 & bh7_w89_7_c0 & bh7_w89_6_c0;
   bh7_w89_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_c0(0);
   bh7_w90_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid493: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid493_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_copy494_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid493_Out0_copy494_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid495_In0_c0 <= "" & bh7_w90_8_c0 & bh7_w90_9_c0 & bh7_w90_7_c0;
   bh7_w90_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_c0(0);
   bh7_w91_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid495: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid495_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_copy496_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid495_Out0_copy496_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid497_In0_c0 <= "" & bh7_w91_7_c0 & bh7_w91_8_c0 & bh7_w91_10_c0 & bh7_w91_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid497_In1_c0 <= "" & "0";
   bh7_w91_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0(0);
   bh7_w92_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0(1);
   bh7_w93_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid497: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid497_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid497_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_copy498_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid497_Out0_copy498_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid499_In0_c0 <= "" & bh7_w92_8_c0 & bh7_w92_7_c0 & bh7_w92_6_c0;
   bh7_w92_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_c0(0);
   bh7_w93_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid499: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid499_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_copy500_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid499_Out0_copy500_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid501_In0_c0 <= "" & bh7_w93_8_c0 & bh7_w93_9_c0 & bh7_w93_7_c0;
   bh7_w93_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_c0(0);
   bh7_w94_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid501: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid501_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_copy502_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid501_Out0_copy502_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid503_In0_c0 <= "" & bh7_w94_7_c0 & bh7_w94_8_c0 & bh7_w94_10_c0 & bh7_w94_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid503_In1_c0 <= "" & "0";
   bh7_w94_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0(0);
   bh7_w95_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0(1);
   bh7_w96_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid503: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid503_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid503_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_copy504_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid503_Out0_copy504_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid505_In0_c0 <= "" & bh7_w95_8_c0 & bh7_w95_7_c0 & bh7_w95_6_c0;
   bh7_w95_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_c0(0);
   bh7_w96_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid505: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid505_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_copy506_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid505_Out0_copy506_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid507_In0_c0 <= "" & bh7_w96_8_c0 & bh7_w96_9_c0 & bh7_w96_7_c0;
   bh7_w96_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_c0(0);
   bh7_w97_11_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid507: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid507_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_copy508_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid507_Out0_copy508_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid509_In0_c0 <= "" & bh7_w97_7_c0 & bh7_w97_8_c0 & bh7_w97_10_c0 & bh7_w97_9_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid509_In1_c0 <= "" & "0";
   bh7_w97_12_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0(0);
   bh7_w98_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0(1);
   bh7_w99_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid509: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid509_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid509_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_copy510_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid509_Out0_copy510_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid511_In0_c0 <= "" & bh7_w98_8_c0 & bh7_w98_7_c0 & bh7_w98_6_c0;
   bh7_w98_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_c0(0);
   bh7_w99_10_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid511: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid511_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_copy512_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid511_Out0_copy512_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid513_In0_c0 <= "" & bh7_w99_7_c0 & bh7_w99_8_c0 & bh7_w99_6_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid513_In1_c0 <= "" & bh7_w100_6_c0 & bh7_w100_8_c0;
   bh7_w99_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0(0);
   bh7_w100_9_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0(1);
   bh7_w101_6_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid513: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid513_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid513_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_copy514_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid513_Out0_copy514_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid515_In0_c0 <= "" & bh7_w101_5_c0 & bh7_w101_4_c0 & bh7_w101_3_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid515_In1_c0 <= "" & bh7_w102_6_c0 & bh7_w102_5_c0;
   bh7_w101_7_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0(0);
   bh7_w102_7_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0(1);
   bh7_w103_3_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid515: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid515_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid515_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_copy516_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid515_Out0_copy516_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid517_In0_c0 <= "" & bh7_w103_1_c0 & bh7_w103_2_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid517_In1_c0 <= "" & bh7_w104_0_c0 & bh7_w104_1_c0;
   bh7_w103_4_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0(0);
   bh7_w104_2_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0(1);
   bh7_w105_1_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid517: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid517_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid517_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_copy518_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid517_Out0_copy518_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid519_In0_c0 <= "" & bh7_w53_13_c0 & bh7_w53_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid519_In1_c0 <= "" & bh7_w54_13_c0 & bh7_w54_14_c0;
   bh7_w53_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0(0);
   bh7_w54_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0(1);
   bh7_w55_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid519: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid519_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid519_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_copy520_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid519_Out0_copy520_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid521_In0_c0 <= "" & bh7_w55_13_c0 & bh7_w55_14_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid521_In1_c0 <= "" & bh7_w56_13_c0 & bh7_w56_12_c0;
   bh7_w55_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0(0);
   bh7_w56_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0(1);
   bh7_w57_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid521: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid521_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid521_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_copy522_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid521_Out0_copy522_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid523_In0_c0 <= "" & bh7_w57_14_c0 & bh7_w57_15_c0 & "0";
   bh7_w57_17_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_c0(0);
   bh7_w58_16_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid523: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid523_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_copy524_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid523_Out0_copy524_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid525_In0_c0 <= "" & bh7_w58_13_c0 & bh7_w58_15_c0 & bh7_w58_14_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid525_In1_c0 <= "" & bh7_w59_13_c0 & bh7_w59_12_c0;
   bh7_w58_17_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0(0);
   bh7_w59_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0(1);
   bh7_w60_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid525: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid525_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid525_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_copy526_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid525_Out0_copy526_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid527_In0_c0 <= "" & bh7_w60_14_c0 & bh7_w60_15_c0 & "0";
   bh7_w60_17_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_c0(0);
   bh7_w61_16_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid527: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid527_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_copy528_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid527_Out0_copy528_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid529_In0_c0 <= "" & bh7_w61_13_c0 & bh7_w61_15_c0 & bh7_w61_14_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid529_In1_c0 <= "" & bh7_w62_13_c0 & bh7_w62_12_c0;
   bh7_w61_17_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0(0);
   bh7_w62_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0(1);
   bh7_w63_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid529: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid529_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid529_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_copy530_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid529_Out0_copy530_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid531_In0_c0 <= "" & bh7_w63_14_c0 & bh7_w63_15_c0 & "0";
   bh7_w63_17_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_c0(0);
   bh7_w64_16_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid531: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid531_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_copy532_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid531_Out0_copy532_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid533_In0_c0 <= "" & bh7_w64_13_c0 & bh7_w64_15_c0 & bh7_w64_14_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid533_In1_c0 <= "" & bh7_w65_9_c0 & bh7_w65_12_c0;
   bh7_w64_17_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0(0);
   bh7_w65_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0(1);
   bh7_w66_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid533: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid533_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid533_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_copy534_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid533_Out0_copy534_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid535_In0_c0 <= "" & bh7_w66_14_c0 & bh7_w66_13_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid535_In1_c0 <= "" & bh7_w67_12_c0 & bh7_w67_13_c0;
   bh7_w66_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0(0);
   bh7_w67_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0(1);
   bh7_w68_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid535: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid535_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid535_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_copy536_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid535_Out0_copy536_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid537_In0_c0 <= "" & bh7_w68_12_c0 & bh7_w68_14_c0 & bh7_w68_13_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid537_In1_c0 <= "" & bh7_w69_9_c0 & bh7_w69_12_c0;
   bh7_w68_16_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0(0);
   bh7_w69_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0(1);
   bh7_w70_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid537: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid537_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid537_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_copy538_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid537_Out0_copy538_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid539_In0_c0 <= "" & bh7_w70_13_c0 & bh7_w70_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid539_In1_c0 <= "" & bh7_w71_9_c0 & bh7_w71_12_c0;
   bh7_w70_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0(0);
   bh7_w71_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0(1);
   bh7_w72_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid539: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid539_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid539_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_copy540_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid539_Out0_copy540_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid541_In0_c0 <= "" & bh7_w72_13_c0 & bh7_w72_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid541_In1_c0 <= "" & bh7_w73_9_c0 & bh7_w73_12_c0;
   bh7_w72_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0(0);
   bh7_w73_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0(1);
   bh7_w74_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid541: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid541_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid541_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_copy542_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid541_Out0_copy542_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid543_In0_c0 <= "" & bh7_w74_13_c0 & bh7_w74_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid543_In1_c0 <= "" & bh7_w75_8_c0 & bh7_w75_11_c0;
   bh7_w74_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0(0);
   bh7_w75_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0(1);
   bh7_w76_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid543: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid543_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid543_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_copy544_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid543_Out0_copy544_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid545_In0_c0 <= "" & bh7_w76_12_c0 & bh7_w76_11_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid545_In1_c0 <= "" & bh7_w77_8_c0 & bh7_w77_11_c0;
   bh7_w76_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0(0);
   bh7_w77_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0(1);
   bh7_w78_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid545: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid545_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid545_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_copy546_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid545_Out0_copy546_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid547_In0_c0 <= "" & bh7_w78_12_c0 & bh7_w78_11_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid547_In1_c0 <= "" & bh7_w79_8_c0 & bh7_w79_11_c0;
   bh7_w78_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0(0);
   bh7_w79_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0(1);
   bh7_w80_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid547: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid547_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid547_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_copy548_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid547_Out0_copy548_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid549_In0_c0 <= "" & bh7_w80_12_c0 & bh7_w80_11_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid549_In1_c0 <= "" & bh7_w81_8_c0 & bh7_w81_11_c0;
   bh7_w80_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0(0);
   bh7_w81_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0(1);
   bh7_w82_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid549: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid549_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid549_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_copy550_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid549_Out0_copy550_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid551_In0_c0 <= "" & bh7_w82_12_c0 & bh7_w82_11_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid551_In1_c0 <= "" & bh7_w83_10_c0 & bh7_w83_11_c0;
   bh7_w82_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0(0);
   bh7_w83_12_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0(1);
   bh7_w84_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid551: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid551_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid551_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_copy552_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid551_Out0_copy552_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid553_In0_c0 <= "" & bh7_w84_10_c0 & bh7_w84_12_c0 & bh7_w84_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid553_In1_c0 <= "" & bh7_w85_12_c0 & bh7_w85_11_c0;
   bh7_w84_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0(0);
   bh7_w85_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0(1);
   bh7_w86_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid553: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid553_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid553_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_copy554_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid553_Out0_copy554_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid555_In0_c0 <= "" & bh7_w86_9_c0 & bh7_w86_10_c0 & "0";
   bh7_w86_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_c0(0);
   bh7_w87_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid555: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid555_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_copy556_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid555_Out0_copy556_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid557_In0_c0 <= "" & bh7_w87_10_c0 & bh7_w87_12_c0 & bh7_w87_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid557_In1_c0 <= "" & bh7_w88_12_c0 & bh7_w88_11_c0;
   bh7_w87_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0(0);
   bh7_w88_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0(1);
   bh7_w89_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid557: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid557_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid557_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_copy558_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid557_Out0_copy558_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid559_In0_c0 <= "" & bh7_w89_9_c0 & bh7_w89_10_c0 & "0";
   bh7_w89_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_c0(0);
   bh7_w90_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid559: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid559_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_copy560_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid559_Out0_copy560_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid561_In0_c0 <= "" & bh7_w90_10_c0 & bh7_w90_12_c0 & bh7_w90_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid561_In1_c0 <= "" & bh7_w91_12_c0 & bh7_w91_11_c0;
   bh7_w90_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0(0);
   bh7_w91_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0(1);
   bh7_w92_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid561: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid561_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid561_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_copy562_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid561_Out0_copy562_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid563_In0_c0 <= "" & bh7_w92_9_c0 & bh7_w92_10_c0 & "0";
   bh7_w92_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_c0(0);
   bh7_w93_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid563: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid563_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_copy564_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid563_Out0_copy564_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid565_In0_c0 <= "" & bh7_w93_10_c0 & bh7_w93_12_c0 & bh7_w93_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid565_In1_c0 <= "" & bh7_w94_12_c0 & bh7_w94_11_c0;
   bh7_w93_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0(0);
   bh7_w94_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0(1);
   bh7_w95_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid565: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid565_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid565_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_copy566_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid565_Out0_copy566_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid567_In0_c0 <= "" & bh7_w95_9_c0 & bh7_w95_10_c0 & "0";
   bh7_w95_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_c0(0);
   bh7_w96_13_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid567: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid567_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_copy568_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid567_Out0_copy568_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid569_In0_c0 <= "" & bh7_w96_10_c0 & bh7_w96_12_c0 & bh7_w96_11_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid569_In1_c0 <= "" & bh7_w97_12_c0 & bh7_w97_11_c0;
   bh7_w96_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0(0);
   bh7_w97_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0(1);
   bh7_w98_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid569: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid569_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid569_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_copy570_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid569_Out0_copy570_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid571_In0_c0 <= "" & bh7_w98_9_c0 & bh7_w98_10_c0 & "0";
   bh7_w98_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_c0(0);
   bh7_w99_12_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_c0(1);
   Compressor_3_2_Freq300_uid432_uid571: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid571_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_copy572_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid571_Out0_copy572_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid573_In0_c0 <= "" & bh7_w99_9_c0 & bh7_w99_11_c0 & bh7_w99_10_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid573_In1_c0 <= "" & bh7_w100_7_c0 & bh7_w100_9_c0;
   bh7_w99_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0(0);
   bh7_w100_10_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0(1);
   bh7_w101_8_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid573: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid573_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid573_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_copy574_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid573_Out0_copy574_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid575_In0_c0 <= "" & bh7_w101_7_c0 & bh7_w101_6_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid575_In1_c0 <= "" & bh7_w102_4_c0 & bh7_w102_7_c0;
   bh7_w101_9_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0(0);
   bh7_w102_8_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0(1);
   bh7_w103_5_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid575: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid575_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid575_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_copy576_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid575_Out0_copy576_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid577_In0_c0 <= "" & bh7_w103_4_c0 & bh7_w103_3_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid577_In1_c0 <= "" & bh7_w104_2_c0;
   bh7_w103_6_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0(0);
   bh7_w104_3_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0(1);
   bh7_w105_2_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid577: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid577_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid577_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_copy578_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid577_Out0_copy578_c0; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid579_In0_c0 <= "" & bh7_w105_0_c0 & bh7_w105_1_c0 & "0";
   bh7_w105_3_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_c0(0);
   Compressor_3_2_Freq300_uid432_uid579: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid579_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_copy580_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_c0 <= Compressor_3_2_Freq300_uid432_bh7_uid579_Out0_copy580_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid581_In0_c0 <= "" & bh7_w55_16_c0 & bh7_w55_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid581_In1_c0 <= "" & bh7_w56_14_c0;
   bh7_w55_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0(0);
   bh7_w56_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0(1);
   bh7_w57_18_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid581: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid581_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid581_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_copy582_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid581_Out0_copy582_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid583_In0_c0 <= "" & bh7_w57_16_c0 & bh7_w57_17_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid583_In1_c0 <= "" & bh7_w58_16_c0 & bh7_w58_17_c0;
   bh7_w57_19_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0(0);
   bh7_w58_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0(1);
   bh7_w59_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid583: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid583_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid583_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_copy584_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid583_Out0_copy584_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid585_In0_c0 <= "" & bh7_w60_16_c0 & bh7_w60_17_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid585_In1_c0 <= "" & bh7_w61_16_c0 & bh7_w61_17_c0;
   bh7_w60_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0(0);
   bh7_w61_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0(1);
   bh7_w62_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid585: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid585_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid585_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_copy586_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid585_Out0_copy586_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid587_In0_c0 <= "" & bh7_w63_16_c0 & bh7_w63_17_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid587_In1_c0 <= "" & bh7_w64_16_c0 & bh7_w64_17_c0;
   bh7_w63_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0(0);
   bh7_w64_18_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0(1);
   bh7_w65_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid587: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid587_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid587_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_copy588_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid587_Out0_copy588_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid589_In0_c0 <= "" & bh7_w66_15_c0 & bh7_w66_16_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid589_In1_c0 <= "" & bh7_w67_14_c0;
   bh7_w66_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0(0);
   bh7_w67_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0(1);
   bh7_w68_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid589: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid589_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid589_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_copy590_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid589_Out0_copy590_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid591_In0_c0 <= "" & bh7_w68_15_c0 & bh7_w68_16_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid591_In1_c0 <= "" & bh7_w69_13_c0;
   bh7_w68_18_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0(0);
   bh7_w69_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0(1);
   bh7_w70_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid591: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid591_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid591_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_copy592_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid591_Out0_copy592_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid593_In0_c0 <= "" & bh7_w70_14_c0 & bh7_w70_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid593_In1_c0 <= "" & bh7_w71_13_c0;
   bh7_w70_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0(0);
   bh7_w71_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0(1);
   bh7_w72_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid593: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid593_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid593_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_copy594_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid593_Out0_copy594_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid595_In0_c0 <= "" & bh7_w72_15_c0 & bh7_w72_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid595_In1_c0 <= "" & bh7_w73_13_c0;
   bh7_w72_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0(0);
   bh7_w73_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0(1);
   bh7_w74_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid595: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid595_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid595_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_copy596_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid595_Out0_copy596_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid597_In0_c0 <= "" & bh7_w74_15_c0 & bh7_w74_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid597_In1_c0 <= "" & bh7_w75_12_c0;
   bh7_w74_17_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0(0);
   bh7_w75_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0(1);
   bh7_w76_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid597: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid597_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid597_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_copy598_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid597_Out0_copy598_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid599_In0_c0 <= "" & bh7_w76_14_c0 & bh7_w76_13_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid599_In1_c0 <= "" & bh7_w77_12_c0;
   bh7_w76_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0(0);
   bh7_w77_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0(1);
   bh7_w78_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid599: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid599_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid599_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_copy600_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid599_Out0_copy600_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid601_In0_c0 <= "" & bh7_w78_14_c0 & bh7_w78_13_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid601_In1_c0 <= "" & bh7_w79_12_c0;
   bh7_w78_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0(0);
   bh7_w79_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0(1);
   bh7_w80_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid601: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid601_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid601_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_copy602_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid601_Out0_copy602_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid603_In0_c0 <= "" & bh7_w80_14_c0 & bh7_w80_13_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid603_In1_c0 <= "" & bh7_w81_12_c0;
   bh7_w80_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0(0);
   bh7_w81_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0(1);
   bh7_w82_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid603: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid603_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid603_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_copy604_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid603_Out0_copy604_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid605_In0_c0 <= "" & bh7_w82_14_c0 & bh7_w82_13_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid605_In1_c0 <= "" & bh7_w83_12_c0;
   bh7_w82_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0(0);
   bh7_w83_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0(1);
   bh7_w84_15_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid605: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid605_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid605_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_copy606_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid605_Out0_copy606_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid607_In0_c0 <= "" & bh7_w84_13_c0 & bh7_w84_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid607_In1_c0 <= "" & bh7_w85_13_c0;
   bh7_w84_16_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0(0);
   bh7_w85_14_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0(1);
   bh7_w86_13_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid607: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid607_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid607_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_copy608_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid607_Out0_copy608_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid609_In0_c0 <= "" & bh7_w86_11_c0 & bh7_w86_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid609_In1_c0 <= "" & bh7_w87_13_c0 & bh7_w87_14_c0;
   bh7_w86_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0(0);
   bh7_w87_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0(1);
   bh7_w88_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid609: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid609_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid609_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_copy610_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid609_Out0_copy610_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid611_In0_c0 <= "" & bh7_w89_11_c0 & bh7_w89_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid611_In1_c0 <= "" & bh7_w90_13_c0 & bh7_w90_14_c0;
   bh7_w89_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0(0);
   bh7_w90_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0(1);
   bh7_w91_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid611: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid611_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid611_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_copy612_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid611_Out0_copy612_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid613_In0_c0 <= "" & bh7_w92_11_c0 & bh7_w92_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid613_In1_c0 <= "" & bh7_w93_13_c0 & bh7_w93_14_c0;
   bh7_w92_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0(0);
   bh7_w93_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0(1);
   bh7_w94_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid613: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid613_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid613_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_copy614_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid613_Out0_copy614_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid615_In0_c0 <= "" & bh7_w95_11_c0 & bh7_w95_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid615_In1_c0 <= "" & bh7_w96_13_c0 & bh7_w96_14_c0;
   bh7_w95_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0(0);
   bh7_w96_15_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0(1);
   bh7_w97_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid615: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid615_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid615_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_copy616_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid615_Out0_copy616_c0; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid617_In0_c0 <= "" & bh7_w98_11_c0 & bh7_w98_12_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid617_In1_c0 <= "" & bh7_w99_12_c0 & bh7_w99_13_c0;
   bh7_w98_13_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0(0);
   bh7_w99_14_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0(1);
   bh7_w100_11_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0(2);
   Compressor_23_3_Freq300_uid322_uid617: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid617_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid617_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_copy618_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_c0 <= Compressor_23_3_Freq300_uid322_bh7_uid617_Out0_copy618_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid619_In0_c0 <= "" & bh7_w101_8_c0 & bh7_w101_9_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid619_In1_c0 <= "" & bh7_w102_8_c0;
   bh7_w101_10_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0(0);
   bh7_w102_9_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0(1);
   bh7_w103_7_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid619: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid619_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid619_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_copy620_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid619_Out0_copy620_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid621_In0_c0 <= "" & bh7_w103_6_c0 & bh7_w103_5_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid621_In1_c0 <= "" & bh7_w104_3_c0;
   bh7_w103_8_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0(0);
   bh7_w104_4_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0(1);
   bh7_w105_4_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0(2);
   Compressor_14_3_Freq300_uid326_uid621: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid621_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid621_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_copy622_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid621_Out0_copy622_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid623_In0_c0 <= "" & bh7_w105_3_c0 & bh7_w105_2_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid623_In1_c0 <= "" & "0";
   bh7_w105_5_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_c0(0);
   Compressor_14_3_Freq300_uid326_uid623: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid623_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid623_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_copy624_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_c0 <= Compressor_14_3_Freq300_uid326_bh7_uid623_Out0_copy624_c0; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid625_In0_c0 <= "" & bh7_w57_18_c0 & bh7_w57_19_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid625_In1_c0 <= "" & bh7_w58_18_c0;
   bh7_w57_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1(0);
   bh7_w58_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1(1);
   bh7_w59_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid625: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid625_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid625_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid625_Out0_copy626_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid627_In0_c0 <= "" & bh7_w59_14_c0 & bh7_w59_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid627_In1_c0 <= "" & bh7_w60_18_c0;
   bh7_w59_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1(0);
   bh7_w60_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1(1);
   bh7_w61_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid627: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid627_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid627_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid627_Out0_copy628_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid629_In0_c0 <= "" & bh7_w62_14_c0 & bh7_w62_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid629_In1_c0 <= "" & bh7_w63_18_c0;
   bh7_w62_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1(0);
   bh7_w63_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1(1);
   bh7_w64_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid629: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid629_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid629_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid629_Out0_copy630_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid631_In0_c0 <= "" & bh7_w65_13_c0 & bh7_w65_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid631_In1_c0 <= "" & bh7_w66_17_c0;
   bh7_w65_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1(0);
   bh7_w66_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1(1);
   bh7_w67_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid631: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid631_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid631_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid631_Out0_copy632_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid633_In0_c0 <= "" & bh7_w68_17_c0 & bh7_w68_18_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid633_In1_c0 <= "" & bh7_w69_14_c0;
   bh7_w68_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1(0);
   bh7_w69_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1(1);
   bh7_w70_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid633: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid633_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid633_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid633_Out0_copy634_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid635_In0_c0 <= "" & bh7_w70_16_c0 & bh7_w70_17_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid635_In1_c0 <= "" & bh7_w71_14_c0;
   bh7_w70_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1(0);
   bh7_w71_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1(1);
   bh7_w72_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid635: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid635_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid635_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid635_Out0_copy636_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid637_In0_c0 <= "" & bh7_w72_16_c0 & bh7_w72_17_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid637_In1_c0 <= "" & bh7_w73_14_c0;
   bh7_w72_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1(0);
   bh7_w73_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1(1);
   bh7_w74_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid637: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid637_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid637_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid637_Out0_copy638_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid639_In0_c0 <= "" & bh7_w74_17_c0 & bh7_w74_16_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid639_In1_c0 <= "" & bh7_w75_13_c0;
   bh7_w74_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1(0);
   bh7_w75_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1(1);
   bh7_w76_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid639: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid639_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid639_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid639_Out0_copy640_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid641_In0_c0 <= "" & bh7_w76_16_c0 & bh7_w76_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid641_In1_c0 <= "" & bh7_w77_13_c0;
   bh7_w76_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1(0);
   bh7_w77_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1(1);
   bh7_w78_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid641: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid641_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid641_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid641_Out0_copy642_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid643_In0_c0 <= "" & bh7_w78_16_c0 & bh7_w78_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid643_In1_c0 <= "" & bh7_w79_13_c0;
   bh7_w78_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1(0);
   bh7_w79_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1(1);
   bh7_w80_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid643: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid643_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid643_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid643_Out0_copy644_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid645_In0_c0 <= "" & bh7_w80_16_c0 & bh7_w80_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid645_In1_c0 <= "" & bh7_w81_13_c0;
   bh7_w80_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1(0);
   bh7_w81_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1(1);
   bh7_w82_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid645: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid645_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid645_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid645_Out0_copy646_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid647_In0_c0 <= "" & bh7_w82_16_c0 & bh7_w82_15_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid647_In1_c0 <= "" & bh7_w83_13_c0;
   bh7_w82_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1(0);
   bh7_w83_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1(1);
   bh7_w84_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid647: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid647_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid647_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid647_Out0_copy648_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid649_In0_c0 <= "" & bh7_w84_15_c0 & bh7_w84_16_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid649_In1_c0 <= "" & bh7_w85_14_c0;
   bh7_w84_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1(0);
   bh7_w85_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1(1);
   bh7_w86_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid649: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid649_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid649_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid649_Out0_copy650_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid651_In0_c0 <= "" & bh7_w86_13_c0 & bh7_w86_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid651_In1_c0 <= "" & bh7_w87_15_c0;
   bh7_w86_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1(0);
   bh7_w87_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1(1);
   bh7_w88_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid651: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid651_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid651_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid651_Out0_copy652_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid653_In0_c0 <= "" & bh7_w88_13_c0 & bh7_w88_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid653_In1_c0 <= "" & bh7_w89_13_c0;
   bh7_w88_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1(0);
   bh7_w89_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1(1);
   bh7_w90_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid653: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid653_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid653_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid653_Out0_copy654_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid655_In0_c0 <= "" & bh7_w91_13_c0 & bh7_w91_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid655_In1_c0 <= "" & bh7_w92_13_c0;
   bh7_w91_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1(0);
   bh7_w92_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1(1);
   bh7_w93_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid655: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid655_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid655_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid655_Out0_copy656_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid657_In0_c0 <= "" & bh7_w94_13_c0 & bh7_w94_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid657_In1_c0 <= "" & bh7_w95_13_c0;
   bh7_w94_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1(0);
   bh7_w95_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1(1);
   bh7_w96_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid657: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid657_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid657_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid657_Out0_copy658_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid659_In0_c0 <= "" & bh7_w97_13_c0 & bh7_w97_14_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid659_In1_c0 <= "" & bh7_w98_13_c0;
   bh7_w97_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1(0);
   bh7_w98_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1(1);
   bh7_w99_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid659: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid659_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid659_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid659_Out0_copy660_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid661_In0_c0 <= "" & bh7_w100_10_c0 & bh7_w100_11_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid661_In1_c0 <= "" & bh7_w101_10_c0;
   bh7_w100_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1(0);
   bh7_w101_11_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1(1);
   bh7_w102_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid661: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid661_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid661_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid661_Out0_copy662_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid663_In0_c0 <= "" & bh7_w103_7_c0 & bh7_w103_8_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid663_In1_c0 <= "" & bh7_w104_4_c0;
   bh7_w103_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1(0);
   bh7_w104_5_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1(1);
   bh7_w105_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid663: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid663_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid663_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid663_Out0_copy664_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid665_In0_c0 <= "" & bh7_w105_5_c0 & bh7_w105_4_c0 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid665_In1_c0 <= "" & "0";
   bh7_w105_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_c1(0);
   Compressor_14_3_Freq300_uid326_uid665: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid665_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid665_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid665_Out0_copy666_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid667_In0_c0 <= "" & bh7_w17_0_c0 & bh7_w17_1_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid667_In1_c0 <= "" & bh7_w18_0_c0 & bh7_w18_1_c0;
   bh7_w17_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1(0);
   bh7_w18_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1(1);
   bh7_w19_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid667: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid667_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid667_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid667_Out0_copy668_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid669_In0_c0 <= "" & bh7_w19_0_c0 & bh7_w19_1_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid669_In1_c0 <= "" & bh7_w20_0_c0 & bh7_w20_1_c0;
   bh7_w19_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1(0);
   bh7_w20_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1(1);
   bh7_w21_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid669: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid669_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid669_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid669_Out0_copy670_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid671_In0_c0 <= "" & bh7_w21_0_c0 & bh7_w21_1_c0 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid671_In1_c0 <= "" & bh7_w22_0_c0 & bh7_w22_1_c0;
   bh7_w21_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1(0);
   bh7_w22_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1(1);
   bh7_w23_2_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid671: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid671_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid671_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid671_Out0_copy672_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid673_In0_c0 <= "" & bh7_w23_0_c0 & bh7_w23_1_c0 & "0";
   bh7_w23_3_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_c1(0);
   bh7_w24_3_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid673: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid673_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid673_Out0_copy674_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid675_In0_c0 <= "" & bh7_w24_0_c0 & bh7_w24_1_c0 & bh7_w24_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid675_In1_c0 <= "" & bh7_w25_0_c0 & bh7_w25_1_c0;
   bh7_w24_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1(0);
   bh7_w25_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1(1);
   bh7_w26_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid675: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid675_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid675_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid675_Out0_copy676_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid677_In0_c0 <= "" & bh7_w26_0_c0 & bh7_w26_1_c0 & bh7_w26_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid677_In1_c0 <= "" & bh7_w27_0_c0 & bh7_w27_1_c0;
   bh7_w26_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1(0);
   bh7_w27_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1(1);
   bh7_w28_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid677: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid677_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid677_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid677_Out0_copy678_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid679_In0_c0 <= "" & bh7_w28_0_c0 & bh7_w28_1_c0 & bh7_w28_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid679_In1_c0 <= "" & bh7_w29_0_c0 & bh7_w29_1_c0;
   bh7_w28_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1(0);
   bh7_w29_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1(1);
   bh7_w30_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid679: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid679_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid679_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid679_Out0_copy680_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid681_In0_c0 <= "" & bh7_w30_0_c0 & bh7_w30_1_c0 & bh7_w30_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid681_In1_c0 <= "" & bh7_w31_0_c0 & bh7_w31_1_c0;
   bh7_w30_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1(0);
   bh7_w31_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1(1);
   bh7_w32_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid681: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid681_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid681_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid681_Out0_copy682_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid683_In0_c0 <= "" & bh7_w32_0_c0 & bh7_w32_1_c0 & bh7_w32_2_c0;
   Compressor_23_3_Freq300_uid322_bh7_uid683_In1_c0 <= "" & bh7_w33_0_c0 & bh7_w33_1_c0;
   bh7_w32_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1(0);
   bh7_w33_3_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1(1);
   bh7_w34_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid683: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid683_In0_c0,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid683_In1_c0,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c0);
   Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid683_Out0_copy684_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid685_In0_c0 <= "" & bh7_w34_0_c0 & bh7_w34_1_c0 & bh7_w34_2_c0 & bh7_w34_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid685_In1_c0 <= "" & bh7_w35_0_c0;
   bh7_w34_5_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1(0);
   bh7_w35_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1(1);
   bh7_w36_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid685: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid685_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid685_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid685_Out0_copy686_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid687_In0_c0 <= "" & bh7_w35_1_c0 & bh7_w35_2_c0 & bh7_w35_3_c0;
   bh7_w35_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_c1(0);
   bh7_w36_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid687: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid687_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid687_Out0_copy688_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid689_In0_c0 <= "" & bh7_w36_0_c0 & bh7_w36_1_c0 & bh7_w36_2_c0 & bh7_w36_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid689_In1_c0 <= "" & bh7_w37_0_c0;
   bh7_w36_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1(0);
   bh7_w37_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1(1);
   bh7_w38_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid689: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid689_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid689_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid689_Out0_copy690_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid691_In0_c0 <= "" & bh7_w37_1_c0 & bh7_w37_2_c0 & bh7_w37_3_c0;
   bh7_w37_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_c1(0);
   bh7_w38_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid691: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid691_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid691_Out0_copy692_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid693_In0_c0 <= "" & bh7_w38_0_c0 & bh7_w38_1_c0 & bh7_w38_2_c0 & bh7_w38_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid693_In1_c0 <= "" & bh7_w39_0_c0;
   bh7_w38_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1(0);
   bh7_w39_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1(1);
   bh7_w40_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid693: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid693_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid693_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid693_Out0_copy694_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid695_In0_c0 <= "" & bh7_w39_1_c0 & bh7_w39_2_c0 & bh7_w39_3_c0;
   bh7_w39_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_c1(0);
   bh7_w40_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid695: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid695_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid695_Out0_copy696_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid697_In0_c0 <= "" & bh7_w40_0_c0 & bh7_w40_1_c0 & bh7_w40_2_c0 & bh7_w40_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid697_In1_c0 <= "" & bh7_w41_0_c0;
   bh7_w40_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1(0);
   bh7_w41_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1(1);
   bh7_w42_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid697: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid697_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid697_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid697_Out0_copy698_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid699_In0_c0 <= "" & bh7_w41_1_c0 & bh7_w41_2_c0 & bh7_w41_3_c0;
   bh7_w41_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_c1(0);
   bh7_w42_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid699: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid699_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid699_Out0_copy700_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid701_In0_c0 <= "" & bh7_w42_0_c0 & bh7_w42_1_c0 & bh7_w42_2_c0 & bh7_w42_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid701_In1_c0 <= "" & bh7_w43_0_c0;
   bh7_w42_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1(0);
   bh7_w43_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1(1);
   bh7_w44_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid701: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid701_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid701_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid701_Out0_copy702_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid703_In0_c0 <= "" & bh7_w43_1_c0 & bh7_w43_2_c0 & bh7_w43_3_c0;
   bh7_w43_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_c1(0);
   bh7_w44_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid703: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid703_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid703_Out0_copy704_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid705_In0_c0 <= "" & bh7_w44_0_c0 & bh7_w44_1_c0 & bh7_w44_2_c0 & bh7_w44_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid705_In1_c0 <= "" & bh7_w45_0_c0;
   bh7_w44_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1(0);
   bh7_w45_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1(1);
   bh7_w46_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid705: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid705_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid705_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid705_Out0_copy706_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid707_In0_c0 <= "" & bh7_w45_1_c0 & bh7_w45_2_c0 & bh7_w45_3_c0;
   bh7_w45_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_c1(0);
   bh7_w46_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid707: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid707_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid707_Out0_copy708_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid709_In0_c0 <= "" & bh7_w46_0_c0 & bh7_w46_1_c0 & bh7_w46_2_c0 & bh7_w46_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid709_In1_c0 <= "" & bh7_w47_0_c0;
   bh7_w46_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1(0);
   bh7_w47_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1(1);
   bh7_w48_5_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid709: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid709_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid709_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid709_Out0_copy710_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid711_In0_c0 <= "" & bh7_w47_1_c0 & bh7_w47_2_c0 & bh7_w47_3_c0;
   bh7_w47_5_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_c1(0);
   bh7_w48_6_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid711: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid711_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid711_Out0_copy712_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid713_In0_c0 <= "" & bh7_w48_4_c0 & bh7_w48_0_c0 & bh7_w48_1_c0 & bh7_w48_2_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid713_In1_c0 <= "" & bh7_w49_5_c0;
   bh7_w48_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1(0);
   bh7_w49_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1(1);
   bh7_w50_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid713: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid713_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid713_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid713_Out0_copy714_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid715_In0_c0 <= "" & bh7_w49_0_c0 & bh7_w49_1_c0 & bh7_w49_2_c0 & bh7_w49_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid715_In1_c0 <= "" & bh7_w50_6_c0;
   bh7_w49_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1(0);
   bh7_w50_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1(1);
   bh7_w51_11_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid715: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid715_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid715_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid715_Out0_copy716_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid717_In0_c0 <= "" & bh7_w50_0_c0 & bh7_w50_1_c0 & bh7_w50_2_c0 & bh7_w50_3_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid717_In1_c0 <= "" & bh7_w51_10_c0;
   bh7_w50_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1(0);
   bh7_w51_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1(1);
   bh7_w52_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid717: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid717_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid717_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid717_Out0_copy718_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid719_In0_c0 <= "" & bh7_w51_0_c0 & bh7_w51_1_c0 & bh7_w51_3_c0 & bh7_w51_4_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid719_In1_c0 <= "" & bh7_w52_11_c0;
   bh7_w51_13_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1(0);
   bh7_w52_13_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1(1);
   bh7_w53_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid719: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid719_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid719_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid719_Out0_copy720_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid721_In0_c0 <= "" & bh7_w52_0_c0 & bh7_w52_1_c0 & bh7_w52_3_c0 & bh7_w52_4_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid721_In1_c0 <= "" & bh7_w53_14_c0;
   bh7_w52_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1(0);
   bh7_w53_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1(1);
   bh7_w54_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid721: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid721_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid721_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid721_Out0_copy722_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid723_In0_c0 <= "" & bh7_w53_0_c0 & bh7_w53_1_c0 & bh7_w53_3_c0 & bh7_w53_4_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid723_In1_c0 <= "" & bh7_w54_15_c0;
   bh7_w53_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1(0);
   bh7_w54_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1(1);
   bh7_w55_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid723: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid723_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid723_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid723_Out0_copy724_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid725_In0_c0 <= "" & bh7_w54_0_c0 & bh7_w54_1_c0 & bh7_w54_4_c0 & bh7_w54_5_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid725_In1_c0 <= "" & bh7_w55_17_c0;
   bh7_w54_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1(0);
   bh7_w55_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1(1);
   bh7_w56_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid725: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid725_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid725_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid725_Out0_copy726_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid727_In0_c0 <= "" & bh7_w55_0_c0 & bh7_w55_1_c0 & bh7_w55_4_c0 & bh7_w55_5_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid727_In1_c0 <= "" & bh7_w56_15_c0;
   bh7_w55_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1(0);
   bh7_w56_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1(1);
   bh7_w57_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid727: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid727_In0_c0,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid727_In1_c0,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c0);
   Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid727_Out0_copy728_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c0 <= "" & bh7_w56_0_c0 & bh7_w56_1_c0 & bh7_w56_3_c0 & bh7_w56_4_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid729_In1_c1 <= "" & bh7_w57_20_c1;
   bh7_w56_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1(0);
   bh7_w57_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1(1);
   bh7_w58_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid729: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid729_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid729_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_copy730_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid729_Out0_copy730_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c0 <= "" & bh7_w57_0_c0 & bh7_w57_1_c0 & bh7_w57_4_c0 & bh7_w57_5_c0;
   Compressor_14_3_Freq300_uid326_bh7_uid731_In1_c1 <= "" & bh7_w58_19_c1;
   bh7_w57_23_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1(0);
   bh7_w58_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1(1);
   bh7_w59_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid731: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid731_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid731_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_copy732_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid731_Out0_copy732_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid733_In0_c0 <= "" & bh7_w58_0_c0 & bh7_w58_3_c0 & bh7_w58_4_c0;
   bh7_w58_22_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_c1(0);
   bh7_w59_19_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid733: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid733_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid733_Out0_copy734_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid735_In0_c1 <= "" & bh7_w59_16_c1 & bh7_w59_17_c1 & bh7_w59_0_c1 & bh7_w59_2_c1 & bh7_w59_3_c1 & bh7_w59_4_c1;
   bh7_w59_20_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1(0);
   bh7_w60_20_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1(1);
   bh7_w61_20_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1(2);
   Compressor_6_3_Freq300_uid334_uid735: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid735_In0_c1,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_copy736_c1);
   Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid735_Out0_copy736_c1; -- output copy to hold a pipeline register if needed


   Compressor_5_3_Freq300_uid400_bh7_uid737_In0_c1 <= "" & bh7_w60_19_c1 & bh7_w60_0_c1 & bh7_w60_3_c1 & bh7_w60_4_c1 & bh7_w60_5_c1;
   bh7_w60_21_c1 <= Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1(0);
   bh7_w61_21_c1 <= Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1(1);
   bh7_w62_17_c1 <= Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1(2);
   Compressor_5_3_Freq300_uid400_uid737: Compressor_5_3_Freq300_uid400
      port map ( X0 => Compressor_5_3_Freq300_uid400_bh7_uid737_In0_c1,
                 R => Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_copy738_c1);
   Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_c1 <= Compressor_5_3_Freq300_uid400_bh7_uid737_Out0_copy738_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid739_In0_c1 <= "" & bh7_w61_18_c1 & bh7_w61_19_c1 & bh7_w61_0_c1 & bh7_w61_3_c1 & bh7_w61_4_c1 & bh7_w61_5_c1;
   bh7_w61_22_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1(0);
   bh7_w62_18_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1(1);
   bh7_w63_20_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1(2);
   Compressor_6_3_Freq300_uid334_uid739: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid739_In0_c1,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_copy740_c1);
   Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid739_Out0_copy740_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid741_In0_c1 <= "" & bh7_w62_16_c1 & bh7_w62_0_c1 & bh7_w62_2_c1 & bh7_w62_3_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid741_In1_c1 <= "" & bh7_w63_19_c1;
   bh7_w62_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1(0);
   bh7_w63_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1(1);
   bh7_w64_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid741: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid741_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid741_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_copy742_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid741_Out0_copy742_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid743_In0_c0 <= "" & bh7_w63_0_c0 & bh7_w63_3_c0 & bh7_w63_4_c0;
   bh7_w63_22_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_c1(0);
   bh7_w64_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid743: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid743_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid743_Out0_copy744_c1; -- output copy to hold a pipeline register if needed


   Compressor_6_3_Freq300_uid334_bh7_uid745_In0_c1 <= "" & bh7_w64_18_c1 & bh7_w64_19_c1 & bh7_w64_0_c1 & bh7_w64_3_c1 & bh7_w64_4_c1 & bh7_w64_5_c1;
   bh7_w64_22_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1(0);
   bh7_w65_16_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1(1);
   bh7_w66_19_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1(2);
   Compressor_6_3_Freq300_uid334_uid745: Compressor_6_3_Freq300_uid334
      port map ( X0 => Compressor_6_3_Freq300_uid334_bh7_uid745_In0_c1,
                 R => Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_copy746_c1);
   Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_c1 <= Compressor_6_3_Freq300_uid334_bh7_uid745_Out0_copy746_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid747_In0_c1 <= "" & bh7_w65_15_c1 & bh7_w65_0_c1 & bh7_w65_2_c1 & bh7_w65_3_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid747_In1_c1 <= "" & bh7_w66_18_c1;
   bh7_w65_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1(0);
   bh7_w66_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1(1);
   bh7_w67_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid747: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid747_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid747_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_copy748_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid747_Out0_copy748_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid749_In0_c0 <= "" & bh7_w66_0_c0 & bh7_w66_3_c0 & bh7_w66_4_c0;
   bh7_w66_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_c1(0);
   bh7_w67_18_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid749: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid749_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid749_Out0_copy750_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid751_In0_c1 <= "" & bh7_w67_15_c1 & bh7_w67_16_c1 & bh7_w67_0_c1 & bh7_w67_3_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid751_In1_c1 <= "" & bh7_w68_19_c1;
   bh7_w67_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1(0);
   bh7_w68_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1(1);
   bh7_w69_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid751: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid751_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid751_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_copy752_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid751_Out0_copy752_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid753_In0_c0 <= "" & bh7_w68_0_c0 & bh7_w68_2_c0 & bh7_w68_3_c0;
   bh7_w68_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_c1(0);
   bh7_w69_17_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid753: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid753_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid753_Out0_copy754_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid755_In0_c1 <= "" & bh7_w69_15_c1 & bh7_w69_0_c1 & bh7_w69_3_c1 & bh7_w69_4_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid755_In1_c1 <= "" & bh7_w70_18_c1;
   bh7_w69_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1(0);
   bh7_w70_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1(1);
   bh7_w71_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid755: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid755_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid755_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_copy756_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid755_Out0_copy756_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid757_In0_c1 <= "" & bh7_w70_19_c1 & bh7_w70_0_c1 & bh7_w70_3_c1 & bh7_w70_4_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid757_In1_c1 <= "" & bh7_w71_15_c1;
   bh7_w70_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1(0);
   bh7_w71_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1(1);
   bh7_w72_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid757: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid757_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid757_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_copy758_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid757_Out0_copy758_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid759_In0_c0 <= "" & bh7_w71_0_c0 & bh7_w71_2_c0 & bh7_w71_3_c0;
   bh7_w71_18_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_c1(0);
   bh7_w72_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid759: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid759_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid759_Out0_copy760_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid761_In0_c1 <= "" & bh7_w72_18_c1 & bh7_w72_19_c1 & bh7_w72_0_c1 & bh7_w72_3_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid761_In1_c1 <= "" & bh7_w73_15_c1;
   bh7_w72_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1(0);
   bh7_w73_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1(1);
   bh7_w74_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid761: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid761_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid761_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_copy762_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid761_Out0_copy762_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid763_In0_c0 <= "" & bh7_w73_0_c0 & bh7_w73_3_c0 & bh7_w73_4_c0;
   bh7_w73_17_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_c1(0);
   bh7_w74_21_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid763: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid763_In0_c0,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c0);
   Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid763_Out0_copy764_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid765_In0_c1 <= "" & bh7_w74_18_c1 & bh7_w74_0_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c0 <= "" & bh7_w75_1_c0;
   bh7_w74_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1(0);
   bh7_w75_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1(1);
   bh7_w76_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid765: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid765_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid765_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_copy766_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid765_Out0_copy766_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid767_In0_c1 <= "" & bh7_w74_2_c1 & bh7_w74_3_c1 & bh7_w74_19_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid767_In1_c1 <= "" & bh7_w75_2_c1 & bh7_w75_14_c1;
   bh7_w74_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1(0);
   bh7_w75_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1(1);
   bh7_w76_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid767: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid767_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid767_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_copy768_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid767_Out0_copy768_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid769_In0_c1 <= "" & bh7_w76_1_c1 & bh7_w76_2_c1 & bh7_w76_18_c1 & bh7_w76_17_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c0 <= "" & "0";
   bh7_w76_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1(0);
   bh7_w77_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1(1);
   bh7_w78_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid769: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid769_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid769_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_copy770_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid769_Out0_copy770_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid771_In0_c1 <= "" & bh7_w77_0_c1 & bh7_w77_1_c1 & bh7_w77_14_c1;
   bh7_w77_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_c1(0);
   bh7_w78_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid771: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid771_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_copy772_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid771_Out0_copy772_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid773_In0_c1 <= "" & bh7_w78_0_c1 & bh7_w78_1_c1 & bh7_w78_18_c1 & bh7_w78_17_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c0 <= "" & "0";
   bh7_w78_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1(0);
   bh7_w79_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1(1);
   bh7_w80_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid773: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid773_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid773_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_copy774_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid773_Out0_copy774_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid775_In0_c1 <= "" & bh7_w79_0_c1 & bh7_w79_1_c1 & bh7_w79_14_c1;
   bh7_w79_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_c1(0);
   bh7_w80_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid775: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid775_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_copy776_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid775_Out0_copy776_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid777_In0_c1 <= "" & bh7_w80_0_c1 & bh7_w80_1_c1 & bh7_w80_18_c1 & bh7_w80_17_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c0 <= "" & "0";
   bh7_w80_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1(0);
   bh7_w81_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1(1);
   bh7_w82_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid777: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid777_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid777_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_copy778_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid777_Out0_copy778_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid779_In0_c1 <= "" & bh7_w81_0_c1 & bh7_w81_1_c1 & bh7_w81_14_c1;
   bh7_w81_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_c1(0);
   bh7_w82_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid779: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid779_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_copy780_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid779_Out0_copy780_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid781_In0_c1 <= "" & bh7_w82_18_c1 & bh7_w82_0_c1 & bh7_w82_17_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid781_In1_c1 <= "" & bh7_w83_14_c1 & bh7_w83_0_c1;
   bh7_w82_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1(0);
   bh7_w83_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1(1);
   bh7_w84_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid781: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid781_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid781_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_copy782_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid781_Out0_copy782_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid783_In0_c1 <= "" & bh7_w84_17_c1 & bh7_w84_18_c1 & bh7_w84_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid783_In1_c1 <= "" & bh7_w85_15_c1 & bh7_w85_0_c1;
   bh7_w84_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1(0);
   bh7_w85_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1(1);
   bh7_w86_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid783: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid783_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid783_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_copy784_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid783_Out0_copy784_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid785_In0_c1 <= "" & bh7_w86_15_c1 & bh7_w86_16_c1 & bh7_w86_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid785_In1_c1 <= "" & bh7_w87_16_c1 & bh7_w87_0_c1;
   bh7_w86_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1(0);
   bh7_w87_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1(1);
   bh7_w88_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid785: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid785_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid785_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_copy786_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid785_Out0_copy786_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid787_In0_c1 <= "" & bh7_w88_15_c1 & bh7_w88_16_c1 & bh7_w88_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid787_In1_c1 <= "" & bh7_w89_14_c1 & bh7_w89_0_c1;
   bh7_w88_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1(0);
   bh7_w89_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1(1);
   bh7_w90_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid787: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid787_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid787_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_copy788_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid787_Out0_copy788_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid789_In0_c1 <= "" & bh7_w90_15_c1 & bh7_w90_16_c1 & bh7_w90_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid789_In1_c1 <= "" & bh7_w91_15_c1 & bh7_w91_0_c1;
   bh7_w90_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1(0);
   bh7_w91_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1(1);
   bh7_w92_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid789: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid789_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid789_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_copy790_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid789_Out0_copy790_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid791_In0_c1 <= "" & bh7_w92_14_c1 & bh7_w92_0_c1 & "0";
   bh7_w92_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_c1(0);
   bh7_w93_17_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid791: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid791_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_copy792_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid791_Out0_copy792_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid793_In0_c1 <= "" & bh7_w93_15_c1 & bh7_w93_16_c1 & bh7_w93_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid793_In1_c1 <= "" & bh7_w94_15_c1 & bh7_w94_0_c1;
   bh7_w93_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1(0);
   bh7_w94_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1(1);
   bh7_w95_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid793: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid793_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid793_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_copy794_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid793_Out0_copy794_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid795_In0_c1 <= "" & bh7_w95_14_c1 & bh7_w95_0_c1 & "0";
   bh7_w95_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_c1(0);
   bh7_w96_17_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid795: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid795_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_copy796_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid795_Out0_copy796_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid797_In0_c1 <= "" & bh7_w96_15_c1 & bh7_w96_16_c1 & bh7_w96_0_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid797_In1_c1 <= "" & bh7_w97_15_c1 & bh7_w97_0_c1;
   bh7_w96_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1(0);
   bh7_w97_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1(1);
   bh7_w98_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid797: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid797_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid797_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_copy798_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid797_Out0_copy798_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid799_In0_c1 <= "" & bh7_w98_14_c1 & bh7_w98_0_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid799_In1_c1 <= "" & bh7_w99_14_c1 & bh7_w99_15_c1;
   bh7_w98_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1(0);
   bh7_w99_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1(1);
   bh7_w100_13_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid799: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid799_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid799_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_copy800_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid799_Out0_copy800_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid801_In0_c1 <= "" & bh7_w102_9_c1 & bh7_w102_10_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid801_In1_c1 <= "" & bh7_w103_9_c1;
   bh7_w102_11_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1(0);
   bh7_w103_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1(1);
   bh7_w104_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid801: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid801_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid801_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_copy802_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid801_Out0_copy802_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid803_In0_c1 <= "" & bh7_w105_6_c1 & bh7_w105_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c0 <= "" & "0";
   bh7_w105_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_c1(0);
   Compressor_14_3_Freq300_uid326_uid803: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid803_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid803_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_copy804_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid803_Out0_copy804_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid805_In0_c1 <= "" & bh7_w19_3_c1 & bh7_w19_2_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid805_In1_c1 <= "" & bh7_w20_2_c1;
   bh7_w19_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1(0);
   bh7_w20_3_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1(1);
   bh7_w21_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid805: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid805_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid805_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_copy806_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid805_Out0_copy806_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid807_In0_c1 <= "" & bh7_w21_3_c1 & bh7_w21_2_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid807_In1_c1 <= "" & bh7_w22_2_c1;
   bh7_w21_5_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1(0);
   bh7_w22_3_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1(1);
   bh7_w23_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid807: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid807_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid807_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_copy808_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid807_Out0_copy808_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid809_In0_c1 <= "" & bh7_w23_3_c1 & bh7_w23_2_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid809_In1_c1 <= "" & bh7_w24_4_c1 & bh7_w24_3_c1;
   bh7_w23_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1(0);
   bh7_w24_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1(1);
   bh7_w25_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid809: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid809_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid809_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_copy810_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid809_Out0_copy810_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid811_In0_c1 <= "" & bh7_w25_2_c1 & bh7_w25_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid811_In1_c1 <= "" & bh7_w26_4_c1 & bh7_w26_3_c1;
   bh7_w25_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1(0);
   bh7_w26_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1(1);
   bh7_w27_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid811: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid811_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid811_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_copy812_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid811_Out0_copy812_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid813_In0_c1 <= "" & bh7_w27_2_c1 & bh7_w27_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid813_In1_c1 <= "" & bh7_w28_4_c1 & bh7_w28_3_c1;
   bh7_w27_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1(0);
   bh7_w28_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1(1);
   bh7_w29_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid813: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid813_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid813_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_copy814_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid813_Out0_copy814_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid815_In0_c1 <= "" & bh7_w29_2_c1 & bh7_w29_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid815_In1_c1 <= "" & bh7_w30_4_c1 & bh7_w30_3_c1;
   bh7_w29_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1(0);
   bh7_w30_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1(1);
   bh7_w31_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid815: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid815_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid815_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_copy816_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid815_Out0_copy816_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid817_In0_c1 <= "" & bh7_w31_2_c1 & bh7_w31_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid817_In1_c1 <= "" & bh7_w32_4_c1 & bh7_w32_3_c1;
   bh7_w31_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1(0);
   bh7_w32_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1(1);
   bh7_w33_4_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid817: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid817_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid817_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_copy818_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid817_Out0_copy818_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid819_In0_c1 <= "" & bh7_w33_2_c1 & bh7_w33_3_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid819_In1_c1 <= "" & bh7_w34_5_c1 & bh7_w34_4_c1;
   bh7_w33_5_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1(0);
   bh7_w34_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1(1);
   bh7_w35_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid819: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid819_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid819_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_copy820_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid819_Out0_copy820_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid821_In0_c1 <= "" & bh7_w35_5_c1 & bh7_w35_4_c1 & "0";
   bh7_w35_7_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_c1(0);
   bh7_w36_7_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid821: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid821_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_copy822_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid821_Out0_copy822_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid823_In0_c1 <= "" & bh7_w36_6_c1 & bh7_w36_5_c1 & bh7_w36_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid823_In1_c1 <= "" & bh7_w37_5_c1 & bh7_w37_4_c1;
   bh7_w36_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1(0);
   bh7_w37_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1(1);
   bh7_w38_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid823: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid823_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid823_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_copy824_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid823_Out0_copy824_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid825_In0_c1 <= "" & bh7_w38_6_c1 & bh7_w38_5_c1 & bh7_w38_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid825_In1_c1 <= "" & bh7_w39_5_c1 & bh7_w39_4_c1;
   bh7_w38_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1(0);
   bh7_w39_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1(1);
   bh7_w40_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid825: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid825_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid825_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_copy826_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid825_Out0_copy826_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid827_In0_c1 <= "" & bh7_w40_6_c1 & bh7_w40_5_c1 & bh7_w40_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid827_In1_c1 <= "" & bh7_w41_5_c1 & bh7_w41_4_c1;
   bh7_w40_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1(0);
   bh7_w41_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1(1);
   bh7_w42_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid827: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid827_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid827_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_copy828_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid827_Out0_copy828_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid829_In0_c1 <= "" & bh7_w42_6_c1 & bh7_w42_5_c1 & bh7_w42_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid829_In1_c1 <= "" & bh7_w43_5_c1 & bh7_w43_4_c1;
   bh7_w42_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1(0);
   bh7_w43_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1(1);
   bh7_w44_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid829: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid829_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid829_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_copy830_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid829_Out0_copy830_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid831_In0_c1 <= "" & bh7_w44_6_c1 & bh7_w44_5_c1 & bh7_w44_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid831_In1_c1 <= "" & bh7_w45_5_c1 & bh7_w45_4_c1;
   bh7_w44_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1(0);
   bh7_w45_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1(1);
   bh7_w46_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid831: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid831_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid831_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_copy832_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid831_Out0_copy832_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid833_In0_c1 <= "" & bh7_w46_6_c1 & bh7_w46_5_c1 & bh7_w46_4_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid833_In1_c1 <= "" & bh7_w47_5_c1 & bh7_w47_4_c1;
   bh7_w46_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1(0);
   bh7_w47_6_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1(1);
   bh7_w48_8_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid833: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid833_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid833_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_copy834_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid833_Out0_copy834_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid835_In0_c1 <= "" & bh7_w48_3_c1 & bh7_w48_7_c1 & bh7_w48_6_c1 & bh7_w48_5_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid835_In1_c1 <= "" & bh7_w49_7_c1;
   bh7_w48_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1(0);
   bh7_w49_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1(1);
   bh7_w50_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid835: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid835_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid835_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_copy836_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid835_Out0_copy836_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid837_In0_c1 <= "" & bh7_w50_9_c1 & bh7_w50_8_c1 & bh7_w50_7_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid837_In1_c1 <= "" & bh7_w51_13_c1 & bh7_w51_12_c1;
   bh7_w50_11_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1(0);
   bh7_w51_14_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1(1);
   bh7_w52_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid837: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid837_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid837_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_copy838_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid837_Out0_copy838_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid839_In0_c1 <= "" & bh7_w52_14_c1 & bh7_w52_13_c1 & bh7_w52_12_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid839_In1_c1 <= "" & bh7_w53_17_c1 & bh7_w53_16_c1;
   bh7_w52_16_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1(0);
   bh7_w53_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1(1);
   bh7_w54_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid839: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid839_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid839_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_copy840_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid839_Out0_copy840_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid841_In0_c1 <= "" & bh7_w54_18_c1 & bh7_w54_17_c1 & bh7_w54_16_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid841_In1_c1 <= "" & bh7_w55_19_c1 & bh7_w55_20_c1;
   bh7_w54_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1(0);
   bh7_w55_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1(1);
   bh7_w56_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid841: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid841_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid841_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_copy842_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid841_Out0_copy842_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid843_In0_c1 <= "" & bh7_w56_16_c1 & bh7_w56_17_c1 & bh7_w56_18_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid843_In1_c1 <= "" & bh7_w57_21_c1 & bh7_w57_22_c1;
   bh7_w56_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1(0);
   bh7_w57_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1(1);
   bh7_w58_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid843: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid843_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid843_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_copy844_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid843_Out0_copy844_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid845_In0_c1 <= "" & bh7_w58_20_c1 & bh7_w58_21_c1 & bh7_w58_5_c1 & bh7_w58_22_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c0 <= "" & "0";
   bh7_w58_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1(0);
   bh7_w59_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1(1);
   bh7_w60_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid845: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid845_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid845_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_copy846_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid845_Out0_copy846_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid847_In0_c1 <= "" & bh7_w59_18_c1 & bh7_w59_20_c1 & bh7_w59_19_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid847_In1_c1 <= "" & bh7_w60_20_c1 & bh7_w60_21_c1;
   bh7_w59_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1(0);
   bh7_w60_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1(1);
   bh7_w61_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid847: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid847_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid847_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_copy848_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid847_Out0_copy848_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid849_In0_c1 <= "" & bh7_w61_20_c1 & bh7_w61_21_c1 & bh7_w61_22_c1;
   bh7_w61_24_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_c1(0);
   bh7_w62_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid849: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid849_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_copy850_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid849_Out0_copy850_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid851_In0_c1 <= "" & bh7_w62_17_c1 & bh7_w62_18_c1 & bh7_w62_19_c1 & bh7_w62_4_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid851_In1_c1 <= "" & bh7_w63_20_c1;
   bh7_w62_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1(0);
   bh7_w63_23_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1(1);
   bh7_w64_23_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid851: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid851_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid851_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_copy852_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid851_Out0_copy852_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid853_In0_c1 <= "" & bh7_w63_21_c1 & bh7_w63_5_c1 & bh7_w63_22_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c0 <= "" & "0" & "0";
   bh7_w63_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1(0);
   bh7_w64_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1(1);
   bh7_w65_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid853: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid853_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid853_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_copy854_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid853_Out0_copy854_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid855_In0_c1 <= "" & bh7_w64_20_c1 & bh7_w64_22_c1 & bh7_w64_21_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid855_In1_c1 <= "" & bh7_w65_16_c1 & bh7_w65_17_c1;
   bh7_w64_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1(0);
   bh7_w65_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1(1);
   bh7_w66_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid855: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid855_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid855_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_copy856_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid855_Out0_copy856_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid857_In0_c1 <= "" & bh7_w66_19_c1 & bh7_w66_20_c1 & bh7_w66_21_c1;
   bh7_w66_23_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_c1(0);
   bh7_w67_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid857: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid857_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_copy858_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid857_Out0_copy858_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid859_In0_c1 <= "" & bh7_w67_17_c1 & bh7_w67_19_c1 & bh7_w67_4_c1 & bh7_w67_18_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid859_In1_c1 <= "" & bh7_w68_20_c1;
   bh7_w67_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1(0);
   bh7_w68_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1(1);
   bh7_w69_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid859: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid859_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid859_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_copy860_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid859_Out0_copy860_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid861_In0_c1 <= "" & bh7_w69_16_c1 & bh7_w69_18_c1 & bh7_w69_17_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid861_In1_c1 <= "" & bh7_w70_20_c1 & bh7_w70_21_c1;
   bh7_w69_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1(0);
   bh7_w70_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1(1);
   bh7_w71_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid861: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid861_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid861_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_copy862_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid861_Out0_copy862_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid863_In0_c1 <= "" & bh7_w71_16_c1 & bh7_w71_17_c1 & bh7_w71_18_c1;
   bh7_w71_20_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_c1(0);
   bh7_w72_23_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid863: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid863_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_copy864_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid863_Out0_copy864_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid865_In0_c1 <= "" & bh7_w72_20_c1 & bh7_w72_22_c1 & bh7_w72_4_c1 & bh7_w72_21_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid865_In1_c1 <= "" & bh7_w73_16_c1;
   bh7_w72_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1(0);
   bh7_w73_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1(1);
   bh7_w74_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid865: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid865_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid865_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_copy866_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid865_Out0_copy866_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid867_In0_c1 <= "" & bh7_w74_20_c1 & bh7_w74_22_c1 & bh7_w74_21_c1 & bh7_w74_23_c1;
   Compressor_14_3_Freq300_uid326_bh7_uid867_In1_c1 <= "" & bh7_w75_15_c1;
   bh7_w74_25_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1(0);
   bh7_w75_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1(1);
   bh7_w76_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid867: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid867_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid867_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_copy868_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid867_Out0_copy868_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid869_In0_c1 <= "" & bh7_w76_19_c1 & bh7_w76_21_c1 & bh7_w76_20_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid869_In1_c1 <= "" & bh7_w77_15_c1 & bh7_w77_16_c1;
   bh7_w76_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1(0);
   bh7_w77_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1(1);
   bh7_w78_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid869: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid869_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid869_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_copy870_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid869_Out0_copy870_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid871_In0_c1 <= "" & bh7_w78_19_c1 & bh7_w78_21_c1 & bh7_w78_20_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid871_In1_c1 <= "" & bh7_w79_15_c1 & bh7_w79_16_c1;
   bh7_w78_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1(0);
   bh7_w79_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1(1);
   bh7_w80_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid871: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid871_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid871_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_copy872_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid871_Out0_copy872_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid873_In0_c1 <= "" & bh7_w80_19_c1 & bh7_w80_21_c1 & bh7_w80_20_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid873_In1_c1 <= "" & bh7_w81_15_c1 & bh7_w81_16_c1;
   bh7_w80_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1(0);
   bh7_w81_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1(1);
   bh7_w82_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid873: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid873_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid873_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_copy874_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid873_Out0_copy874_c1; -- output copy to hold a pipeline register if needed


   Compressor_3_2_Freq300_uid432_bh7_uid875_In0_c1 <= "" & bh7_w82_19_c1 & bh7_w82_21_c1 & bh7_w82_20_c1;
   bh7_w82_23_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_c1(0);
   bh7_w83_16_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_c1(1);
   Compressor_3_2_Freq300_uid432_uid875: Compressor_3_2_Freq300_uid432
      port map ( X0 => Compressor_3_2_Freq300_uid432_bh7_uid875_In0_c1,
                 R => Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_copy876_c1);
   Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_c1 <= Compressor_3_2_Freq300_uid432_bh7_uid875_Out0_copy876_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid877_In0_c1 <= "" & bh7_w84_19_c1 & bh7_w84_20_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid877_In1_c1 <= "" & bh7_w85_16_c1;
   bh7_w84_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1(0);
   bh7_w85_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1(1);
   bh7_w86_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid877: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid877_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid877_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_copy878_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid877_Out0_copy878_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid879_In0_c1 <= "" & bh7_w86_17_c1 & bh7_w86_18_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid879_In1_c1 <= "" & bh7_w87_17_c1;
   bh7_w86_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1(0);
   bh7_w87_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1(1);
   bh7_w88_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid879: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid879_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid879_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_copy880_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid879_Out0_copy880_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid881_In0_c1 <= "" & bh7_w88_17_c1 & bh7_w88_18_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid881_In1_c1 <= "" & bh7_w89_15_c1;
   bh7_w88_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1(0);
   bh7_w89_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1(1);
   bh7_w90_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid881: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid881_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid881_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_copy882_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid881_Out0_copy882_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid883_In0_c1 <= "" & bh7_w90_17_c1 & bh7_w90_18_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid883_In1_c1 <= "" & bh7_w91_16_c1;
   bh7_w90_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1(0);
   bh7_w91_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1(1);
   bh7_w92_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid883: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid883_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid883_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_copy884_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid883_Out0_copy884_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid885_In0_c1 <= "" & bh7_w92_15_c1 & bh7_w92_16_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid885_In1_c1 <= "" & bh7_w93_17_c1 & bh7_w93_18_c1;
   bh7_w92_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1(0);
   bh7_w93_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1(1);
   bh7_w94_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid885: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid885_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid885_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_copy886_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid885_Out0_copy886_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid887_In0_c1 <= "" & bh7_w95_15_c1 & bh7_w95_16_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid887_In1_c1 <= "" & bh7_w96_17_c1 & bh7_w96_18_c1;
   bh7_w95_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1(0);
   bh7_w96_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1(1);
   bh7_w97_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid887: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid887_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid887_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_copy888_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid887_Out0_copy888_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid889_In0_c1 <= "" & bh7_w98_15_c1 & bh7_w98_16_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid889_In1_c1 <= "" & bh7_w99_16_c1;
   bh7_w98_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1(0);
   bh7_w99_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1(1);
   bh7_w100_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid889: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid889_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid889_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_copy890_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid889_Out0_copy890_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid891_In0_c1 <= "" & bh7_w100_12_c1 & bh7_w100_13_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid891_In1_c1 <= "" & bh7_w101_11_c1;
   bh7_w100_15_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1(0);
   bh7_w101_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1(1);
   bh7_w102_12_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid891: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid891_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid891_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_copy892_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid891_Out0_copy892_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid893_In0_c1 <= "" & bh7_w104_5_c1 & bh7_w104_6_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid893_In1_c1 <= "" & bh7_w105_8_c1;
   bh7_w104_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_c1(0);
   bh7_w105_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_c1(1);
   Compressor_14_3_Freq300_uid326_uid893: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid893_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid893_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_copy894_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid893_Out0_copy894_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid895_In0_c1 <= "" & bh7_w21_5_c1 & bh7_w21_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid895_In1_c1 <= "" & bh7_w22_3_c1;
   bh7_w21_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1(0);
   bh7_w22_4_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1(1);
   bh7_w23_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid895: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid895_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid895_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_copy896_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid895_Out0_copy896_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid897_In0_c1 <= "" & bh7_w23_5_c1 & bh7_w23_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid897_In1_c1 <= "" & bh7_w24_5_c1;
   bh7_w23_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1(0);
   bh7_w24_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1(1);
   bh7_w25_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid897: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid897_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid897_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_copy898_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid897_Out0_copy898_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid899_In0_c1 <= "" & bh7_w25_5_c1 & bh7_w25_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid899_In1_c1 <= "" & bh7_w26_5_c1;
   bh7_w25_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1(0);
   bh7_w26_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1(1);
   bh7_w27_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid899: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid899_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid899_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_copy900_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid899_Out0_copy900_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid901_In0_c1 <= "" & bh7_w27_5_c1 & bh7_w27_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid901_In1_c1 <= "" & bh7_w28_5_c1;
   bh7_w27_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1(0);
   bh7_w28_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1(1);
   bh7_w29_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid901: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid901_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid901_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_copy902_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid901_Out0_copy902_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid903_In0_c1 <= "" & bh7_w29_5_c1 & bh7_w29_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid903_In1_c1 <= "" & bh7_w30_5_c1;
   bh7_w29_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1(0);
   bh7_w30_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1(1);
   bh7_w31_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid903: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid903_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid903_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_copy904_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid903_Out0_copy904_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid905_In0_c1 <= "" & bh7_w31_5_c1 & bh7_w31_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid905_In1_c1 <= "" & bh7_w32_5_c1;
   bh7_w31_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1(0);
   bh7_w32_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1(1);
   bh7_w33_6_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid905: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid905_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid905_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_copy906_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid905_Out0_copy906_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid907_In0_c1 <= "" & bh7_w33_5_c1 & bh7_w33_4_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid907_In1_c1 <= "" & bh7_w34_6_c1;
   bh7_w33_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1(0);
   bh7_w34_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1(1);
   bh7_w35_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid907: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid907_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid907_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_copy908_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid907_Out0_copy908_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid909_In0_c1 <= "" & bh7_w35_7_c1 & bh7_w35_6_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid909_In1_c1 <= "" & bh7_w36_8_c1 & bh7_w36_7_c1;
   bh7_w35_9_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1(0);
   bh7_w36_9_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1(1);
   bh7_w37_7_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid909: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid909_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid909_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_copy910_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid909_Out0_copy910_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid911_In0_c1 <= "" & bh7_w38_8_c1 & bh7_w38_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid911_In1_c1 <= "" & bh7_w39_6_c1;
   bh7_w38_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1(0);
   bh7_w39_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1(1);
   bh7_w40_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid911: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid911_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid911_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_copy912_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid911_Out0_copy912_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid913_In0_c1 <= "" & bh7_w40_8_c1 & bh7_w40_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid913_In1_c1 <= "" & bh7_w41_6_c1;
   bh7_w40_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1(0);
   bh7_w41_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1(1);
   bh7_w42_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid913: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid913_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid913_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_copy914_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid913_Out0_copy914_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid915_In0_c1 <= "" & bh7_w42_8_c1 & bh7_w42_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid915_In1_c1 <= "" & bh7_w43_6_c1;
   bh7_w42_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1(0);
   bh7_w43_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1(1);
   bh7_w44_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid915: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid915_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid915_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_copy916_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid915_Out0_copy916_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid917_In0_c1 <= "" & bh7_w44_8_c1 & bh7_w44_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid917_In1_c1 <= "" & bh7_w45_6_c1;
   bh7_w44_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1(0);
   bh7_w45_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1(1);
   bh7_w46_9_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid917: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid917_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid917_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_copy918_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid917_Out0_copy918_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid919_In0_c1 <= "" & bh7_w46_8_c1 & bh7_w46_7_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid919_In1_c1 <= "" & bh7_w47_6_c1;
   bh7_w46_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1(0);
   bh7_w47_7_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1(1);
   bh7_w48_10_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid919: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid919_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid919_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_copy920_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid919_Out0_copy920_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid921_In0_c1 <= "" & bh7_w48_9_c1 & bh7_w48_8_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid921_In1_c1 <= "" & bh7_w49_6_c1 & bh7_w49_8_c1;
   bh7_w48_11_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1(0);
   bh7_w49_9_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1(1);
   bh7_w50_12_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid921: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid921_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid921_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_copy922_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid921_Out0_copy922_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid923_In0_c1 <= "" & bh7_w50_11_c1 & bh7_w50_10_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid923_In1_c1 <= "" & bh7_w51_11_c1 & bh7_w51_14_c1;
   bh7_w50_13_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1(0);
   bh7_w51_15_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1(1);
   bh7_w52_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid923: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid923_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid923_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_copy924_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid923_Out0_copy924_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid925_In0_c1 <= "" & bh7_w52_16_c1 & bh7_w52_15_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid925_In1_c1 <= "" & bh7_w53_15_c1 & bh7_w53_18_c1;
   bh7_w52_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1(0);
   bh7_w53_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1(1);
   bh7_w54_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid925: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid925_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid925_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_copy926_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid925_Out0_copy926_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid927_In0_c1 <= "" & bh7_w54_20_c1 & bh7_w54_19_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid927_In1_c1 <= "" & bh7_w55_21_c1 & bh7_w55_18_c1;
   bh7_w54_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1(0);
   bh7_w55_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1(1);
   bh7_w56_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid927: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid927_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid927_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_copy928_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid927_Out0_copy928_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid929_In0_c1 <= "" & bh7_w56_19_c1 & bh7_w56_20_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid929_In1_c1 <= "" & bh7_w57_23_c1 & bh7_w57_24_c1;
   bh7_w56_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1(0);
   bh7_w57_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1(1);
   bh7_w58_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid929: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid929_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid929_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_copy930_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid929_Out0_copy930_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid931_In0_c1 <= "" & bh7_w58_23_c1 & bh7_w58_24_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid931_In1_c1 <= "" & bh7_w59_21_c1 & bh7_w59_22_c1;
   bh7_w58_26_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1(0);
   bh7_w59_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1(1);
   bh7_w60_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid931: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid931_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid931_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_copy932_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid931_Out0_copy932_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid933_In0_c1 <= "" & bh7_w60_22_c1 & bh7_w60_23_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid933_In1_c1 <= "" & bh7_w61_23_c1 & bh7_w61_24_c1;
   bh7_w60_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1(0);
   bh7_w61_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1(1);
   bh7_w62_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid933: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid933_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid933_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_copy934_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid933_Out0_copy934_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid935_In0_c1 <= "" & bh7_w62_20_c1 & bh7_w62_21_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid935_In1_c1 <= "" & bh7_w63_23_c1 & bh7_w63_24_c1;
   bh7_w62_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1(0);
   bh7_w63_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1(1);
   bh7_w64_26_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid935: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid935_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid935_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_copy936_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid935_Out0_copy936_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid937_In0_c1 <= "" & bh7_w64_23_c1 & bh7_w64_24_c1 & bh7_w64_25_c1;
   Compressor_23_3_Freq300_uid322_bh7_uid937_In1_c1 <= "" & bh7_w65_18_c1 & bh7_w65_19_c1;
   bh7_w64_27_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1(0);
   bh7_w65_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1(1);
   bh7_w66_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid937: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid937_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid937_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_copy938_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid937_Out0_copy938_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid939_In0_c1 <= "" & bh7_w66_22_c1 & bh7_w66_23_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid939_In1_c1 <= "" & bh7_w67_20_c1 & bh7_w67_21_c1;
   bh7_w66_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1(0);
   bh7_w67_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1(1);
   bh7_w68_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid939: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid939_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid939_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_copy940_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid939_Out0_copy940_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid941_In0_c1 <= "" & bh7_w68_22_c1 & bh7_w68_21_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid941_In1_c1 <= "" & bh7_w69_19_c1 & bh7_w69_20_c1;
   bh7_w68_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1(0);
   bh7_w69_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1(1);
   bh7_w70_23_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid941: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid941_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid941_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_copy942_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid941_Out0_copy942_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid943_In0_c1 <= "" & bh7_w71_19_c1 & bh7_w71_20_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid943_In1_c1 <= "" & bh7_w72_23_c1 & bh7_w72_24_c1;
   bh7_w71_21_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1(0);
   bh7_w72_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1(1);
   bh7_w73_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid943: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid943_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid943_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_copy944_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid943_Out0_copy944_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid945_In0_c1 <= "" & bh7_w73_18_c1 & bh7_w73_17_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid945_In1_c1 <= "" & bh7_w74_24_c1 & bh7_w74_25_c1;
   bh7_w73_20_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1(0);
   bh7_w74_26_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1(1);
   bh7_w75_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid945: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid945_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid945_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_copy946_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid945_Out0_copy946_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid947_In0_c1 <= "" & bh7_w75_17_c1 & bh7_w75_16_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid947_In1_c1 <= "" & bh7_w76_22_c1 & bh7_w76_23_c1;
   bh7_w75_19_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1(0);
   bh7_w76_24_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1(1);
   bh7_w77_18_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid947: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid947_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid947_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_copy948_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid947_Out0_copy948_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid949_In0_c1 <= "" & bh7_w78_22_c1 & bh7_w78_23_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid949_In1_c1 <= "" & bh7_w79_17_c1;
   bh7_w78_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1(0);
   bh7_w79_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1(1);
   bh7_w80_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid949: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid949_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid949_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_copy950_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid949_Out0_copy950_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid951_In0_c1 <= "" & bh7_w80_22_c1 & bh7_w80_23_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid951_In1_c1 <= "" & bh7_w81_17_c1;
   bh7_w80_25_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1(0);
   bh7_w81_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1(1);
   bh7_w82_24_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid951: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid951_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid951_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_copy952_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid951_Out0_copy952_c1; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq300_uid322_bh7_uid953_In0_c1 <= "" & bh7_w82_22_c1 & bh7_w82_23_c1 & "0";
   Compressor_23_3_Freq300_uid322_bh7_uid953_In1_c1 <= "" & bh7_w83_15_c1 & bh7_w83_16_c1;
   bh7_w82_25_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1(0);
   bh7_w83_17_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1(1);
   bh7_w84_22_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1(2);
   Compressor_23_3_Freq300_uid322_uid953: Compressor_23_3_Freq300_uid322
      port map ( X0 => Compressor_23_3_Freq300_uid322_bh7_uid953_In0_c1,
                 X1 => Compressor_23_3_Freq300_uid322_bh7_uid953_In1_c1,
                 R => Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_copy954_c1);
   Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_c1 <= Compressor_23_3_Freq300_uid322_bh7_uid953_Out0_copy954_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid955_In0_c1 <= "" & bh7_w86_19_c1 & bh7_w86_20_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid955_In1_c1 <= "" & bh7_w87_18_c1;
   bh7_w86_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1(0);
   bh7_w87_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1(1);
   bh7_w88_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid955: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid955_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid955_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_copy956_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid955_Out0_copy956_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid957_In0_c1 <= "" & bh7_w88_19_c1 & bh7_w88_20_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid957_In1_c1 <= "" & bh7_w89_16_c1;
   bh7_w88_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1(0);
   bh7_w89_17_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1(1);
   bh7_w90_21_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid957: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid957_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid957_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_copy958_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid957_Out0_copy958_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid959_In0_c1 <= "" & bh7_w90_19_c1 & bh7_w90_20_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid959_In1_c1 <= "" & bh7_w91_17_c1;
   bh7_w90_22_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1(0);
   bh7_w91_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1(1);
   bh7_w92_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid959: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid959_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid959_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_copy960_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid959_Out0_copy960_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid961_In0_c1 <= "" & bh7_w92_17_c1 & bh7_w92_18_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid961_In1_c1 <= "" & bh7_w93_19_c1;
   bh7_w92_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1(0);
   bh7_w93_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1(1);
   bh7_w94_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid961: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid961_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid961_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_copy962_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid961_Out0_copy962_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid963_In0_c1 <= "" & bh7_w94_16_c1 & bh7_w94_17_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid963_In1_c1 <= "" & bh7_w95_17_c1;
   bh7_w94_19_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1(0);
   bh7_w95_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1(1);
   bh7_w96_20_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid963: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid963_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid963_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_copy964_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid963_Out0_copy964_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid965_In0_c1 <= "" & bh7_w97_16_c1 & bh7_w97_17_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid965_In1_c1 <= "" & bh7_w98_17_c1;
   bh7_w97_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1(0);
   bh7_w98_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1(1);
   bh7_w99_18_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid965: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid965_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid965_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_copy966_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid965_Out0_copy966_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid967_In0_c1 <= "" & bh7_w100_14_c1 & bh7_w100_15_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid967_In1_c1 <= "" & bh7_w101_12_c1;
   bh7_w100_16_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1(0);
   bh7_w101_13_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1(1);
   bh7_w102_13_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid967: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid967_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid967_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_copy968_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid967_Out0_copy968_c1; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq300_uid326_bh7_uid969_In0_c1 <= "" & bh7_w102_11_c1 & bh7_w102_12_c1 & "0" & "0";
   Compressor_14_3_Freq300_uid326_bh7_uid969_In1_c1 <= "" & bh7_w103_10_c1;
   bh7_w102_14_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1(0);
   bh7_w103_11_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1(1);
   bh7_w104_8_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1(2);
   Compressor_14_3_Freq300_uid326_uid969: Compressor_14_3_Freq300_uid326
      port map ( X0 => Compressor_14_3_Freq300_uid326_bh7_uid969_In0_c1,
                 X1 => Compressor_14_3_Freq300_uid326_bh7_uid969_In1_c1,
                 R => Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_copy970_c1);
   Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_c1 <= Compressor_14_3_Freq300_uid326_bh7_uid969_Out0_copy970_c1; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh7_22_c1 <= bh7_w22_4_c1 & bh7_w21_6_c1 & bh7_w20_3_c1 & bh7_w19_4_c1 & bh7_w18_2_c1 & bh7_w17_2_c1 & bh7_w16_0_c1 & bh7_w15_0_c1 & bh7_w14_0_c1 & bh7_w13_0_c1 & bh7_w12_0_c1 & bh7_w11_0_c1 & bh7_w10_0_c1 & bh7_w9_0_c1 & bh7_w8_0_c1 & bh7_w7_0_c1 & bh7_w6_0_c1 & bh7_w5_0_c1 & bh7_w4_0_c1 & bh7_w3_0_c1 & bh7_w2_0_c1 & bh7_w1_0_c1 & bh7_w0_0_c1;

   bitheapFinalAdd_bh7_In0_c1 <= "0" & bh7_w105_9_c1 & bh7_w104_7_c1 & bh7_w103_11_c1 & bh7_w102_13_c1 & bh7_w101_13_c1 & bh7_w100_16_c1 & bh7_w99_17_c1 & bh7_w98_18_c1 & bh7_w97_18_c1 & bh7_w96_19_c1 & bh7_w95_18_c1 & bh7_w94_18_c1 & bh7_w93_20_c1 & bh7_w92_19_c1 & bh7_w91_18_c1 & bh7_w90_21_c1 & bh7_w89_17_c1 & bh7_w88_21_c1 & bh7_w87_19_c1 & bh7_w86_21_c1 & bh7_w85_17_c1 & bh7_w84_21_c1 & bh7_w83_17_c1 & bh7_w82_24_c1 & bh7_w81_18_c1 & bh7_w80_24_c1 & bh7_w79_18_c1 & bh7_w78_24_c1 & bh7_w77_17_c1 & bh7_w76_24_c1 & bh7_w75_18_c1 & bh7_w74_26_c1 & bh7_w73_19_c1 & bh7_w72_25_c1 & bh7_w71_21_c1 & bh7_w70_22_c1 & bh7_w69_21_c1 & bh7_w68_23_c1 & bh7_w67_22_c1 & bh7_w66_24_c1 & bh7_w65_20_c1 & bh7_w64_26_c1 & bh7_w63_25_c1 & bh7_w62_22_c1 & bh7_w61_25_c1 & bh7_w60_24_c1 & bh7_w59_23_c1 & bh7_w58_25_c1 & bh7_w57_25_c1 & bh7_w56_21_c1 & bh7_w55_22_c1 & bh7_w54_22_c1 & bh7_w53_19_c1 & bh7_w52_18_c1 & bh7_w51_15_c1 & bh7_w50_13_c1 & bh7_w49_9_c1 & bh7_w48_11_c1 & bh7_w47_7_c1 & bh7_w46_10_c1 & bh7_w45_7_c1 & bh7_w44_10_c1 & bh7_w43_7_c1 & bh7_w42_10_c1 & bh7_w41_7_c1 & bh7_w40_10_c1 & bh7_w39_7_c1 & bh7_w38_9_c1 & bh7_w37_6_c1 & bh7_w36_9_c1 & bh7_w35_9_c1 & bh7_w34_7_c1 & bh7_w33_7_c1 & bh7_w32_6_c1 & bh7_w31_7_c1 & bh7_w30_6_c1 & bh7_w29_7_c1 & bh7_w28_6_c1 & bh7_w27_7_c1 & bh7_w26_6_c1 & bh7_w25_7_c1 & bh7_w24_6_c1 & bh7_w23_7_c1;
   bitheapFinalAdd_bh7_In1_c1 <= "0" & "0" & bh7_w104_8_c1 & "0" & bh7_w102_14_c1 & "0" & "0" & bh7_w99_18_c1 & "0" & "0" & bh7_w96_20_c1 & "0" & bh7_w94_19_c1 & "0" & bh7_w92_20_c1 & "0" & bh7_w90_22_c1 & "0" & bh7_w88_22_c1 & "0" & "0" & "0" & bh7_w84_22_c1 & "0" & bh7_w82_25_c1 & "0" & bh7_w80_25_c1 & "0" & "0" & bh7_w77_18_c1 & "0" & bh7_w75_19_c1 & "0" & bh7_w73_20_c1 & "0" & "0" & bh7_w70_23_c1 & "0" & bh7_w68_24_c1 & "0" & bh7_w66_25_c1 & "0" & bh7_w64_27_c1 & "0" & bh7_w62_23_c1 & "0" & bh7_w60_25_c1 & "0" & bh7_w58_26_c1 & "0" & bh7_w56_22_c1 & "0" & bh7_w54_21_c1 & "0" & bh7_w52_17_c1 & "0" & bh7_w50_12_c1 & "0" & bh7_w48_10_c1 & "0" & bh7_w46_9_c1 & "0" & bh7_w44_9_c1 & "0" & bh7_w42_9_c1 & "0" & bh7_w40_9_c1 & "0" & "0" & bh7_w37_7_c1 & "0" & bh7_w35_8_c1 & "0" & bh7_w33_6_c1 & "0" & bh7_w31_6_c1 & "0" & bh7_w29_6_c1 & "0" & bh7_w27_6_c1 & "0" & bh7_w25_6_c1 & "0" & bh7_w23_6_c1;
   bitheapFinalAdd_bh7_Cin_c0 <= '0';

   bitheapFinalAdd_bh7: IntAdder_84_Freq300_uid972
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 Cin => bitheapFinalAdd_bh7_Cin_c0,
                 X => bitheapFinalAdd_bh7_In0_c1,
                 Y => bitheapFinalAdd_bh7_In1_c1,
                 R => bitheapFinalAdd_bh7_Out_c2);
   bitheapResult_bh7_c2 <= bitheapFinalAdd_bh7_Out_c2(82 downto 0) & tmp_bitheapResult_bh7_22_c2;
   R <= bitheapResult_bh7_c2(105 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_65_Freq300_uid975
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_65_Freq300_uid975 is
    port (clk, ce_1, ce_2, ce_3 : in std_logic;
          X : in  std_logic_vector(64 downto 0);
          Y : in  std_logic_vector(64 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(64 downto 0)   );
end entity;

architecture arch of IntAdder_65_Freq300_uid975 is
signal Cin_1_c2, Cin_1_c3 :  std_logic;
signal X_1_c2, X_1_c3 :  std_logic_vector(65 downto 0);
signal Y_1_c0, Y_1_c1, Y_1_c2, Y_1_c3 :  std_logic_vector(65 downto 0);
signal S_1_c3 :  std_logic_vector(65 downto 0);
signal R_1_c3 :  std_logic_vector(64 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               Y_1_c1 <= Y_1_c0;
            end if;
            if ce_2 = '1' then
               Y_1_c2 <= Y_1_c1;
            end if;
            if ce_3 = '1' then
               Cin_1_c3 <= Cin_1_c2;
               X_1_c3 <= X_1_c2;
               Y_1_c3 <= Y_1_c2;
            end if;
         end if;
      end process;
   Cin_1_c2 <= Cin;
   X_1_c2 <= '0' & X(64 downto 0);
   Y_1_c0 <= '0' & Y(64 downto 0);
   S_1_c3 <= X_1_c3 + Y_1_c3 + Cin_1_c3;
   R_1_c3 <= S_1_c3(64 downto 0);
   R <= R_1_c3 ;
end architecture;

--------------------------------------------------------------------------------
--                          FloatingPointMultiplier
--                      (FPMult_11_52_uid2_Freq300_uid3)
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin 2008-2021
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointMultiplier_64_4_242333 is
    port (clk, ce_1, ce_2, ce_3 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointMultiplier_64_4_242333 is
   component IntMultiplier_53x53_106_Freq300_uid5 is
      port ( clk, ce_1, ce_2 : in std_logic;
             X : in  std_logic_vector(52 downto 0);
             Y : in  std_logic_vector(52 downto 0);
             R : out  std_logic_vector(105 downto 0)   );
   end component;

   component IntAdder_65_Freq300_uid975 is
      port ( clk, ce_1, ce_2, ce_3 : in std_logic;
             X : in  std_logic_vector(64 downto 0);
             Y : in  std_logic_vector(64 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(64 downto 0)   );
   end component;

signal sign_c0, sign_c1, sign_c2, sign_c3 :  std_logic;
signal expX_c0 :  std_logic_vector(10 downto 0);
signal expY_c0 :  std_logic_vector(10 downto 0);
signal expSumPreSub_c0 :  std_logic_vector(12 downto 0);
signal bias_c0 :  std_logic_vector(12 downto 0);
signal expSum_c0, expSum_c1, expSum_c2 :  std_logic_vector(12 downto 0);
signal sigX_c0 :  std_logic_vector(52 downto 0);
signal sigY_c0 :  std_logic_vector(52 downto 0);
signal sigProd_c2 :  std_logic_vector(105 downto 0);
signal excSel_c0 :  std_logic_vector(3 downto 0);
signal exc_c0, exc_c1, exc_c2, exc_c3 :  std_logic_vector(1 downto 0);
signal norm_c2 :  std_logic;
signal expPostNorm_c2 :  std_logic_vector(12 downto 0);
signal sigProdExt_c2 :  std_logic_vector(105 downto 0);
signal expSig_c2 :  std_logic_vector(64 downto 0);
signal sticky_c2 :  std_logic;
signal guard_c2 :  std_logic;
signal round_c2 :  std_logic;
signal expSigPostRound_c3 :  std_logic_vector(64 downto 0);
signal excPostNorm_c3 :  std_logic_vector(1 downto 0);
signal finalExc_c3 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               sign_c1 <= sign_c0;
               expSum_c1 <= expSum_c0;
               exc_c1 <= exc_c0;
            end if;
            if ce_2 = '1' then
               sign_c2 <= sign_c1;
               expSum_c2 <= expSum_c1;
               exc_c2 <= exc_c1;
            end if;
            if ce_3 = '1' then
               sign_c3 <= sign_c2;
               exc_c3 <= exc_c2;
            end if;
         end if;
      end process;
   sign_c0 <= X(63) xor Y(63);
   expX_c0 <= X(62 downto 52);
   expY_c0 <= Y(62 downto 52);
   expSumPreSub_c0 <= ("00" & expX_c0) + ("00" & expY_c0);
   bias_c0 <= CONV_STD_LOGIC_VECTOR(1023,13);
   expSum_c0 <= expSumPreSub_c0 - bias_c0;
   sigX_c0 <= "1" & X(51 downto 0);
   sigY_c0 <= "1" & Y(51 downto 0);
   SignificandMultiplication: IntMultiplier_53x53_106_Freq300_uid5
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 X => sigX_c0,
                 Y => sigY_c0,
                 R => sigProd_c2);
   excSel_c0 <= X(65 downto 64) & Y(65 downto 64);
   with excSel_c0  select  
   exc_c0 <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;
   norm_c2 <= sigProd_c2(105);
   -- exponent update
   expPostNorm_c2 <= expSum_c2 + ("000000000000" & norm_c2);
   -- significand normalization shift
   sigProdExt_c2 <= sigProd_c2(104 downto 0) & "0" when norm_c2='1' else
                         sigProd_c2(103 downto 0) & "00";
   expSig_c2 <= expPostNorm_c2 & sigProdExt_c2(105 downto 54);
   sticky_c2 <= sigProdExt_c2(53);
   guard_c2 <= '0' when sigProdExt_c2(52 downto 0)="00000000000000000000000000000000000000000000000000000" else '1';
   round_c2 <= sticky_c2 and ( (guard_c2 and not(sigProdExt_c2(54))) or (sigProdExt_c2(54) ))  ;
   RoundingAdder: IntAdder_65_Freq300_uid975
      port map ( clk  => clk,
                 ce_1 => ce_1,
                 ce_2=> ce_2,
                 ce_3=> ce_3,
                 Cin => round_c2,
                 X => expSig_c2,
                 Y => "00000000000000000000000000000000000000000000000000000000000000000",
                 R => expSigPostRound_c3);
   with expSigPostRound_c3(64 downto 63)  select 
   excPostNorm_c3 <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc_c3  select  
   finalExc_c3 <= exc_c3 when  "11"|"10"|"00",
                       excPostNorm_c3 when others; 
   R <= finalExc_c3 & sign_c3 & expSigPostRound_c3(62 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          selFunction_Freq800_uid4
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity selFunction_Freq800_uid4 is
    port (X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of selFunction_Freq800_uid4 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000000000",
      "000" when "000000001",
      "000" when "000000010",
      "000" when "000000011",
      "000" when "000000100",
      "000" when "000000101",
      "000" when "000000110",
      "000" when "000000111",
      "000" when "000001000",
      "000" when "000001001",
      "000" when "000001010",
      "000" when "000001011",
      "000" when "000001100",
      "000" when "000001101",
      "000" when "000001110",
      "000" when "000001111",
      "001" when "000010000",
      "000" when "000010001",
      "000" when "000010010",
      "000" when "000010011",
      "000" when "000010100",
      "000" when "000010101",
      "000" when "000010110",
      "000" when "000010111",
      "001" when "000011000",
      "001" when "000011001",
      "001" when "000011010",
      "001" when "000011011",
      "000" when "000011100",
      "000" when "000011101",
      "000" when "000011110",
      "000" when "000011111",
      "001" when "000100000",
      "001" when "000100001",
      "001" when "000100010",
      "001" when "000100011",
      "001" when "000100100",
      "001" when "000100101",
      "001" when "000100110",
      "000" when "000100111",
      "001" when "000101000",
      "001" when "000101001",
      "001" when "000101010",
      "001" when "000101011",
      "001" when "000101100",
      "001" when "000101101",
      "001" when "000101110",
      "001" when "000101111",
      "010" when "000110000",
      "001" when "000110001",
      "001" when "000110010",
      "001" when "000110011",
      "001" when "000110100",
      "001" when "000110101",
      "001" when "000110110",
      "001" when "000110111",
      "010" when "000111000",
      "010" when "000111001",
      "001" when "000111010",
      "001" when "000111011",
      "001" when "000111100",
      "001" when "000111101",
      "001" when "000111110",
      "001" when "000111111",
      "010" when "001000000",
      "010" when "001000001",
      "010" when "001000010",
      "001" when "001000011",
      "001" when "001000100",
      "001" when "001000101",
      "001" when "001000110",
      "001" when "001000111",
      "010" when "001001000",
      "010" when "001001001",
      "010" when "001001010",
      "010" when "001001011",
      "001" when "001001100",
      "001" when "001001101",
      "001" when "001001110",
      "001" when "001001111",
      "010" when "001010000",
      "010" when "001010001",
      "010" when "001010010",
      "010" when "001010011",
      "010" when "001010100",
      "010" when "001010101",
      "001" when "001010110",
      "001" when "001010111",
      "010" when "001011000",
      "010" when "001011001",
      "010" when "001011010",
      "010" when "001011011",
      "010" when "001011100",
      "010" when "001011101",
      "010" when "001011110",
      "001" when "001011111",
      "010" when "001100000",
      "010" when "001100001",
      "010" when "001100010",
      "010" when "001100011",
      "010" when "001100100",
      "010" when "001100101",
      "010" when "001100110",
      "010" when "001100111",
      "010" when "001101000",
      "010" when "001101001",
      "010" when "001101010",
      "010" when "001101011",
      "010" when "001101100",
      "010" when "001101101",
      "010" when "001101110",
      "010" when "001101111",
      "010" when "001110000",
      "010" when "001110001",
      "010" when "001110010",
      "010" when "001110011",
      "010" when "001110100",
      "010" when "001110101",
      "010" when "001110110",
      "010" when "001110111",
      "010" when "001111000",
      "010" when "001111001",
      "010" when "001111010",
      "010" when "001111011",
      "010" when "001111100",
      "010" when "001111101",
      "010" when "001111110",
      "010" when "001111111",
      "010" when "010000000",
      "010" when "010000001",
      "010" when "010000010",
      "010" when "010000011",
      "010" when "010000100",
      "010" when "010000101",
      "010" when "010000110",
      "010" when "010000111",
      "010" when "010001000",
      "010" when "010001001",
      "010" when "010001010",
      "010" when "010001011",
      "010" when "010001100",
      "010" when "010001101",
      "010" when "010001110",
      "010" when "010001111",
      "010" when "010010000",
      "010" when "010010001",
      "010" when "010010010",
      "010" when "010010011",
      "010" when "010010100",
      "010" when "010010101",
      "010" when "010010110",
      "010" when "010010111",
      "010" when "010011000",
      "010" when "010011001",
      "010" when "010011010",
      "010" when "010011011",
      "010" when "010011100",
      "010" when "010011101",
      "010" when "010011110",
      "010" when "010011111",
      "010" when "010100000",
      "010" when "010100001",
      "010" when "010100010",
      "010" when "010100011",
      "010" when "010100100",
      "010" when "010100101",
      "010" when "010100110",
      "010" when "010100111",
      "010" when "010101000",
      "010" when "010101001",
      "010" when "010101010",
      "010" when "010101011",
      "010" when "010101100",
      "010" when "010101101",
      "010" when "010101110",
      "010" when "010101111",
      "010" when "010110000",
      "010" when "010110001",
      "010" when "010110010",
      "010" when "010110011",
      "010" when "010110100",
      "010" when "010110101",
      "010" when "010110110",
      "010" when "010110111",
      "010" when "010111000",
      "010" when "010111001",
      "010" when "010111010",
      "010" when "010111011",
      "010" when "010111100",
      "010" when "010111101",
      "010" when "010111110",
      "010" when "010111111",
      "010" when "011000000",
      "010" when "011000001",
      "010" when "011000010",
      "010" when "011000011",
      "010" when "011000100",
      "010" when "011000101",
      "010" when "011000110",
      "010" when "011000111",
      "010" when "011001000",
      "010" when "011001001",
      "010" when "011001010",
      "010" when "011001011",
      "010" when "011001100",
      "010" when "011001101",
      "010" when "011001110",
      "010" when "011001111",
      "010" when "011010000",
      "010" when "011010001",
      "010" when "011010010",
      "010" when "011010011",
      "010" when "011010100",
      "010" when "011010101",
      "010" when "011010110",
      "010" when "011010111",
      "010" when "011011000",
      "010" when "011011001",
      "010" when "011011010",
      "010" when "011011011",
      "010" when "011011100",
      "010" when "011011101",
      "010" when "011011110",
      "010" when "011011111",
      "010" when "011100000",
      "010" when "011100001",
      "010" when "011100010",
      "010" when "011100011",
      "010" when "011100100",
      "010" when "011100101",
      "010" when "011100110",
      "010" when "011100111",
      "010" when "011101000",
      "010" when "011101001",
      "010" when "011101010",
      "010" when "011101011",
      "010" when "011101100",
      "010" when "011101101",
      "010" when "011101110",
      "010" when "011101111",
      "010" when "011110000",
      "010" when "011110001",
      "010" when "011110010",
      "010" when "011110011",
      "010" when "011110100",
      "010" when "011110101",
      "010" when "011110110",
      "010" when "011110111",
      "010" when "011111000",
      "010" when "011111001",
      "010" when "011111010",
      "010" when "011111011",
      "010" when "011111100",
      "010" when "011111101",
      "010" when "011111110",
      "010" when "011111111",
      "110" when "100000000",
      "110" when "100000001",
      "110" when "100000010",
      "110" when "100000011",
      "110" when "100000100",
      "110" when "100000101",
      "110" when "100000110",
      "110" when "100000111",
      "110" when "100001000",
      "110" when "100001001",
      "110" when "100001010",
      "110" when "100001011",
      "110" when "100001100",
      "110" when "100001101",
      "110" when "100001110",
      "110" when "100001111",
      "110" when "100010000",
      "110" when "100010001",
      "110" when "100010010",
      "110" when "100010011",
      "110" when "100010100",
      "110" when "100010101",
      "110" when "100010110",
      "110" when "100010111",
      "110" when "100011000",
      "110" when "100011001",
      "110" when "100011010",
      "110" when "100011011",
      "110" when "100011100",
      "110" when "100011101",
      "110" when "100011110",
      "110" when "100011111",
      "110" when "100100000",
      "110" when "100100001",
      "110" when "100100010",
      "110" when "100100011",
      "110" when "100100100",
      "110" when "100100101",
      "110" when "100100110",
      "110" when "100100111",
      "110" when "100101000",
      "110" when "100101001",
      "110" when "100101010",
      "110" when "100101011",
      "110" when "100101100",
      "110" when "100101101",
      "110" when "100101110",
      "110" when "100101111",
      "110" when "100110000",
      "110" when "100110001",
      "110" when "100110010",
      "110" when "100110011",
      "110" when "100110100",
      "110" when "100110101",
      "110" when "100110110",
      "110" when "100110111",
      "110" when "100111000",
      "110" when "100111001",
      "110" when "100111010",
      "110" when "100111011",
      "110" when "100111100",
      "110" when "100111101",
      "110" when "100111110",
      "110" when "100111111",
      "110" when "101000000",
      "110" when "101000001",
      "110" when "101000010",
      "110" when "101000011",
      "110" when "101000100",
      "110" when "101000101",
      "110" when "101000110",
      "110" when "101000111",
      "110" when "101001000",
      "110" when "101001001",
      "110" when "101001010",
      "110" when "101001011",
      "110" when "101001100",
      "110" when "101001101",
      "110" when "101001110",
      "110" when "101001111",
      "110" when "101010000",
      "110" when "101010001",
      "110" when "101010010",
      "110" when "101010011",
      "110" when "101010100",
      "110" when "101010101",
      "110" when "101010110",
      "110" when "101010111",
      "110" when "101011000",
      "110" when "101011001",
      "110" when "101011010",
      "110" when "101011011",
      "110" when "101011100",
      "110" when "101011101",
      "110" when "101011110",
      "110" when "101011111",
      "110" when "101100000",
      "110" when "101100001",
      "110" when "101100010",
      "110" when "101100011",
      "110" when "101100100",
      "110" when "101100101",
      "110" when "101100110",
      "110" when "101100111",
      "110" when "101101000",
      "110" when "101101001",
      "110" when "101101010",
      "110" when "101101011",
      "110" when "101101100",
      "110" when "101101101",
      "110" when "101101110",
      "110" when "101101111",
      "110" when "101110000",
      "110" when "101110001",
      "110" when "101110010",
      "110" when "101110011",
      "110" when "101110100",
      "110" when "101110101",
      "110" when "101110110",
      "110" when "101110111",
      "110" when "101111000",
      "110" when "101111001",
      "110" when "101111010",
      "110" when "101111011",
      "110" when "101111100",
      "110" when "101111101",
      "110" when "101111110",
      "110" when "101111111",
      "110" when "110000000",
      "110" when "110000001",
      "110" when "110000010",
      "110" when "110000011",
      "110" when "110000100",
      "110" when "110000101",
      "110" when "110000110",
      "110" when "110000111",
      "110" when "110001000",
      "110" when "110001001",
      "110" when "110001010",
      "110" when "110001011",
      "110" when "110001100",
      "110" when "110001101",
      "110" when "110001110",
      "110" when "110001111",
      "110" when "110010000",
      "110" when "110010001",
      "110" when "110010010",
      "110" when "110010011",
      "110" when "110010100",
      "110" when "110010101",
      "110" when "110010110",
      "110" when "110010111",
      "110" when "110011000",
      "110" when "110011001",
      "110" when "110011010",
      "110" when "110011011",
      "110" when "110011100",
      "110" when "110011101",
      "110" when "110011110",
      "110" when "110011111",
      "110" when "110100000",
      "110" when "110100001",
      "110" when "110100010",
      "110" when "110100011",
      "110" when "110100100",
      "110" when "110100101",
      "110" when "110100110",
      "110" when "110100111",
      "110" when "110101000",
      "110" when "110101001",
      "110" when "110101010",
      "110" when "110101011",
      "110" when "110101100",
      "110" when "110101101",
      "110" when "110101110",
      "111" when "110101111",
      "110" when "110110000",
      "110" when "110110001",
      "110" when "110110010",
      "110" when "110110011",
      "110" when "110110100",
      "111" when "110110101",
      "111" when "110110110",
      "111" when "110110111",
      "110" when "110111000",
      "110" when "110111001",
      "110" when "110111010",
      "110" when "110111011",
      "111" when "110111100",
      "111" when "110111101",
      "111" when "110111110",
      "111" when "110111111",
      "110" when "111000000",
      "110" when "111000001",
      "111" when "111000010",
      "111" when "111000011",
      "111" when "111000100",
      "111" when "111000101",
      "111" when "111000110",
      "111" when "111000111",
      "110" when "111001000",
      "111" when "111001001",
      "111" when "111001010",
      "111" when "111001011",
      "111" when "111001100",
      "111" when "111001101",
      "111" when "111001110",
      "111" when "111001111",
      "111" when "111010000",
      "111" when "111010001",
      "111" when "111010010",
      "111" when "111010011",
      "111" when "111010100",
      "111" when "111010101",
      "111" when "111010110",
      "111" when "111010111",
      "111" when "111011000",
      "111" when "111011001",
      "111" when "111011010",
      "111" when "111011011",
      "111" when "111011100",
      "111" when "111011101",
      "111" when "111011110",
      "111" when "111011111",
      "111" when "111100000",
      "111" when "111100001",
      "111" when "111100010",
      "111" when "111100011",
      "111" when "111100100",
      "111" when "111100101",
      "111" when "111100110",
      "111" when "111100111",
      "111" when "111101000",
      "111" when "111101001",
      "111" when "111101010",
      "111" when "111101011",
      "000" when "111101100",
      "000" when "111101101",
      "000" when "111101110",
      "000" when "111101111",
      "000" when "111110000",
      "000" when "111110001",
      "000" when "111110010",
      "000" when "111110011",
      "000" when "111110100",
      "000" when "111110101",
      "000" when "111110110",
      "000" when "111110111",
      "000" when "111111000",
      "000" when "111111001",
      "000" when "111111010",
      "000" when "111111011",
      "000" when "111111100",
      "000" when "111111101",
      "000" when "111111110",
      "000" when "111111111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            FloatingPointDivider
--                         (FPDiv_11_52_Freq800_uid2)
-- VHDL generated for Kintex7 @ 800MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 63 cycles
-- Clock period (ns): 1.25
-- Target frequency (MHz): 800
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointDivider_64_4_345000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36, ce_37, ce_38, ce_39, ce_40, ce_41, ce_42, ce_43, ce_44, ce_45, ce_46, ce_47, ce_48, ce_49, ce_50, ce_51, ce_52, ce_53, ce_54, ce_55, ce_56, ce_57, ce_58, ce_59, ce_60, ce_61, ce_62, ce_63 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointDivider_64_4_345000 is
   component selFunction_Freq800_uid4 is
      port ( X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal fX_c0 :  std_logic_vector(52 downto 0);
signal fY_c0 :  std_logic_vector(52 downto 0);
signal expR0_c0, expR0_c1, expR0_c2, expR0_c3, expR0_c4, expR0_c5, expR0_c6, expR0_c7, expR0_c8, expR0_c9, expR0_c10, expR0_c11, expR0_c12, expR0_c13, expR0_c14, expR0_c15, expR0_c16, expR0_c17, expR0_c18, expR0_c19, expR0_c20, expR0_c21, expR0_c22, expR0_c23, expR0_c24, expR0_c25, expR0_c26, expR0_c27, expR0_c28, expR0_c29, expR0_c30, expR0_c31, expR0_c32, expR0_c33, expR0_c34, expR0_c35, expR0_c36, expR0_c37, expR0_c38, expR0_c39, expR0_c40, expR0_c41, expR0_c42, expR0_c43, expR0_c44, expR0_c45, expR0_c46, expR0_c47, expR0_c48, expR0_c49, expR0_c50, expR0_c51, expR0_c52, expR0_c53, expR0_c54, expR0_c55, expR0_c56, expR0_c57, expR0_c58, expR0_c59, expR0_c60, expR0_c61, expR0_c62 :  std_logic_vector(12 downto 0);
signal sR_c0, sR_c1, sR_c2, sR_c3, sR_c4, sR_c5, sR_c6, sR_c7, sR_c8, sR_c9, sR_c10, sR_c11, sR_c12, sR_c13, sR_c14, sR_c15, sR_c16, sR_c17, sR_c18, sR_c19, sR_c20, sR_c21, sR_c22, sR_c23, sR_c24, sR_c25, sR_c26, sR_c27, sR_c28, sR_c29, sR_c30, sR_c31, sR_c32, sR_c33, sR_c34, sR_c35, sR_c36, sR_c37, sR_c38, sR_c39, sR_c40, sR_c41, sR_c42, sR_c43, sR_c44, sR_c45, sR_c46, sR_c47, sR_c48, sR_c49, sR_c50, sR_c51, sR_c52, sR_c53, sR_c54, sR_c55, sR_c56, sR_c57, sR_c58, sR_c59, sR_c60, sR_c61, sR_c62, sR_c63 :  std_logic;
signal exnXY_c0 :  std_logic_vector(3 downto 0);
signal exnR0_c0, exnR0_c1, exnR0_c2, exnR0_c3, exnR0_c4, exnR0_c5, exnR0_c6, exnR0_c7, exnR0_c8, exnR0_c9, exnR0_c10, exnR0_c11, exnR0_c12, exnR0_c13, exnR0_c14, exnR0_c15, exnR0_c16, exnR0_c17, exnR0_c18, exnR0_c19, exnR0_c20, exnR0_c21, exnR0_c22, exnR0_c23, exnR0_c24, exnR0_c25, exnR0_c26, exnR0_c27, exnR0_c28, exnR0_c29, exnR0_c30, exnR0_c31, exnR0_c32, exnR0_c33, exnR0_c34, exnR0_c35, exnR0_c36, exnR0_c37, exnR0_c38, exnR0_c39, exnR0_c40, exnR0_c41, exnR0_c42, exnR0_c43, exnR0_c44, exnR0_c45, exnR0_c46, exnR0_c47, exnR0_c48, exnR0_c49, exnR0_c50, exnR0_c51, exnR0_c52, exnR0_c53, exnR0_c54, exnR0_c55, exnR0_c56, exnR0_c57, exnR0_c58, exnR0_c59, exnR0_c60, exnR0_c61, exnR0_c62, exnR0_c63 :  std_logic_vector(1 downto 0);
signal D_c0, D_c1, D_c2, D_c3, D_c4, D_c5, D_c6, D_c7, D_c8, D_c9, D_c10, D_c11, D_c12, D_c13, D_c14, D_c15, D_c16, D_c17, D_c18, D_c19, D_c20, D_c21, D_c22, D_c23, D_c24, D_c25, D_c26, D_c27, D_c28, D_c29, D_c30, D_c31, D_c32, D_c33, D_c34, D_c35, D_c36, D_c37, D_c38, D_c39, D_c40, D_c41, D_c42, D_c43, D_c44, D_c45, D_c46, D_c47, D_c48, D_c49, D_c50, D_c51, D_c52, D_c53, D_c54, D_c55, D_c56, D_c57, D_c58 :  std_logic_vector(52 downto 0);
signal psX_c0 :  std_logic_vector(53 downto 0);
signal betaw28_c0, betaw28_c1, betaw28_c2 :  std_logic_vector(55 downto 0);
signal sel28_c0 :  std_logic_vector(8 downto 0);
signal q28_c0, q28_c1, q28_c2 :  std_logic_vector(2 downto 0);
signal q28_copy5_c0 :  std_logic_vector(2 downto 0);
signal absq28D_c0, absq28D_c1, absq28D_c2 :  std_logic_vector(55 downto 0);
signal w27_c2 :  std_logic_vector(55 downto 0);
signal betaw27_c2, betaw27_c3, betaw27_c4 :  std_logic_vector(55 downto 0);
signal sel27_c2 :  std_logic_vector(8 downto 0);
signal q27_c2, q27_c3, q27_c4 :  std_logic_vector(2 downto 0);
signal q27_copy6_c2 :  std_logic_vector(2 downto 0);
signal absq27D_c2, absq27D_c3, absq27D_c4 :  std_logic_vector(55 downto 0);
signal w26_c4 :  std_logic_vector(55 downto 0);
signal betaw26_c4, betaw26_c5, betaw26_c6 :  std_logic_vector(55 downto 0);
signal sel26_c4 :  std_logic_vector(8 downto 0);
signal q26_c4, q26_c5, q26_c6 :  std_logic_vector(2 downto 0);
signal q26_copy7_c4 :  std_logic_vector(2 downto 0);
signal absq26D_c4, absq26D_c5, absq26D_c6 :  std_logic_vector(55 downto 0);
signal w25_c6 :  std_logic_vector(55 downto 0);
signal betaw25_c6, betaw25_c7, betaw25_c8 :  std_logic_vector(55 downto 0);
signal sel25_c6 :  std_logic_vector(8 downto 0);
signal q25_c6, q25_c7, q25_c8 :  std_logic_vector(2 downto 0);
signal q25_copy8_c6 :  std_logic_vector(2 downto 0);
signal absq25D_c6, absq25D_c7, absq25D_c8 :  std_logic_vector(55 downto 0);
signal w24_c8 :  std_logic_vector(55 downto 0);
signal betaw24_c8, betaw24_c9, betaw24_c10 :  std_logic_vector(55 downto 0);
signal sel24_c8 :  std_logic_vector(8 downto 0);
signal q24_c9, q24_c10 :  std_logic_vector(2 downto 0);
signal q24_copy9_c8, q24_copy9_c9 :  std_logic_vector(2 downto 0);
signal absq24D_c9, absq24D_c10 :  std_logic_vector(55 downto 0);
signal w23_c10 :  std_logic_vector(55 downto 0);
signal betaw23_c10, betaw23_c11, betaw23_c12 :  std_logic_vector(55 downto 0);
signal sel23_c10 :  std_logic_vector(8 downto 0);
signal q23_c11, q23_c12 :  std_logic_vector(2 downto 0);
signal q23_copy10_c10, q23_copy10_c11 :  std_logic_vector(2 downto 0);
signal absq23D_c11, absq23D_c12 :  std_logic_vector(55 downto 0);
signal w22_c12 :  std_logic_vector(55 downto 0);
signal betaw22_c12, betaw22_c13, betaw22_c14, betaw22_c15 :  std_logic_vector(55 downto 0);
signal sel22_c12 :  std_logic_vector(8 downto 0);
signal q22_c13, q22_c14, q22_c15 :  std_logic_vector(2 downto 0);
signal q22_copy11_c12, q22_copy11_c13 :  std_logic_vector(2 downto 0);
signal absq22D_c13, absq22D_c14, absq22D_c15 :  std_logic_vector(55 downto 0);
signal w21_c15 :  std_logic_vector(55 downto 0);
signal betaw21_c15, betaw21_c16, betaw21_c17 :  std_logic_vector(55 downto 0);
signal sel21_c15 :  std_logic_vector(8 downto 0);
signal q21_c15, q21_c16, q21_c17 :  std_logic_vector(2 downto 0);
signal q21_copy12_c15 :  std_logic_vector(2 downto 0);
signal absq21D_c15, absq21D_c16, absq21D_c17 :  std_logic_vector(55 downto 0);
signal w20_c17 :  std_logic_vector(55 downto 0);
signal betaw20_c17, betaw20_c18, betaw20_c19 :  std_logic_vector(55 downto 0);
signal sel20_c17 :  std_logic_vector(8 downto 0);
signal q20_c17, q20_c18, q20_c19 :  std_logic_vector(2 downto 0);
signal q20_copy13_c17 :  std_logic_vector(2 downto 0);
signal absq20D_c17, absq20D_c18, absq20D_c19 :  std_logic_vector(55 downto 0);
signal w19_c19 :  std_logic_vector(55 downto 0);
signal betaw19_c19, betaw19_c20, betaw19_c21 :  std_logic_vector(55 downto 0);
signal sel19_c19 :  std_logic_vector(8 downto 0);
signal q19_c19, q19_c20, q19_c21 :  std_logic_vector(2 downto 0);
signal q19_copy14_c19 :  std_logic_vector(2 downto 0);
signal absq19D_c19, absq19D_c20, absq19D_c21 :  std_logic_vector(55 downto 0);
signal w18_c21 :  std_logic_vector(55 downto 0);
signal betaw18_c21, betaw18_c22, betaw18_c23 :  std_logic_vector(55 downto 0);
signal sel18_c21 :  std_logic_vector(8 downto 0);
signal q18_c22, q18_c23 :  std_logic_vector(2 downto 0);
signal q18_copy15_c21, q18_copy15_c22 :  std_logic_vector(2 downto 0);
signal absq18D_c22, absq18D_c23 :  std_logic_vector(55 downto 0);
signal w17_c23 :  std_logic_vector(55 downto 0);
signal betaw17_c23, betaw17_c24, betaw17_c25 :  std_logic_vector(55 downto 0);
signal sel17_c23 :  std_logic_vector(8 downto 0);
signal q17_c24, q17_c25 :  std_logic_vector(2 downto 0);
signal q17_copy16_c23, q17_copy16_c24 :  std_logic_vector(2 downto 0);
signal absq17D_c24, absq17D_c25 :  std_logic_vector(55 downto 0);
signal w16_c25 :  std_logic_vector(55 downto 0);
signal betaw16_c25, betaw16_c26, betaw16_c27 :  std_logic_vector(55 downto 0);
signal sel16_c25 :  std_logic_vector(8 downto 0);
signal q16_c26, q16_c27 :  std_logic_vector(2 downto 0);
signal q16_copy17_c25, q16_copy17_c26 :  std_logic_vector(2 downto 0);
signal absq16D_c26, absq16D_c27 :  std_logic_vector(55 downto 0);
signal w15_c27 :  std_logic_vector(55 downto 0);
signal betaw15_c27, betaw15_c28, betaw15_c29, betaw15_c30 :  std_logic_vector(55 downto 0);
signal sel15_c27 :  std_logic_vector(8 downto 0);
signal q15_c28, q15_c29, q15_c30 :  std_logic_vector(2 downto 0);
signal q15_copy18_c27, q15_copy18_c28 :  std_logic_vector(2 downto 0);
signal absq15D_c28, absq15D_c29, absq15D_c30 :  std_logic_vector(55 downto 0);
signal w14_c30 :  std_logic_vector(55 downto 0);
signal betaw14_c30, betaw14_c31, betaw14_c32 :  std_logic_vector(55 downto 0);
signal sel14_c30 :  std_logic_vector(8 downto 0);
signal q14_c30, q14_c31, q14_c32 :  std_logic_vector(2 downto 0);
signal q14_copy19_c30 :  std_logic_vector(2 downto 0);
signal absq14D_c30, absq14D_c31, absq14D_c32 :  std_logic_vector(55 downto 0);
signal w13_c32 :  std_logic_vector(55 downto 0);
signal betaw13_c32, betaw13_c33, betaw13_c34 :  std_logic_vector(55 downto 0);
signal sel13_c32 :  std_logic_vector(8 downto 0);
signal q13_c32, q13_c33, q13_c34 :  std_logic_vector(2 downto 0);
signal q13_copy20_c32 :  std_logic_vector(2 downto 0);
signal absq13D_c32, absq13D_c33, absq13D_c34 :  std_logic_vector(55 downto 0);
signal w12_c34 :  std_logic_vector(55 downto 0);
signal betaw12_c34, betaw12_c35, betaw12_c36 :  std_logic_vector(55 downto 0);
signal sel12_c34 :  std_logic_vector(8 downto 0);
signal q12_c34, q12_c35, q12_c36 :  std_logic_vector(2 downto 0);
signal q12_copy21_c34 :  std_logic_vector(2 downto 0);
signal absq12D_c34, absq12D_c35, absq12D_c36 :  std_logic_vector(55 downto 0);
signal w11_c36 :  std_logic_vector(55 downto 0);
signal betaw11_c36, betaw11_c37, betaw11_c38 :  std_logic_vector(55 downto 0);
signal sel11_c36 :  std_logic_vector(8 downto 0);
signal q11_c37, q11_c38 :  std_logic_vector(2 downto 0);
signal q11_copy22_c36, q11_copy22_c37 :  std_logic_vector(2 downto 0);
signal absq11D_c37, absq11D_c38 :  std_logic_vector(55 downto 0);
signal w10_c38 :  std_logic_vector(55 downto 0);
signal betaw10_c38, betaw10_c39, betaw10_c40 :  std_logic_vector(55 downto 0);
signal sel10_c38 :  std_logic_vector(8 downto 0);
signal q10_c39, q10_c40 :  std_logic_vector(2 downto 0);
signal q10_copy23_c38, q10_copy23_c39 :  std_logic_vector(2 downto 0);
signal absq10D_c39, absq10D_c40 :  std_logic_vector(55 downto 0);
signal w9_c40 :  std_logic_vector(55 downto 0);
signal betaw9_c40, betaw9_c41, betaw9_c42 :  std_logic_vector(55 downto 0);
signal sel9_c40 :  std_logic_vector(8 downto 0);
signal q9_c41, q9_c42 :  std_logic_vector(2 downto 0);
signal q9_copy24_c40, q9_copy24_c41 :  std_logic_vector(2 downto 0);
signal absq9D_c41, absq9D_c42 :  std_logic_vector(55 downto 0);
signal w8_c42 :  std_logic_vector(55 downto 0);
signal betaw8_c42, betaw8_c43, betaw8_c44, betaw8_c45 :  std_logic_vector(55 downto 0);
signal sel8_c42 :  std_logic_vector(8 downto 0);
signal q8_c43, q8_c44, q8_c45 :  std_logic_vector(2 downto 0);
signal q8_copy25_c42, q8_copy25_c43 :  std_logic_vector(2 downto 0);
signal absq8D_c43, absq8D_c44, absq8D_c45 :  std_logic_vector(55 downto 0);
signal w7_c45 :  std_logic_vector(55 downto 0);
signal betaw7_c45, betaw7_c46, betaw7_c47 :  std_logic_vector(55 downto 0);
signal sel7_c45 :  std_logic_vector(8 downto 0);
signal q7_c45, q7_c46, q7_c47 :  std_logic_vector(2 downto 0);
signal q7_copy26_c45 :  std_logic_vector(2 downto 0);
signal absq7D_c45, absq7D_c46, absq7D_c47 :  std_logic_vector(55 downto 0);
signal w6_c47 :  std_logic_vector(55 downto 0);
signal betaw6_c47, betaw6_c48, betaw6_c49 :  std_logic_vector(55 downto 0);
signal sel6_c47 :  std_logic_vector(8 downto 0);
signal q6_c47, q6_c48, q6_c49 :  std_logic_vector(2 downto 0);
signal q6_copy27_c47 :  std_logic_vector(2 downto 0);
signal absq6D_c47, absq6D_c48, absq6D_c49 :  std_logic_vector(55 downto 0);
signal w5_c49 :  std_logic_vector(55 downto 0);
signal betaw5_c49, betaw5_c50, betaw5_c51 :  std_logic_vector(55 downto 0);
signal sel5_c49 :  std_logic_vector(8 downto 0);
signal q5_c49, q5_c50, q5_c51 :  std_logic_vector(2 downto 0);
signal q5_copy28_c49 :  std_logic_vector(2 downto 0);
signal absq5D_c49, absq5D_c50, absq5D_c51 :  std_logic_vector(55 downto 0);
signal w4_c51 :  std_logic_vector(55 downto 0);
signal betaw4_c51, betaw4_c52, betaw4_c53 :  std_logic_vector(55 downto 0);
signal sel4_c51 :  std_logic_vector(8 downto 0);
signal q4_c52, q4_c53 :  std_logic_vector(2 downto 0);
signal q4_copy29_c51, q4_copy29_c52 :  std_logic_vector(2 downto 0);
signal absq4D_c52, absq4D_c53 :  std_logic_vector(55 downto 0);
signal w3_c53 :  std_logic_vector(55 downto 0);
signal betaw3_c53, betaw3_c54, betaw3_c55 :  std_logic_vector(55 downto 0);
signal sel3_c53 :  std_logic_vector(8 downto 0);
signal q3_c54, q3_c55 :  std_logic_vector(2 downto 0);
signal q3_copy30_c53, q3_copy30_c54 :  std_logic_vector(2 downto 0);
signal absq3D_c54, absq3D_c55 :  std_logic_vector(55 downto 0);
signal w2_c55 :  std_logic_vector(55 downto 0);
signal betaw2_c55, betaw2_c56, betaw2_c57, betaw2_c58 :  std_logic_vector(55 downto 0);
signal sel2_c55 :  std_logic_vector(8 downto 0);
signal q2_c56, q2_c57, q2_c58 :  std_logic_vector(2 downto 0);
signal q2_copy31_c55, q2_copy31_c56 :  std_logic_vector(2 downto 0);
signal absq2D_c56, absq2D_c57, absq2D_c58 :  std_logic_vector(55 downto 0);
signal w1_c58 :  std_logic_vector(55 downto 0);
signal betaw1_c58, betaw1_c59, betaw1_c60 :  std_logic_vector(55 downto 0);
signal sel1_c58 :  std_logic_vector(8 downto 0);
signal q1_c58, q1_c59, q1_c60 :  std_logic_vector(2 downto 0);
signal q1_copy32_c58 :  std_logic_vector(2 downto 0);
signal absq1D_c58, absq1D_c59, absq1D_c60 :  std_logic_vector(55 downto 0);
signal w0_c60 :  std_logic_vector(55 downto 0);
signal wfinal_c60 :  std_logic_vector(53 downto 0);
signal qM0_c60 :  std_logic;
signal qP28_c0, qP28_c1, qP28_c2, qP28_c3, qP28_c4, qP28_c5, qP28_c6, qP28_c7, qP28_c8, qP28_c9, qP28_c10, qP28_c11, qP28_c12, qP28_c13, qP28_c14, qP28_c15, qP28_c16, qP28_c17, qP28_c18, qP28_c19, qP28_c20, qP28_c21, qP28_c22, qP28_c23, qP28_c24, qP28_c25, qP28_c26, qP28_c27, qP28_c28, qP28_c29, qP28_c30, qP28_c31, qP28_c32, qP28_c33, qP28_c34, qP28_c35, qP28_c36, qP28_c37, qP28_c38, qP28_c39, qP28_c40, qP28_c41, qP28_c42, qP28_c43, qP28_c44, qP28_c45, qP28_c46, qP28_c47, qP28_c48, qP28_c49, qP28_c50, qP28_c51, qP28_c52, qP28_c53, qP28_c54, qP28_c55, qP28_c56, qP28_c57, qP28_c58 :  std_logic_vector(1 downto 0);
signal qM28_c0, qM28_c1, qM28_c2, qM28_c3, qM28_c4, qM28_c5, qM28_c6, qM28_c7, qM28_c8, qM28_c9, qM28_c10, qM28_c11, qM28_c12, qM28_c13, qM28_c14, qM28_c15, qM28_c16, qM28_c17, qM28_c18, qM28_c19, qM28_c20, qM28_c21, qM28_c22, qM28_c23, qM28_c24, qM28_c25, qM28_c26, qM28_c27, qM28_c28, qM28_c29, qM28_c30, qM28_c31, qM28_c32, qM28_c33, qM28_c34, qM28_c35, qM28_c36, qM28_c37, qM28_c38, qM28_c39, qM28_c40, qM28_c41, qM28_c42, qM28_c43, qM28_c44, qM28_c45, qM28_c46, qM28_c47, qM28_c48, qM28_c49, qM28_c50, qM28_c51, qM28_c52, qM28_c53, qM28_c54, qM28_c55, qM28_c56, qM28_c57, qM28_c58, qM28_c59, qM28_c60 :  std_logic_vector(1 downto 0);
signal qP27_c2, qP27_c3, qP27_c4, qP27_c5, qP27_c6, qP27_c7, qP27_c8, qP27_c9, qP27_c10, qP27_c11, qP27_c12, qP27_c13, qP27_c14, qP27_c15, qP27_c16, qP27_c17, qP27_c18, qP27_c19, qP27_c20, qP27_c21, qP27_c22, qP27_c23, qP27_c24, qP27_c25, qP27_c26, qP27_c27, qP27_c28, qP27_c29, qP27_c30, qP27_c31, qP27_c32, qP27_c33, qP27_c34, qP27_c35, qP27_c36, qP27_c37, qP27_c38, qP27_c39, qP27_c40, qP27_c41, qP27_c42, qP27_c43, qP27_c44, qP27_c45, qP27_c46, qP27_c47, qP27_c48, qP27_c49, qP27_c50, qP27_c51, qP27_c52, qP27_c53, qP27_c54, qP27_c55, qP27_c56, qP27_c57, qP27_c58 :  std_logic_vector(1 downto 0);
signal qM27_c2, qM27_c3, qM27_c4, qM27_c5, qM27_c6, qM27_c7, qM27_c8, qM27_c9, qM27_c10, qM27_c11, qM27_c12, qM27_c13, qM27_c14, qM27_c15, qM27_c16, qM27_c17, qM27_c18, qM27_c19, qM27_c20, qM27_c21, qM27_c22, qM27_c23, qM27_c24, qM27_c25, qM27_c26, qM27_c27, qM27_c28, qM27_c29, qM27_c30, qM27_c31, qM27_c32, qM27_c33, qM27_c34, qM27_c35, qM27_c36, qM27_c37, qM27_c38, qM27_c39, qM27_c40, qM27_c41, qM27_c42, qM27_c43, qM27_c44, qM27_c45, qM27_c46, qM27_c47, qM27_c48, qM27_c49, qM27_c50, qM27_c51, qM27_c52, qM27_c53, qM27_c54, qM27_c55, qM27_c56, qM27_c57, qM27_c58, qM27_c59, qM27_c60 :  std_logic_vector(1 downto 0);
signal qP26_c4, qP26_c5, qP26_c6, qP26_c7, qP26_c8, qP26_c9, qP26_c10, qP26_c11, qP26_c12, qP26_c13, qP26_c14, qP26_c15, qP26_c16, qP26_c17, qP26_c18, qP26_c19, qP26_c20, qP26_c21, qP26_c22, qP26_c23, qP26_c24, qP26_c25, qP26_c26, qP26_c27, qP26_c28, qP26_c29, qP26_c30, qP26_c31, qP26_c32, qP26_c33, qP26_c34, qP26_c35, qP26_c36, qP26_c37, qP26_c38, qP26_c39, qP26_c40, qP26_c41, qP26_c42, qP26_c43, qP26_c44, qP26_c45, qP26_c46, qP26_c47, qP26_c48, qP26_c49, qP26_c50, qP26_c51, qP26_c52, qP26_c53, qP26_c54, qP26_c55, qP26_c56, qP26_c57, qP26_c58 :  std_logic_vector(1 downto 0);
signal qM26_c4, qM26_c5, qM26_c6, qM26_c7, qM26_c8, qM26_c9, qM26_c10, qM26_c11, qM26_c12, qM26_c13, qM26_c14, qM26_c15, qM26_c16, qM26_c17, qM26_c18, qM26_c19, qM26_c20, qM26_c21, qM26_c22, qM26_c23, qM26_c24, qM26_c25, qM26_c26, qM26_c27, qM26_c28, qM26_c29, qM26_c30, qM26_c31, qM26_c32, qM26_c33, qM26_c34, qM26_c35, qM26_c36, qM26_c37, qM26_c38, qM26_c39, qM26_c40, qM26_c41, qM26_c42, qM26_c43, qM26_c44, qM26_c45, qM26_c46, qM26_c47, qM26_c48, qM26_c49, qM26_c50, qM26_c51, qM26_c52, qM26_c53, qM26_c54, qM26_c55, qM26_c56, qM26_c57, qM26_c58, qM26_c59, qM26_c60 :  std_logic_vector(1 downto 0);
signal qP25_c6, qP25_c7, qP25_c8, qP25_c9, qP25_c10, qP25_c11, qP25_c12, qP25_c13, qP25_c14, qP25_c15, qP25_c16, qP25_c17, qP25_c18, qP25_c19, qP25_c20, qP25_c21, qP25_c22, qP25_c23, qP25_c24, qP25_c25, qP25_c26, qP25_c27, qP25_c28, qP25_c29, qP25_c30, qP25_c31, qP25_c32, qP25_c33, qP25_c34, qP25_c35, qP25_c36, qP25_c37, qP25_c38, qP25_c39, qP25_c40, qP25_c41, qP25_c42, qP25_c43, qP25_c44, qP25_c45, qP25_c46, qP25_c47, qP25_c48, qP25_c49, qP25_c50, qP25_c51, qP25_c52, qP25_c53, qP25_c54, qP25_c55, qP25_c56, qP25_c57, qP25_c58 :  std_logic_vector(1 downto 0);
signal qM25_c6, qM25_c7, qM25_c8, qM25_c9, qM25_c10, qM25_c11, qM25_c12, qM25_c13, qM25_c14, qM25_c15, qM25_c16, qM25_c17, qM25_c18, qM25_c19, qM25_c20, qM25_c21, qM25_c22, qM25_c23, qM25_c24, qM25_c25, qM25_c26, qM25_c27, qM25_c28, qM25_c29, qM25_c30, qM25_c31, qM25_c32, qM25_c33, qM25_c34, qM25_c35, qM25_c36, qM25_c37, qM25_c38, qM25_c39, qM25_c40, qM25_c41, qM25_c42, qM25_c43, qM25_c44, qM25_c45, qM25_c46, qM25_c47, qM25_c48, qM25_c49, qM25_c50, qM25_c51, qM25_c52, qM25_c53, qM25_c54, qM25_c55, qM25_c56, qM25_c57, qM25_c58, qM25_c59, qM25_c60 :  std_logic_vector(1 downto 0);
signal qP24_c9, qP24_c10, qP24_c11, qP24_c12, qP24_c13, qP24_c14, qP24_c15, qP24_c16, qP24_c17, qP24_c18, qP24_c19, qP24_c20, qP24_c21, qP24_c22, qP24_c23, qP24_c24, qP24_c25, qP24_c26, qP24_c27, qP24_c28, qP24_c29, qP24_c30, qP24_c31, qP24_c32, qP24_c33, qP24_c34, qP24_c35, qP24_c36, qP24_c37, qP24_c38, qP24_c39, qP24_c40, qP24_c41, qP24_c42, qP24_c43, qP24_c44, qP24_c45, qP24_c46, qP24_c47, qP24_c48, qP24_c49, qP24_c50, qP24_c51, qP24_c52, qP24_c53, qP24_c54, qP24_c55, qP24_c56, qP24_c57, qP24_c58 :  std_logic_vector(1 downto 0);
signal qM24_c9, qM24_c10, qM24_c11, qM24_c12, qM24_c13, qM24_c14, qM24_c15, qM24_c16, qM24_c17, qM24_c18, qM24_c19, qM24_c20, qM24_c21, qM24_c22, qM24_c23, qM24_c24, qM24_c25, qM24_c26, qM24_c27, qM24_c28, qM24_c29, qM24_c30, qM24_c31, qM24_c32, qM24_c33, qM24_c34, qM24_c35, qM24_c36, qM24_c37, qM24_c38, qM24_c39, qM24_c40, qM24_c41, qM24_c42, qM24_c43, qM24_c44, qM24_c45, qM24_c46, qM24_c47, qM24_c48, qM24_c49, qM24_c50, qM24_c51, qM24_c52, qM24_c53, qM24_c54, qM24_c55, qM24_c56, qM24_c57, qM24_c58, qM24_c59, qM24_c60 :  std_logic_vector(1 downto 0);
signal qP23_c11, qP23_c12, qP23_c13, qP23_c14, qP23_c15, qP23_c16, qP23_c17, qP23_c18, qP23_c19, qP23_c20, qP23_c21, qP23_c22, qP23_c23, qP23_c24, qP23_c25, qP23_c26, qP23_c27, qP23_c28, qP23_c29, qP23_c30, qP23_c31, qP23_c32, qP23_c33, qP23_c34, qP23_c35, qP23_c36, qP23_c37, qP23_c38, qP23_c39, qP23_c40, qP23_c41, qP23_c42, qP23_c43, qP23_c44, qP23_c45, qP23_c46, qP23_c47, qP23_c48, qP23_c49, qP23_c50, qP23_c51, qP23_c52, qP23_c53, qP23_c54, qP23_c55, qP23_c56, qP23_c57, qP23_c58 :  std_logic_vector(1 downto 0);
signal qM23_c11, qM23_c12, qM23_c13, qM23_c14, qM23_c15, qM23_c16, qM23_c17, qM23_c18, qM23_c19, qM23_c20, qM23_c21, qM23_c22, qM23_c23, qM23_c24, qM23_c25, qM23_c26, qM23_c27, qM23_c28, qM23_c29, qM23_c30, qM23_c31, qM23_c32, qM23_c33, qM23_c34, qM23_c35, qM23_c36, qM23_c37, qM23_c38, qM23_c39, qM23_c40, qM23_c41, qM23_c42, qM23_c43, qM23_c44, qM23_c45, qM23_c46, qM23_c47, qM23_c48, qM23_c49, qM23_c50, qM23_c51, qM23_c52, qM23_c53, qM23_c54, qM23_c55, qM23_c56, qM23_c57, qM23_c58, qM23_c59, qM23_c60 :  std_logic_vector(1 downto 0);
signal qP22_c13, qP22_c14, qP22_c15, qP22_c16, qP22_c17, qP22_c18, qP22_c19, qP22_c20, qP22_c21, qP22_c22, qP22_c23, qP22_c24, qP22_c25, qP22_c26, qP22_c27, qP22_c28, qP22_c29, qP22_c30, qP22_c31, qP22_c32, qP22_c33, qP22_c34, qP22_c35, qP22_c36, qP22_c37, qP22_c38, qP22_c39, qP22_c40, qP22_c41, qP22_c42, qP22_c43, qP22_c44, qP22_c45, qP22_c46, qP22_c47, qP22_c48, qP22_c49, qP22_c50, qP22_c51, qP22_c52, qP22_c53, qP22_c54, qP22_c55, qP22_c56, qP22_c57, qP22_c58 :  std_logic_vector(1 downto 0);
signal qM22_c13, qM22_c14, qM22_c15, qM22_c16, qM22_c17, qM22_c18, qM22_c19, qM22_c20, qM22_c21, qM22_c22, qM22_c23, qM22_c24, qM22_c25, qM22_c26, qM22_c27, qM22_c28, qM22_c29, qM22_c30, qM22_c31, qM22_c32, qM22_c33, qM22_c34, qM22_c35, qM22_c36, qM22_c37, qM22_c38, qM22_c39, qM22_c40, qM22_c41, qM22_c42, qM22_c43, qM22_c44, qM22_c45, qM22_c46, qM22_c47, qM22_c48, qM22_c49, qM22_c50, qM22_c51, qM22_c52, qM22_c53, qM22_c54, qM22_c55, qM22_c56, qM22_c57, qM22_c58, qM22_c59, qM22_c60 :  std_logic_vector(1 downto 0);
signal qP21_c15, qP21_c16, qP21_c17, qP21_c18, qP21_c19, qP21_c20, qP21_c21, qP21_c22, qP21_c23, qP21_c24, qP21_c25, qP21_c26, qP21_c27, qP21_c28, qP21_c29, qP21_c30, qP21_c31, qP21_c32, qP21_c33, qP21_c34, qP21_c35, qP21_c36, qP21_c37, qP21_c38, qP21_c39, qP21_c40, qP21_c41, qP21_c42, qP21_c43, qP21_c44, qP21_c45, qP21_c46, qP21_c47, qP21_c48, qP21_c49, qP21_c50, qP21_c51, qP21_c52, qP21_c53, qP21_c54, qP21_c55, qP21_c56, qP21_c57, qP21_c58 :  std_logic_vector(1 downto 0);
signal qM21_c15, qM21_c16, qM21_c17, qM21_c18, qM21_c19, qM21_c20, qM21_c21, qM21_c22, qM21_c23, qM21_c24, qM21_c25, qM21_c26, qM21_c27, qM21_c28, qM21_c29, qM21_c30, qM21_c31, qM21_c32, qM21_c33, qM21_c34, qM21_c35, qM21_c36, qM21_c37, qM21_c38, qM21_c39, qM21_c40, qM21_c41, qM21_c42, qM21_c43, qM21_c44, qM21_c45, qM21_c46, qM21_c47, qM21_c48, qM21_c49, qM21_c50, qM21_c51, qM21_c52, qM21_c53, qM21_c54, qM21_c55, qM21_c56, qM21_c57, qM21_c58, qM21_c59, qM21_c60 :  std_logic_vector(1 downto 0);
signal qP20_c17, qP20_c18, qP20_c19, qP20_c20, qP20_c21, qP20_c22, qP20_c23, qP20_c24, qP20_c25, qP20_c26, qP20_c27, qP20_c28, qP20_c29, qP20_c30, qP20_c31, qP20_c32, qP20_c33, qP20_c34, qP20_c35, qP20_c36, qP20_c37, qP20_c38, qP20_c39, qP20_c40, qP20_c41, qP20_c42, qP20_c43, qP20_c44, qP20_c45, qP20_c46, qP20_c47, qP20_c48, qP20_c49, qP20_c50, qP20_c51, qP20_c52, qP20_c53, qP20_c54, qP20_c55, qP20_c56, qP20_c57, qP20_c58 :  std_logic_vector(1 downto 0);
signal qM20_c17, qM20_c18, qM20_c19, qM20_c20, qM20_c21, qM20_c22, qM20_c23, qM20_c24, qM20_c25, qM20_c26, qM20_c27, qM20_c28, qM20_c29, qM20_c30, qM20_c31, qM20_c32, qM20_c33, qM20_c34, qM20_c35, qM20_c36, qM20_c37, qM20_c38, qM20_c39, qM20_c40, qM20_c41, qM20_c42, qM20_c43, qM20_c44, qM20_c45, qM20_c46, qM20_c47, qM20_c48, qM20_c49, qM20_c50, qM20_c51, qM20_c52, qM20_c53, qM20_c54, qM20_c55, qM20_c56, qM20_c57, qM20_c58, qM20_c59, qM20_c60 :  std_logic_vector(1 downto 0);
signal qP19_c19, qP19_c20, qP19_c21, qP19_c22, qP19_c23, qP19_c24, qP19_c25, qP19_c26, qP19_c27, qP19_c28, qP19_c29, qP19_c30, qP19_c31, qP19_c32, qP19_c33, qP19_c34, qP19_c35, qP19_c36, qP19_c37, qP19_c38, qP19_c39, qP19_c40, qP19_c41, qP19_c42, qP19_c43, qP19_c44, qP19_c45, qP19_c46, qP19_c47, qP19_c48, qP19_c49, qP19_c50, qP19_c51, qP19_c52, qP19_c53, qP19_c54, qP19_c55, qP19_c56, qP19_c57, qP19_c58 :  std_logic_vector(1 downto 0);
signal qM19_c19, qM19_c20, qM19_c21, qM19_c22, qM19_c23, qM19_c24, qM19_c25, qM19_c26, qM19_c27, qM19_c28, qM19_c29, qM19_c30, qM19_c31, qM19_c32, qM19_c33, qM19_c34, qM19_c35, qM19_c36, qM19_c37, qM19_c38, qM19_c39, qM19_c40, qM19_c41, qM19_c42, qM19_c43, qM19_c44, qM19_c45, qM19_c46, qM19_c47, qM19_c48, qM19_c49, qM19_c50, qM19_c51, qM19_c52, qM19_c53, qM19_c54, qM19_c55, qM19_c56, qM19_c57, qM19_c58, qM19_c59, qM19_c60 :  std_logic_vector(1 downto 0);
signal qP18_c22, qP18_c23, qP18_c24, qP18_c25, qP18_c26, qP18_c27, qP18_c28, qP18_c29, qP18_c30, qP18_c31, qP18_c32, qP18_c33, qP18_c34, qP18_c35, qP18_c36, qP18_c37, qP18_c38, qP18_c39, qP18_c40, qP18_c41, qP18_c42, qP18_c43, qP18_c44, qP18_c45, qP18_c46, qP18_c47, qP18_c48, qP18_c49, qP18_c50, qP18_c51, qP18_c52, qP18_c53, qP18_c54, qP18_c55, qP18_c56, qP18_c57, qP18_c58 :  std_logic_vector(1 downto 0);
signal qM18_c22, qM18_c23, qM18_c24, qM18_c25, qM18_c26, qM18_c27, qM18_c28, qM18_c29, qM18_c30, qM18_c31, qM18_c32, qM18_c33, qM18_c34, qM18_c35, qM18_c36, qM18_c37, qM18_c38, qM18_c39, qM18_c40, qM18_c41, qM18_c42, qM18_c43, qM18_c44, qM18_c45, qM18_c46, qM18_c47, qM18_c48, qM18_c49, qM18_c50, qM18_c51, qM18_c52, qM18_c53, qM18_c54, qM18_c55, qM18_c56, qM18_c57, qM18_c58, qM18_c59, qM18_c60 :  std_logic_vector(1 downto 0);
signal qP17_c24, qP17_c25, qP17_c26, qP17_c27, qP17_c28, qP17_c29, qP17_c30, qP17_c31, qP17_c32, qP17_c33, qP17_c34, qP17_c35, qP17_c36, qP17_c37, qP17_c38, qP17_c39, qP17_c40, qP17_c41, qP17_c42, qP17_c43, qP17_c44, qP17_c45, qP17_c46, qP17_c47, qP17_c48, qP17_c49, qP17_c50, qP17_c51, qP17_c52, qP17_c53, qP17_c54, qP17_c55, qP17_c56, qP17_c57, qP17_c58 :  std_logic_vector(1 downto 0);
signal qM17_c24, qM17_c25, qM17_c26, qM17_c27, qM17_c28, qM17_c29, qM17_c30, qM17_c31, qM17_c32, qM17_c33, qM17_c34, qM17_c35, qM17_c36, qM17_c37, qM17_c38, qM17_c39, qM17_c40, qM17_c41, qM17_c42, qM17_c43, qM17_c44, qM17_c45, qM17_c46, qM17_c47, qM17_c48, qM17_c49, qM17_c50, qM17_c51, qM17_c52, qM17_c53, qM17_c54, qM17_c55, qM17_c56, qM17_c57, qM17_c58, qM17_c59, qM17_c60 :  std_logic_vector(1 downto 0);
signal qP16_c26, qP16_c27, qP16_c28, qP16_c29, qP16_c30, qP16_c31, qP16_c32, qP16_c33, qP16_c34, qP16_c35, qP16_c36, qP16_c37, qP16_c38, qP16_c39, qP16_c40, qP16_c41, qP16_c42, qP16_c43, qP16_c44, qP16_c45, qP16_c46, qP16_c47, qP16_c48, qP16_c49, qP16_c50, qP16_c51, qP16_c52, qP16_c53, qP16_c54, qP16_c55, qP16_c56, qP16_c57, qP16_c58 :  std_logic_vector(1 downto 0);
signal qM16_c26, qM16_c27, qM16_c28, qM16_c29, qM16_c30, qM16_c31, qM16_c32, qM16_c33, qM16_c34, qM16_c35, qM16_c36, qM16_c37, qM16_c38, qM16_c39, qM16_c40, qM16_c41, qM16_c42, qM16_c43, qM16_c44, qM16_c45, qM16_c46, qM16_c47, qM16_c48, qM16_c49, qM16_c50, qM16_c51, qM16_c52, qM16_c53, qM16_c54, qM16_c55, qM16_c56, qM16_c57, qM16_c58, qM16_c59, qM16_c60 :  std_logic_vector(1 downto 0);
signal qP15_c28, qP15_c29, qP15_c30, qP15_c31, qP15_c32, qP15_c33, qP15_c34, qP15_c35, qP15_c36, qP15_c37, qP15_c38, qP15_c39, qP15_c40, qP15_c41, qP15_c42, qP15_c43, qP15_c44, qP15_c45, qP15_c46, qP15_c47, qP15_c48, qP15_c49, qP15_c50, qP15_c51, qP15_c52, qP15_c53, qP15_c54, qP15_c55, qP15_c56, qP15_c57, qP15_c58 :  std_logic_vector(1 downto 0);
signal qM15_c28, qM15_c29, qM15_c30, qM15_c31, qM15_c32, qM15_c33, qM15_c34, qM15_c35, qM15_c36, qM15_c37, qM15_c38, qM15_c39, qM15_c40, qM15_c41, qM15_c42, qM15_c43, qM15_c44, qM15_c45, qM15_c46, qM15_c47, qM15_c48, qM15_c49, qM15_c50, qM15_c51, qM15_c52, qM15_c53, qM15_c54, qM15_c55, qM15_c56, qM15_c57, qM15_c58, qM15_c59, qM15_c60 :  std_logic_vector(1 downto 0);
signal qP14_c30, qP14_c31, qP14_c32, qP14_c33, qP14_c34, qP14_c35, qP14_c36, qP14_c37, qP14_c38, qP14_c39, qP14_c40, qP14_c41, qP14_c42, qP14_c43, qP14_c44, qP14_c45, qP14_c46, qP14_c47, qP14_c48, qP14_c49, qP14_c50, qP14_c51, qP14_c52, qP14_c53, qP14_c54, qP14_c55, qP14_c56, qP14_c57, qP14_c58 :  std_logic_vector(1 downto 0);
signal qM14_c30, qM14_c31, qM14_c32, qM14_c33, qM14_c34, qM14_c35, qM14_c36, qM14_c37, qM14_c38, qM14_c39, qM14_c40, qM14_c41, qM14_c42, qM14_c43, qM14_c44, qM14_c45, qM14_c46, qM14_c47, qM14_c48, qM14_c49, qM14_c50, qM14_c51, qM14_c52, qM14_c53, qM14_c54, qM14_c55, qM14_c56, qM14_c57, qM14_c58, qM14_c59, qM14_c60 :  std_logic_vector(1 downto 0);
signal qP13_c32, qP13_c33, qP13_c34, qP13_c35, qP13_c36, qP13_c37, qP13_c38, qP13_c39, qP13_c40, qP13_c41, qP13_c42, qP13_c43, qP13_c44, qP13_c45, qP13_c46, qP13_c47, qP13_c48, qP13_c49, qP13_c50, qP13_c51, qP13_c52, qP13_c53, qP13_c54, qP13_c55, qP13_c56, qP13_c57, qP13_c58 :  std_logic_vector(1 downto 0);
signal qM13_c32, qM13_c33, qM13_c34, qM13_c35, qM13_c36, qM13_c37, qM13_c38, qM13_c39, qM13_c40, qM13_c41, qM13_c42, qM13_c43, qM13_c44, qM13_c45, qM13_c46, qM13_c47, qM13_c48, qM13_c49, qM13_c50, qM13_c51, qM13_c52, qM13_c53, qM13_c54, qM13_c55, qM13_c56, qM13_c57, qM13_c58, qM13_c59, qM13_c60 :  std_logic_vector(1 downto 0);
signal qP12_c34, qP12_c35, qP12_c36, qP12_c37, qP12_c38, qP12_c39, qP12_c40, qP12_c41, qP12_c42, qP12_c43, qP12_c44, qP12_c45, qP12_c46, qP12_c47, qP12_c48, qP12_c49, qP12_c50, qP12_c51, qP12_c52, qP12_c53, qP12_c54, qP12_c55, qP12_c56, qP12_c57, qP12_c58 :  std_logic_vector(1 downto 0);
signal qM12_c34, qM12_c35, qM12_c36, qM12_c37, qM12_c38, qM12_c39, qM12_c40, qM12_c41, qM12_c42, qM12_c43, qM12_c44, qM12_c45, qM12_c46, qM12_c47, qM12_c48, qM12_c49, qM12_c50, qM12_c51, qM12_c52, qM12_c53, qM12_c54, qM12_c55, qM12_c56, qM12_c57, qM12_c58, qM12_c59, qM12_c60 :  std_logic_vector(1 downto 0);
signal qP11_c37, qP11_c38, qP11_c39, qP11_c40, qP11_c41, qP11_c42, qP11_c43, qP11_c44, qP11_c45, qP11_c46, qP11_c47, qP11_c48, qP11_c49, qP11_c50, qP11_c51, qP11_c52, qP11_c53, qP11_c54, qP11_c55, qP11_c56, qP11_c57, qP11_c58 :  std_logic_vector(1 downto 0);
signal qM11_c37, qM11_c38, qM11_c39, qM11_c40, qM11_c41, qM11_c42, qM11_c43, qM11_c44, qM11_c45, qM11_c46, qM11_c47, qM11_c48, qM11_c49, qM11_c50, qM11_c51, qM11_c52, qM11_c53, qM11_c54, qM11_c55, qM11_c56, qM11_c57, qM11_c58, qM11_c59, qM11_c60 :  std_logic_vector(1 downto 0);
signal qP10_c39, qP10_c40, qP10_c41, qP10_c42, qP10_c43, qP10_c44, qP10_c45, qP10_c46, qP10_c47, qP10_c48, qP10_c49, qP10_c50, qP10_c51, qP10_c52, qP10_c53, qP10_c54, qP10_c55, qP10_c56, qP10_c57, qP10_c58 :  std_logic_vector(1 downto 0);
signal qM10_c39, qM10_c40, qM10_c41, qM10_c42, qM10_c43, qM10_c44, qM10_c45, qM10_c46, qM10_c47, qM10_c48, qM10_c49, qM10_c50, qM10_c51, qM10_c52, qM10_c53, qM10_c54, qM10_c55, qM10_c56, qM10_c57, qM10_c58, qM10_c59, qM10_c60 :  std_logic_vector(1 downto 0);
signal qP9_c41, qP9_c42, qP9_c43, qP9_c44, qP9_c45, qP9_c46, qP9_c47, qP9_c48, qP9_c49, qP9_c50, qP9_c51, qP9_c52, qP9_c53, qP9_c54, qP9_c55, qP9_c56, qP9_c57, qP9_c58 :  std_logic_vector(1 downto 0);
signal qM9_c41, qM9_c42, qM9_c43, qM9_c44, qM9_c45, qM9_c46, qM9_c47, qM9_c48, qM9_c49, qM9_c50, qM9_c51, qM9_c52, qM9_c53, qM9_c54, qM9_c55, qM9_c56, qM9_c57, qM9_c58, qM9_c59, qM9_c60 :  std_logic_vector(1 downto 0);
signal qP8_c43, qP8_c44, qP8_c45, qP8_c46, qP8_c47, qP8_c48, qP8_c49, qP8_c50, qP8_c51, qP8_c52, qP8_c53, qP8_c54, qP8_c55, qP8_c56, qP8_c57, qP8_c58 :  std_logic_vector(1 downto 0);
signal qM8_c43, qM8_c44, qM8_c45, qM8_c46, qM8_c47, qM8_c48, qM8_c49, qM8_c50, qM8_c51, qM8_c52, qM8_c53, qM8_c54, qM8_c55, qM8_c56, qM8_c57, qM8_c58, qM8_c59, qM8_c60 :  std_logic_vector(1 downto 0);
signal qP7_c45, qP7_c46, qP7_c47, qP7_c48, qP7_c49, qP7_c50, qP7_c51, qP7_c52, qP7_c53, qP7_c54, qP7_c55, qP7_c56, qP7_c57, qP7_c58 :  std_logic_vector(1 downto 0);
signal qM7_c45, qM7_c46, qM7_c47, qM7_c48, qM7_c49, qM7_c50, qM7_c51, qM7_c52, qM7_c53, qM7_c54, qM7_c55, qM7_c56, qM7_c57, qM7_c58, qM7_c59, qM7_c60 :  std_logic_vector(1 downto 0);
signal qP6_c47, qP6_c48, qP6_c49, qP6_c50, qP6_c51, qP6_c52, qP6_c53, qP6_c54, qP6_c55, qP6_c56, qP6_c57, qP6_c58 :  std_logic_vector(1 downto 0);
signal qM6_c47, qM6_c48, qM6_c49, qM6_c50, qM6_c51, qM6_c52, qM6_c53, qM6_c54, qM6_c55, qM6_c56, qM6_c57, qM6_c58, qM6_c59, qM6_c60 :  std_logic_vector(1 downto 0);
signal qP5_c49, qP5_c50, qP5_c51, qP5_c52, qP5_c53, qP5_c54, qP5_c55, qP5_c56, qP5_c57, qP5_c58 :  std_logic_vector(1 downto 0);
signal qM5_c49, qM5_c50, qM5_c51, qM5_c52, qM5_c53, qM5_c54, qM5_c55, qM5_c56, qM5_c57, qM5_c58, qM5_c59, qM5_c60 :  std_logic_vector(1 downto 0);
signal qP4_c52, qP4_c53, qP4_c54, qP4_c55, qP4_c56, qP4_c57, qP4_c58 :  std_logic_vector(1 downto 0);
signal qM4_c52, qM4_c53, qM4_c54, qM4_c55, qM4_c56, qM4_c57, qM4_c58, qM4_c59, qM4_c60 :  std_logic_vector(1 downto 0);
signal qP3_c54, qP3_c55, qP3_c56, qP3_c57, qP3_c58 :  std_logic_vector(1 downto 0);
signal qM3_c54, qM3_c55, qM3_c56, qM3_c57, qM3_c58, qM3_c59, qM3_c60 :  std_logic_vector(1 downto 0);
signal qP2_c56, qP2_c57, qP2_c58 :  std_logic_vector(1 downto 0);
signal qM2_c56, qM2_c57, qM2_c58, qM2_c59, qM2_c60 :  std_logic_vector(1 downto 0);
signal qP1_c58 :  std_logic_vector(1 downto 0);
signal qM1_c58, qM1_c59, qM1_c60 :  std_logic_vector(1 downto 0);
signal qP_c58, qP_c59, qP_c60, qP_c61 :  std_logic_vector(55 downto 0);
signal qM_c60, qM_c61 :  std_logic_vector(55 downto 0);
signal quotient_c61 :  std_logic_vector(55 downto 0);
signal mR_c61, mR_c62 :  std_logic_vector(54 downto 0);
signal fRnorm_c61, fRnorm_c62 :  std_logic_vector(52 downto 0);
signal round_c61, round_c62 :  std_logic;
signal expR1_c62 :  std_logic_vector(12 downto 0);
signal expfrac_c62 :  std_logic_vector(64 downto 0);
signal expfracR_c62, expfracR_c63 :  std_logic_vector(64 downto 0);
signal exnR_c63 :  std_logic_vector(1 downto 0);
signal exnRfinal_c63 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               expR0_c1 <= expR0_c0;
               sR_c1 <= sR_c0;
               exnR0_c1 <= exnR0_c0;
               D_c1 <= D_c0;
               betaw28_c1 <= betaw28_c0;
               q28_c1 <= q28_c0;
               absq28D_c1 <= absq28D_c0;
               qP28_c1 <= qP28_c0;
               qM28_c1 <= qM28_c0;
            end if;
            if ce_2 = '1' then
               expR0_c2 <= expR0_c1;
               sR_c2 <= sR_c1;
               exnR0_c2 <= exnR0_c1;
               D_c2 <= D_c1;
               betaw28_c2 <= betaw28_c1;
               q28_c2 <= q28_c1;
               absq28D_c2 <= absq28D_c1;
               qP28_c2 <= qP28_c1;
               qM28_c2 <= qM28_c1;
            end if;
            if ce_3 = '1' then
               expR0_c3 <= expR0_c2;
               sR_c3 <= sR_c2;
               exnR0_c3 <= exnR0_c2;
               D_c3 <= D_c2;
               betaw27_c3 <= betaw27_c2;
               q27_c3 <= q27_c2;
               absq27D_c3 <= absq27D_c2;
               qP28_c3 <= qP28_c2;
               qM28_c3 <= qM28_c2;
               qP27_c3 <= qP27_c2;
               qM27_c3 <= qM27_c2;
            end if;
            if ce_4 = '1' then
               expR0_c4 <= expR0_c3;
               sR_c4 <= sR_c3;
               exnR0_c4 <= exnR0_c3;
               D_c4 <= D_c3;
               betaw27_c4 <= betaw27_c3;
               q27_c4 <= q27_c3;
               absq27D_c4 <= absq27D_c3;
               qP28_c4 <= qP28_c3;
               qM28_c4 <= qM28_c3;
               qP27_c4 <= qP27_c3;
               qM27_c4 <= qM27_c3;
            end if;
            if ce_5 = '1' then
               expR0_c5 <= expR0_c4;
               sR_c5 <= sR_c4;
               exnR0_c5 <= exnR0_c4;
               D_c5 <= D_c4;
               betaw26_c5 <= betaw26_c4;
               q26_c5 <= q26_c4;
               absq26D_c5 <= absq26D_c4;
               qP28_c5 <= qP28_c4;
               qM28_c5 <= qM28_c4;
               qP27_c5 <= qP27_c4;
               qM27_c5 <= qM27_c4;
               qP26_c5 <= qP26_c4;
               qM26_c5 <= qM26_c4;
            end if;
            if ce_6 = '1' then
               expR0_c6 <= expR0_c5;
               sR_c6 <= sR_c5;
               exnR0_c6 <= exnR0_c5;
               D_c6 <= D_c5;
               betaw26_c6 <= betaw26_c5;
               q26_c6 <= q26_c5;
               absq26D_c6 <= absq26D_c5;
               qP28_c6 <= qP28_c5;
               qM28_c6 <= qM28_c5;
               qP27_c6 <= qP27_c5;
               qM27_c6 <= qM27_c5;
               qP26_c6 <= qP26_c5;
               qM26_c6 <= qM26_c5;
            end if;
            if ce_7 = '1' then
               expR0_c7 <= expR0_c6;
               sR_c7 <= sR_c6;
               exnR0_c7 <= exnR0_c6;
               D_c7 <= D_c6;
               betaw25_c7 <= betaw25_c6;
               q25_c7 <= q25_c6;
               absq25D_c7 <= absq25D_c6;
               qP28_c7 <= qP28_c6;
               qM28_c7 <= qM28_c6;
               qP27_c7 <= qP27_c6;
               qM27_c7 <= qM27_c6;
               qP26_c7 <= qP26_c6;
               qM26_c7 <= qM26_c6;
               qP25_c7 <= qP25_c6;
               qM25_c7 <= qM25_c6;
            end if;
            if ce_8 = '1' then
               expR0_c8 <= expR0_c7;
               sR_c8 <= sR_c7;
               exnR0_c8 <= exnR0_c7;
               D_c8 <= D_c7;
               betaw25_c8 <= betaw25_c7;
               q25_c8 <= q25_c7;
               absq25D_c8 <= absq25D_c7;
               qP28_c8 <= qP28_c7;
               qM28_c8 <= qM28_c7;
               qP27_c8 <= qP27_c7;
               qM27_c8 <= qM27_c7;
               qP26_c8 <= qP26_c7;
               qM26_c8 <= qM26_c7;
               qP25_c8 <= qP25_c7;
               qM25_c8 <= qM25_c7;
            end if;
            if ce_9 = '1' then
               expR0_c9 <= expR0_c8;
               sR_c9 <= sR_c8;
               exnR0_c9 <= exnR0_c8;
               D_c9 <= D_c8;
               betaw24_c9 <= betaw24_c8;
               q24_copy9_c9 <= q24_copy9_c8;
               qP28_c9 <= qP28_c8;
               qM28_c9 <= qM28_c8;
               qP27_c9 <= qP27_c8;
               qM27_c9 <= qM27_c8;
               qP26_c9 <= qP26_c8;
               qM26_c9 <= qM26_c8;
               qP25_c9 <= qP25_c8;
               qM25_c9 <= qM25_c8;
            end if;
            if ce_10 = '1' then
               expR0_c10 <= expR0_c9;
               sR_c10 <= sR_c9;
               exnR0_c10 <= exnR0_c9;
               D_c10 <= D_c9;
               betaw24_c10 <= betaw24_c9;
               q24_c10 <= q24_c9;
               absq24D_c10 <= absq24D_c9;
               qP28_c10 <= qP28_c9;
               qM28_c10 <= qM28_c9;
               qP27_c10 <= qP27_c9;
               qM27_c10 <= qM27_c9;
               qP26_c10 <= qP26_c9;
               qM26_c10 <= qM26_c9;
               qP25_c10 <= qP25_c9;
               qM25_c10 <= qM25_c9;
               qP24_c10 <= qP24_c9;
               qM24_c10 <= qM24_c9;
            end if;
            if ce_11 = '1' then
               expR0_c11 <= expR0_c10;
               sR_c11 <= sR_c10;
               exnR0_c11 <= exnR0_c10;
               D_c11 <= D_c10;
               betaw23_c11 <= betaw23_c10;
               q23_copy10_c11 <= q23_copy10_c10;
               qP28_c11 <= qP28_c10;
               qM28_c11 <= qM28_c10;
               qP27_c11 <= qP27_c10;
               qM27_c11 <= qM27_c10;
               qP26_c11 <= qP26_c10;
               qM26_c11 <= qM26_c10;
               qP25_c11 <= qP25_c10;
               qM25_c11 <= qM25_c10;
               qP24_c11 <= qP24_c10;
               qM24_c11 <= qM24_c10;
            end if;
            if ce_12 = '1' then
               expR0_c12 <= expR0_c11;
               sR_c12 <= sR_c11;
               exnR0_c12 <= exnR0_c11;
               D_c12 <= D_c11;
               betaw23_c12 <= betaw23_c11;
               q23_c12 <= q23_c11;
               absq23D_c12 <= absq23D_c11;
               qP28_c12 <= qP28_c11;
               qM28_c12 <= qM28_c11;
               qP27_c12 <= qP27_c11;
               qM27_c12 <= qM27_c11;
               qP26_c12 <= qP26_c11;
               qM26_c12 <= qM26_c11;
               qP25_c12 <= qP25_c11;
               qM25_c12 <= qM25_c11;
               qP24_c12 <= qP24_c11;
               qM24_c12 <= qM24_c11;
               qP23_c12 <= qP23_c11;
               qM23_c12 <= qM23_c11;
            end if;
            if ce_13 = '1' then
               expR0_c13 <= expR0_c12;
               sR_c13 <= sR_c12;
               exnR0_c13 <= exnR0_c12;
               D_c13 <= D_c12;
               betaw22_c13 <= betaw22_c12;
               q22_copy11_c13 <= q22_copy11_c12;
               qP28_c13 <= qP28_c12;
               qM28_c13 <= qM28_c12;
               qP27_c13 <= qP27_c12;
               qM27_c13 <= qM27_c12;
               qP26_c13 <= qP26_c12;
               qM26_c13 <= qM26_c12;
               qP25_c13 <= qP25_c12;
               qM25_c13 <= qM25_c12;
               qP24_c13 <= qP24_c12;
               qM24_c13 <= qM24_c12;
               qP23_c13 <= qP23_c12;
               qM23_c13 <= qM23_c12;
            end if;
            if ce_14 = '1' then
               expR0_c14 <= expR0_c13;
               sR_c14 <= sR_c13;
               exnR0_c14 <= exnR0_c13;
               D_c14 <= D_c13;
               betaw22_c14 <= betaw22_c13;
               q22_c14 <= q22_c13;
               absq22D_c14 <= absq22D_c13;
               qP28_c14 <= qP28_c13;
               qM28_c14 <= qM28_c13;
               qP27_c14 <= qP27_c13;
               qM27_c14 <= qM27_c13;
               qP26_c14 <= qP26_c13;
               qM26_c14 <= qM26_c13;
               qP25_c14 <= qP25_c13;
               qM25_c14 <= qM25_c13;
               qP24_c14 <= qP24_c13;
               qM24_c14 <= qM24_c13;
               qP23_c14 <= qP23_c13;
               qM23_c14 <= qM23_c13;
               qP22_c14 <= qP22_c13;
               qM22_c14 <= qM22_c13;
            end if;
            if ce_15 = '1' then
               expR0_c15 <= expR0_c14;
               sR_c15 <= sR_c14;
               exnR0_c15 <= exnR0_c14;
               D_c15 <= D_c14;
               betaw22_c15 <= betaw22_c14;
               q22_c15 <= q22_c14;
               absq22D_c15 <= absq22D_c14;
               qP28_c15 <= qP28_c14;
               qM28_c15 <= qM28_c14;
               qP27_c15 <= qP27_c14;
               qM27_c15 <= qM27_c14;
               qP26_c15 <= qP26_c14;
               qM26_c15 <= qM26_c14;
               qP25_c15 <= qP25_c14;
               qM25_c15 <= qM25_c14;
               qP24_c15 <= qP24_c14;
               qM24_c15 <= qM24_c14;
               qP23_c15 <= qP23_c14;
               qM23_c15 <= qM23_c14;
               qP22_c15 <= qP22_c14;
               qM22_c15 <= qM22_c14;
            end if;
            if ce_16 = '1' then
               expR0_c16 <= expR0_c15;
               sR_c16 <= sR_c15;
               exnR0_c16 <= exnR0_c15;
               D_c16 <= D_c15;
               betaw21_c16 <= betaw21_c15;
               q21_c16 <= q21_c15;
               absq21D_c16 <= absq21D_c15;
               qP28_c16 <= qP28_c15;
               qM28_c16 <= qM28_c15;
               qP27_c16 <= qP27_c15;
               qM27_c16 <= qM27_c15;
               qP26_c16 <= qP26_c15;
               qM26_c16 <= qM26_c15;
               qP25_c16 <= qP25_c15;
               qM25_c16 <= qM25_c15;
               qP24_c16 <= qP24_c15;
               qM24_c16 <= qM24_c15;
               qP23_c16 <= qP23_c15;
               qM23_c16 <= qM23_c15;
               qP22_c16 <= qP22_c15;
               qM22_c16 <= qM22_c15;
               qP21_c16 <= qP21_c15;
               qM21_c16 <= qM21_c15;
            end if;
            if ce_17 = '1' then
               expR0_c17 <= expR0_c16;
               sR_c17 <= sR_c16;
               exnR0_c17 <= exnR0_c16;
               D_c17 <= D_c16;
               betaw21_c17 <= betaw21_c16;
               q21_c17 <= q21_c16;
               absq21D_c17 <= absq21D_c16;
               qP28_c17 <= qP28_c16;
               qM28_c17 <= qM28_c16;
               qP27_c17 <= qP27_c16;
               qM27_c17 <= qM27_c16;
               qP26_c17 <= qP26_c16;
               qM26_c17 <= qM26_c16;
               qP25_c17 <= qP25_c16;
               qM25_c17 <= qM25_c16;
               qP24_c17 <= qP24_c16;
               qM24_c17 <= qM24_c16;
               qP23_c17 <= qP23_c16;
               qM23_c17 <= qM23_c16;
               qP22_c17 <= qP22_c16;
               qM22_c17 <= qM22_c16;
               qP21_c17 <= qP21_c16;
               qM21_c17 <= qM21_c16;
            end if;
            if ce_18 = '1' then
               expR0_c18 <= expR0_c17;
               sR_c18 <= sR_c17;
               exnR0_c18 <= exnR0_c17;
               D_c18 <= D_c17;
               betaw20_c18 <= betaw20_c17;
               q20_c18 <= q20_c17;
               absq20D_c18 <= absq20D_c17;
               qP28_c18 <= qP28_c17;
               qM28_c18 <= qM28_c17;
               qP27_c18 <= qP27_c17;
               qM27_c18 <= qM27_c17;
               qP26_c18 <= qP26_c17;
               qM26_c18 <= qM26_c17;
               qP25_c18 <= qP25_c17;
               qM25_c18 <= qM25_c17;
               qP24_c18 <= qP24_c17;
               qM24_c18 <= qM24_c17;
               qP23_c18 <= qP23_c17;
               qM23_c18 <= qM23_c17;
               qP22_c18 <= qP22_c17;
               qM22_c18 <= qM22_c17;
               qP21_c18 <= qP21_c17;
               qM21_c18 <= qM21_c17;
               qP20_c18 <= qP20_c17;
               qM20_c18 <= qM20_c17;
            end if;
            if ce_19 = '1' then
               expR0_c19 <= expR0_c18;
               sR_c19 <= sR_c18;
               exnR0_c19 <= exnR0_c18;
               D_c19 <= D_c18;
               betaw20_c19 <= betaw20_c18;
               q20_c19 <= q20_c18;
               absq20D_c19 <= absq20D_c18;
               qP28_c19 <= qP28_c18;
               qM28_c19 <= qM28_c18;
               qP27_c19 <= qP27_c18;
               qM27_c19 <= qM27_c18;
               qP26_c19 <= qP26_c18;
               qM26_c19 <= qM26_c18;
               qP25_c19 <= qP25_c18;
               qM25_c19 <= qM25_c18;
               qP24_c19 <= qP24_c18;
               qM24_c19 <= qM24_c18;
               qP23_c19 <= qP23_c18;
               qM23_c19 <= qM23_c18;
               qP22_c19 <= qP22_c18;
               qM22_c19 <= qM22_c18;
               qP21_c19 <= qP21_c18;
               qM21_c19 <= qM21_c18;
               qP20_c19 <= qP20_c18;
               qM20_c19 <= qM20_c18;
            end if;
            if ce_20 = '1' then
               expR0_c20 <= expR0_c19;
               sR_c20 <= sR_c19;
               exnR0_c20 <= exnR0_c19;
               D_c20 <= D_c19;
               betaw19_c20 <= betaw19_c19;
               q19_c20 <= q19_c19;
               absq19D_c20 <= absq19D_c19;
               qP28_c20 <= qP28_c19;
               qM28_c20 <= qM28_c19;
               qP27_c20 <= qP27_c19;
               qM27_c20 <= qM27_c19;
               qP26_c20 <= qP26_c19;
               qM26_c20 <= qM26_c19;
               qP25_c20 <= qP25_c19;
               qM25_c20 <= qM25_c19;
               qP24_c20 <= qP24_c19;
               qM24_c20 <= qM24_c19;
               qP23_c20 <= qP23_c19;
               qM23_c20 <= qM23_c19;
               qP22_c20 <= qP22_c19;
               qM22_c20 <= qM22_c19;
               qP21_c20 <= qP21_c19;
               qM21_c20 <= qM21_c19;
               qP20_c20 <= qP20_c19;
               qM20_c20 <= qM20_c19;
               qP19_c20 <= qP19_c19;
               qM19_c20 <= qM19_c19;
            end if;
            if ce_21 = '1' then
               expR0_c21 <= expR0_c20;
               sR_c21 <= sR_c20;
               exnR0_c21 <= exnR0_c20;
               D_c21 <= D_c20;
               betaw19_c21 <= betaw19_c20;
               q19_c21 <= q19_c20;
               absq19D_c21 <= absq19D_c20;
               qP28_c21 <= qP28_c20;
               qM28_c21 <= qM28_c20;
               qP27_c21 <= qP27_c20;
               qM27_c21 <= qM27_c20;
               qP26_c21 <= qP26_c20;
               qM26_c21 <= qM26_c20;
               qP25_c21 <= qP25_c20;
               qM25_c21 <= qM25_c20;
               qP24_c21 <= qP24_c20;
               qM24_c21 <= qM24_c20;
               qP23_c21 <= qP23_c20;
               qM23_c21 <= qM23_c20;
               qP22_c21 <= qP22_c20;
               qM22_c21 <= qM22_c20;
               qP21_c21 <= qP21_c20;
               qM21_c21 <= qM21_c20;
               qP20_c21 <= qP20_c20;
               qM20_c21 <= qM20_c20;
               qP19_c21 <= qP19_c20;
               qM19_c21 <= qM19_c20;
            end if;
            if ce_22 = '1' then
               expR0_c22 <= expR0_c21;
               sR_c22 <= sR_c21;
               exnR0_c22 <= exnR0_c21;
               D_c22 <= D_c21;
               betaw18_c22 <= betaw18_c21;
               q18_copy15_c22 <= q18_copy15_c21;
               qP28_c22 <= qP28_c21;
               qM28_c22 <= qM28_c21;
               qP27_c22 <= qP27_c21;
               qM27_c22 <= qM27_c21;
               qP26_c22 <= qP26_c21;
               qM26_c22 <= qM26_c21;
               qP25_c22 <= qP25_c21;
               qM25_c22 <= qM25_c21;
               qP24_c22 <= qP24_c21;
               qM24_c22 <= qM24_c21;
               qP23_c22 <= qP23_c21;
               qM23_c22 <= qM23_c21;
               qP22_c22 <= qP22_c21;
               qM22_c22 <= qM22_c21;
               qP21_c22 <= qP21_c21;
               qM21_c22 <= qM21_c21;
               qP20_c22 <= qP20_c21;
               qM20_c22 <= qM20_c21;
               qP19_c22 <= qP19_c21;
               qM19_c22 <= qM19_c21;
            end if;
            if ce_23 = '1' then
               expR0_c23 <= expR0_c22;
               sR_c23 <= sR_c22;
               exnR0_c23 <= exnR0_c22;
               D_c23 <= D_c22;
               betaw18_c23 <= betaw18_c22;
               q18_c23 <= q18_c22;
               absq18D_c23 <= absq18D_c22;
               qP28_c23 <= qP28_c22;
               qM28_c23 <= qM28_c22;
               qP27_c23 <= qP27_c22;
               qM27_c23 <= qM27_c22;
               qP26_c23 <= qP26_c22;
               qM26_c23 <= qM26_c22;
               qP25_c23 <= qP25_c22;
               qM25_c23 <= qM25_c22;
               qP24_c23 <= qP24_c22;
               qM24_c23 <= qM24_c22;
               qP23_c23 <= qP23_c22;
               qM23_c23 <= qM23_c22;
               qP22_c23 <= qP22_c22;
               qM22_c23 <= qM22_c22;
               qP21_c23 <= qP21_c22;
               qM21_c23 <= qM21_c22;
               qP20_c23 <= qP20_c22;
               qM20_c23 <= qM20_c22;
               qP19_c23 <= qP19_c22;
               qM19_c23 <= qM19_c22;
               qP18_c23 <= qP18_c22;
               qM18_c23 <= qM18_c22;
            end if;
            if ce_24 = '1' then
               expR0_c24 <= expR0_c23;
               sR_c24 <= sR_c23;
               exnR0_c24 <= exnR0_c23;
               D_c24 <= D_c23;
               betaw17_c24 <= betaw17_c23;
               q17_copy16_c24 <= q17_copy16_c23;
               qP28_c24 <= qP28_c23;
               qM28_c24 <= qM28_c23;
               qP27_c24 <= qP27_c23;
               qM27_c24 <= qM27_c23;
               qP26_c24 <= qP26_c23;
               qM26_c24 <= qM26_c23;
               qP25_c24 <= qP25_c23;
               qM25_c24 <= qM25_c23;
               qP24_c24 <= qP24_c23;
               qM24_c24 <= qM24_c23;
               qP23_c24 <= qP23_c23;
               qM23_c24 <= qM23_c23;
               qP22_c24 <= qP22_c23;
               qM22_c24 <= qM22_c23;
               qP21_c24 <= qP21_c23;
               qM21_c24 <= qM21_c23;
               qP20_c24 <= qP20_c23;
               qM20_c24 <= qM20_c23;
               qP19_c24 <= qP19_c23;
               qM19_c24 <= qM19_c23;
               qP18_c24 <= qP18_c23;
               qM18_c24 <= qM18_c23;
            end if;
            if ce_25 = '1' then
               expR0_c25 <= expR0_c24;
               sR_c25 <= sR_c24;
               exnR0_c25 <= exnR0_c24;
               D_c25 <= D_c24;
               betaw17_c25 <= betaw17_c24;
               q17_c25 <= q17_c24;
               absq17D_c25 <= absq17D_c24;
               qP28_c25 <= qP28_c24;
               qM28_c25 <= qM28_c24;
               qP27_c25 <= qP27_c24;
               qM27_c25 <= qM27_c24;
               qP26_c25 <= qP26_c24;
               qM26_c25 <= qM26_c24;
               qP25_c25 <= qP25_c24;
               qM25_c25 <= qM25_c24;
               qP24_c25 <= qP24_c24;
               qM24_c25 <= qM24_c24;
               qP23_c25 <= qP23_c24;
               qM23_c25 <= qM23_c24;
               qP22_c25 <= qP22_c24;
               qM22_c25 <= qM22_c24;
               qP21_c25 <= qP21_c24;
               qM21_c25 <= qM21_c24;
               qP20_c25 <= qP20_c24;
               qM20_c25 <= qM20_c24;
               qP19_c25 <= qP19_c24;
               qM19_c25 <= qM19_c24;
               qP18_c25 <= qP18_c24;
               qM18_c25 <= qM18_c24;
               qP17_c25 <= qP17_c24;
               qM17_c25 <= qM17_c24;
            end if;
            if ce_26 = '1' then
               expR0_c26 <= expR0_c25;
               sR_c26 <= sR_c25;
               exnR0_c26 <= exnR0_c25;
               D_c26 <= D_c25;
               betaw16_c26 <= betaw16_c25;
               q16_copy17_c26 <= q16_copy17_c25;
               qP28_c26 <= qP28_c25;
               qM28_c26 <= qM28_c25;
               qP27_c26 <= qP27_c25;
               qM27_c26 <= qM27_c25;
               qP26_c26 <= qP26_c25;
               qM26_c26 <= qM26_c25;
               qP25_c26 <= qP25_c25;
               qM25_c26 <= qM25_c25;
               qP24_c26 <= qP24_c25;
               qM24_c26 <= qM24_c25;
               qP23_c26 <= qP23_c25;
               qM23_c26 <= qM23_c25;
               qP22_c26 <= qP22_c25;
               qM22_c26 <= qM22_c25;
               qP21_c26 <= qP21_c25;
               qM21_c26 <= qM21_c25;
               qP20_c26 <= qP20_c25;
               qM20_c26 <= qM20_c25;
               qP19_c26 <= qP19_c25;
               qM19_c26 <= qM19_c25;
               qP18_c26 <= qP18_c25;
               qM18_c26 <= qM18_c25;
               qP17_c26 <= qP17_c25;
               qM17_c26 <= qM17_c25;
            end if;
            if ce_27 = '1' then
               expR0_c27 <= expR0_c26;
               sR_c27 <= sR_c26;
               exnR0_c27 <= exnR0_c26;
               D_c27 <= D_c26;
               betaw16_c27 <= betaw16_c26;
               q16_c27 <= q16_c26;
               absq16D_c27 <= absq16D_c26;
               qP28_c27 <= qP28_c26;
               qM28_c27 <= qM28_c26;
               qP27_c27 <= qP27_c26;
               qM27_c27 <= qM27_c26;
               qP26_c27 <= qP26_c26;
               qM26_c27 <= qM26_c26;
               qP25_c27 <= qP25_c26;
               qM25_c27 <= qM25_c26;
               qP24_c27 <= qP24_c26;
               qM24_c27 <= qM24_c26;
               qP23_c27 <= qP23_c26;
               qM23_c27 <= qM23_c26;
               qP22_c27 <= qP22_c26;
               qM22_c27 <= qM22_c26;
               qP21_c27 <= qP21_c26;
               qM21_c27 <= qM21_c26;
               qP20_c27 <= qP20_c26;
               qM20_c27 <= qM20_c26;
               qP19_c27 <= qP19_c26;
               qM19_c27 <= qM19_c26;
               qP18_c27 <= qP18_c26;
               qM18_c27 <= qM18_c26;
               qP17_c27 <= qP17_c26;
               qM17_c27 <= qM17_c26;
               qP16_c27 <= qP16_c26;
               qM16_c27 <= qM16_c26;
            end if;
            if ce_28 = '1' then
               expR0_c28 <= expR0_c27;
               sR_c28 <= sR_c27;
               exnR0_c28 <= exnR0_c27;
               D_c28 <= D_c27;
               betaw15_c28 <= betaw15_c27;
               q15_copy18_c28 <= q15_copy18_c27;
               qP28_c28 <= qP28_c27;
               qM28_c28 <= qM28_c27;
               qP27_c28 <= qP27_c27;
               qM27_c28 <= qM27_c27;
               qP26_c28 <= qP26_c27;
               qM26_c28 <= qM26_c27;
               qP25_c28 <= qP25_c27;
               qM25_c28 <= qM25_c27;
               qP24_c28 <= qP24_c27;
               qM24_c28 <= qM24_c27;
               qP23_c28 <= qP23_c27;
               qM23_c28 <= qM23_c27;
               qP22_c28 <= qP22_c27;
               qM22_c28 <= qM22_c27;
               qP21_c28 <= qP21_c27;
               qM21_c28 <= qM21_c27;
               qP20_c28 <= qP20_c27;
               qM20_c28 <= qM20_c27;
               qP19_c28 <= qP19_c27;
               qM19_c28 <= qM19_c27;
               qP18_c28 <= qP18_c27;
               qM18_c28 <= qM18_c27;
               qP17_c28 <= qP17_c27;
               qM17_c28 <= qM17_c27;
               qP16_c28 <= qP16_c27;
               qM16_c28 <= qM16_c27;
            end if;
            if ce_29 = '1' then
               expR0_c29 <= expR0_c28;
               sR_c29 <= sR_c28;
               exnR0_c29 <= exnR0_c28;
               D_c29 <= D_c28;
               betaw15_c29 <= betaw15_c28;
               q15_c29 <= q15_c28;
               absq15D_c29 <= absq15D_c28;
               qP28_c29 <= qP28_c28;
               qM28_c29 <= qM28_c28;
               qP27_c29 <= qP27_c28;
               qM27_c29 <= qM27_c28;
               qP26_c29 <= qP26_c28;
               qM26_c29 <= qM26_c28;
               qP25_c29 <= qP25_c28;
               qM25_c29 <= qM25_c28;
               qP24_c29 <= qP24_c28;
               qM24_c29 <= qM24_c28;
               qP23_c29 <= qP23_c28;
               qM23_c29 <= qM23_c28;
               qP22_c29 <= qP22_c28;
               qM22_c29 <= qM22_c28;
               qP21_c29 <= qP21_c28;
               qM21_c29 <= qM21_c28;
               qP20_c29 <= qP20_c28;
               qM20_c29 <= qM20_c28;
               qP19_c29 <= qP19_c28;
               qM19_c29 <= qM19_c28;
               qP18_c29 <= qP18_c28;
               qM18_c29 <= qM18_c28;
               qP17_c29 <= qP17_c28;
               qM17_c29 <= qM17_c28;
               qP16_c29 <= qP16_c28;
               qM16_c29 <= qM16_c28;
               qP15_c29 <= qP15_c28;
               qM15_c29 <= qM15_c28;
            end if;
            if ce_30 = '1' then
               expR0_c30 <= expR0_c29;
               sR_c30 <= sR_c29;
               exnR0_c30 <= exnR0_c29;
               D_c30 <= D_c29;
               betaw15_c30 <= betaw15_c29;
               q15_c30 <= q15_c29;
               absq15D_c30 <= absq15D_c29;
               qP28_c30 <= qP28_c29;
               qM28_c30 <= qM28_c29;
               qP27_c30 <= qP27_c29;
               qM27_c30 <= qM27_c29;
               qP26_c30 <= qP26_c29;
               qM26_c30 <= qM26_c29;
               qP25_c30 <= qP25_c29;
               qM25_c30 <= qM25_c29;
               qP24_c30 <= qP24_c29;
               qM24_c30 <= qM24_c29;
               qP23_c30 <= qP23_c29;
               qM23_c30 <= qM23_c29;
               qP22_c30 <= qP22_c29;
               qM22_c30 <= qM22_c29;
               qP21_c30 <= qP21_c29;
               qM21_c30 <= qM21_c29;
               qP20_c30 <= qP20_c29;
               qM20_c30 <= qM20_c29;
               qP19_c30 <= qP19_c29;
               qM19_c30 <= qM19_c29;
               qP18_c30 <= qP18_c29;
               qM18_c30 <= qM18_c29;
               qP17_c30 <= qP17_c29;
               qM17_c30 <= qM17_c29;
               qP16_c30 <= qP16_c29;
               qM16_c30 <= qM16_c29;
               qP15_c30 <= qP15_c29;
               qM15_c30 <= qM15_c29;
            end if;
            if ce_31 = '1' then
               expR0_c31 <= expR0_c30;
               sR_c31 <= sR_c30;
               exnR0_c31 <= exnR0_c30;
               D_c31 <= D_c30;
               betaw14_c31 <= betaw14_c30;
               q14_c31 <= q14_c30;
               absq14D_c31 <= absq14D_c30;
               qP28_c31 <= qP28_c30;
               qM28_c31 <= qM28_c30;
               qP27_c31 <= qP27_c30;
               qM27_c31 <= qM27_c30;
               qP26_c31 <= qP26_c30;
               qM26_c31 <= qM26_c30;
               qP25_c31 <= qP25_c30;
               qM25_c31 <= qM25_c30;
               qP24_c31 <= qP24_c30;
               qM24_c31 <= qM24_c30;
               qP23_c31 <= qP23_c30;
               qM23_c31 <= qM23_c30;
               qP22_c31 <= qP22_c30;
               qM22_c31 <= qM22_c30;
               qP21_c31 <= qP21_c30;
               qM21_c31 <= qM21_c30;
               qP20_c31 <= qP20_c30;
               qM20_c31 <= qM20_c30;
               qP19_c31 <= qP19_c30;
               qM19_c31 <= qM19_c30;
               qP18_c31 <= qP18_c30;
               qM18_c31 <= qM18_c30;
               qP17_c31 <= qP17_c30;
               qM17_c31 <= qM17_c30;
               qP16_c31 <= qP16_c30;
               qM16_c31 <= qM16_c30;
               qP15_c31 <= qP15_c30;
               qM15_c31 <= qM15_c30;
               qP14_c31 <= qP14_c30;
               qM14_c31 <= qM14_c30;
            end if;
            if ce_32 = '1' then
               expR0_c32 <= expR0_c31;
               sR_c32 <= sR_c31;
               exnR0_c32 <= exnR0_c31;
               D_c32 <= D_c31;
               betaw14_c32 <= betaw14_c31;
               q14_c32 <= q14_c31;
               absq14D_c32 <= absq14D_c31;
               qP28_c32 <= qP28_c31;
               qM28_c32 <= qM28_c31;
               qP27_c32 <= qP27_c31;
               qM27_c32 <= qM27_c31;
               qP26_c32 <= qP26_c31;
               qM26_c32 <= qM26_c31;
               qP25_c32 <= qP25_c31;
               qM25_c32 <= qM25_c31;
               qP24_c32 <= qP24_c31;
               qM24_c32 <= qM24_c31;
               qP23_c32 <= qP23_c31;
               qM23_c32 <= qM23_c31;
               qP22_c32 <= qP22_c31;
               qM22_c32 <= qM22_c31;
               qP21_c32 <= qP21_c31;
               qM21_c32 <= qM21_c31;
               qP20_c32 <= qP20_c31;
               qM20_c32 <= qM20_c31;
               qP19_c32 <= qP19_c31;
               qM19_c32 <= qM19_c31;
               qP18_c32 <= qP18_c31;
               qM18_c32 <= qM18_c31;
               qP17_c32 <= qP17_c31;
               qM17_c32 <= qM17_c31;
               qP16_c32 <= qP16_c31;
               qM16_c32 <= qM16_c31;
               qP15_c32 <= qP15_c31;
               qM15_c32 <= qM15_c31;
               qP14_c32 <= qP14_c31;
               qM14_c32 <= qM14_c31;
            end if;
            if ce_33 = '1' then
               expR0_c33 <= expR0_c32;
               sR_c33 <= sR_c32;
               exnR0_c33 <= exnR0_c32;
               D_c33 <= D_c32;
               betaw13_c33 <= betaw13_c32;
               q13_c33 <= q13_c32;
               absq13D_c33 <= absq13D_c32;
               qP28_c33 <= qP28_c32;
               qM28_c33 <= qM28_c32;
               qP27_c33 <= qP27_c32;
               qM27_c33 <= qM27_c32;
               qP26_c33 <= qP26_c32;
               qM26_c33 <= qM26_c32;
               qP25_c33 <= qP25_c32;
               qM25_c33 <= qM25_c32;
               qP24_c33 <= qP24_c32;
               qM24_c33 <= qM24_c32;
               qP23_c33 <= qP23_c32;
               qM23_c33 <= qM23_c32;
               qP22_c33 <= qP22_c32;
               qM22_c33 <= qM22_c32;
               qP21_c33 <= qP21_c32;
               qM21_c33 <= qM21_c32;
               qP20_c33 <= qP20_c32;
               qM20_c33 <= qM20_c32;
               qP19_c33 <= qP19_c32;
               qM19_c33 <= qM19_c32;
               qP18_c33 <= qP18_c32;
               qM18_c33 <= qM18_c32;
               qP17_c33 <= qP17_c32;
               qM17_c33 <= qM17_c32;
               qP16_c33 <= qP16_c32;
               qM16_c33 <= qM16_c32;
               qP15_c33 <= qP15_c32;
               qM15_c33 <= qM15_c32;
               qP14_c33 <= qP14_c32;
               qM14_c33 <= qM14_c32;
               qP13_c33 <= qP13_c32;
               qM13_c33 <= qM13_c32;
            end if;
            if ce_34 = '1' then
               expR0_c34 <= expR0_c33;
               sR_c34 <= sR_c33;
               exnR0_c34 <= exnR0_c33;
               D_c34 <= D_c33;
               betaw13_c34 <= betaw13_c33;
               q13_c34 <= q13_c33;
               absq13D_c34 <= absq13D_c33;
               qP28_c34 <= qP28_c33;
               qM28_c34 <= qM28_c33;
               qP27_c34 <= qP27_c33;
               qM27_c34 <= qM27_c33;
               qP26_c34 <= qP26_c33;
               qM26_c34 <= qM26_c33;
               qP25_c34 <= qP25_c33;
               qM25_c34 <= qM25_c33;
               qP24_c34 <= qP24_c33;
               qM24_c34 <= qM24_c33;
               qP23_c34 <= qP23_c33;
               qM23_c34 <= qM23_c33;
               qP22_c34 <= qP22_c33;
               qM22_c34 <= qM22_c33;
               qP21_c34 <= qP21_c33;
               qM21_c34 <= qM21_c33;
               qP20_c34 <= qP20_c33;
               qM20_c34 <= qM20_c33;
               qP19_c34 <= qP19_c33;
               qM19_c34 <= qM19_c33;
               qP18_c34 <= qP18_c33;
               qM18_c34 <= qM18_c33;
               qP17_c34 <= qP17_c33;
               qM17_c34 <= qM17_c33;
               qP16_c34 <= qP16_c33;
               qM16_c34 <= qM16_c33;
               qP15_c34 <= qP15_c33;
               qM15_c34 <= qM15_c33;
               qP14_c34 <= qP14_c33;
               qM14_c34 <= qM14_c33;
               qP13_c34 <= qP13_c33;
               qM13_c34 <= qM13_c33;
            end if;
            if ce_35 = '1' then
               expR0_c35 <= expR0_c34;
               sR_c35 <= sR_c34;
               exnR0_c35 <= exnR0_c34;
               D_c35 <= D_c34;
               betaw12_c35 <= betaw12_c34;
               q12_c35 <= q12_c34;
               absq12D_c35 <= absq12D_c34;
               qP28_c35 <= qP28_c34;
               qM28_c35 <= qM28_c34;
               qP27_c35 <= qP27_c34;
               qM27_c35 <= qM27_c34;
               qP26_c35 <= qP26_c34;
               qM26_c35 <= qM26_c34;
               qP25_c35 <= qP25_c34;
               qM25_c35 <= qM25_c34;
               qP24_c35 <= qP24_c34;
               qM24_c35 <= qM24_c34;
               qP23_c35 <= qP23_c34;
               qM23_c35 <= qM23_c34;
               qP22_c35 <= qP22_c34;
               qM22_c35 <= qM22_c34;
               qP21_c35 <= qP21_c34;
               qM21_c35 <= qM21_c34;
               qP20_c35 <= qP20_c34;
               qM20_c35 <= qM20_c34;
               qP19_c35 <= qP19_c34;
               qM19_c35 <= qM19_c34;
               qP18_c35 <= qP18_c34;
               qM18_c35 <= qM18_c34;
               qP17_c35 <= qP17_c34;
               qM17_c35 <= qM17_c34;
               qP16_c35 <= qP16_c34;
               qM16_c35 <= qM16_c34;
               qP15_c35 <= qP15_c34;
               qM15_c35 <= qM15_c34;
               qP14_c35 <= qP14_c34;
               qM14_c35 <= qM14_c34;
               qP13_c35 <= qP13_c34;
               qM13_c35 <= qM13_c34;
               qP12_c35 <= qP12_c34;
               qM12_c35 <= qM12_c34;
            end if;
            if ce_36 = '1' then
               expR0_c36 <= expR0_c35;
               sR_c36 <= sR_c35;
               exnR0_c36 <= exnR0_c35;
               D_c36 <= D_c35;
               betaw12_c36 <= betaw12_c35;
               q12_c36 <= q12_c35;
               absq12D_c36 <= absq12D_c35;
               qP28_c36 <= qP28_c35;
               qM28_c36 <= qM28_c35;
               qP27_c36 <= qP27_c35;
               qM27_c36 <= qM27_c35;
               qP26_c36 <= qP26_c35;
               qM26_c36 <= qM26_c35;
               qP25_c36 <= qP25_c35;
               qM25_c36 <= qM25_c35;
               qP24_c36 <= qP24_c35;
               qM24_c36 <= qM24_c35;
               qP23_c36 <= qP23_c35;
               qM23_c36 <= qM23_c35;
               qP22_c36 <= qP22_c35;
               qM22_c36 <= qM22_c35;
               qP21_c36 <= qP21_c35;
               qM21_c36 <= qM21_c35;
               qP20_c36 <= qP20_c35;
               qM20_c36 <= qM20_c35;
               qP19_c36 <= qP19_c35;
               qM19_c36 <= qM19_c35;
               qP18_c36 <= qP18_c35;
               qM18_c36 <= qM18_c35;
               qP17_c36 <= qP17_c35;
               qM17_c36 <= qM17_c35;
               qP16_c36 <= qP16_c35;
               qM16_c36 <= qM16_c35;
               qP15_c36 <= qP15_c35;
               qM15_c36 <= qM15_c35;
               qP14_c36 <= qP14_c35;
               qM14_c36 <= qM14_c35;
               qP13_c36 <= qP13_c35;
               qM13_c36 <= qM13_c35;
               qP12_c36 <= qP12_c35;
               qM12_c36 <= qM12_c35;
            end if;
            if ce_37 = '1' then
               expR0_c37 <= expR0_c36;
               sR_c37 <= sR_c36;
               exnR0_c37 <= exnR0_c36;
               D_c37 <= D_c36;
               betaw11_c37 <= betaw11_c36;
               q11_copy22_c37 <= q11_copy22_c36;
               qP28_c37 <= qP28_c36;
               qM28_c37 <= qM28_c36;
               qP27_c37 <= qP27_c36;
               qM27_c37 <= qM27_c36;
               qP26_c37 <= qP26_c36;
               qM26_c37 <= qM26_c36;
               qP25_c37 <= qP25_c36;
               qM25_c37 <= qM25_c36;
               qP24_c37 <= qP24_c36;
               qM24_c37 <= qM24_c36;
               qP23_c37 <= qP23_c36;
               qM23_c37 <= qM23_c36;
               qP22_c37 <= qP22_c36;
               qM22_c37 <= qM22_c36;
               qP21_c37 <= qP21_c36;
               qM21_c37 <= qM21_c36;
               qP20_c37 <= qP20_c36;
               qM20_c37 <= qM20_c36;
               qP19_c37 <= qP19_c36;
               qM19_c37 <= qM19_c36;
               qP18_c37 <= qP18_c36;
               qM18_c37 <= qM18_c36;
               qP17_c37 <= qP17_c36;
               qM17_c37 <= qM17_c36;
               qP16_c37 <= qP16_c36;
               qM16_c37 <= qM16_c36;
               qP15_c37 <= qP15_c36;
               qM15_c37 <= qM15_c36;
               qP14_c37 <= qP14_c36;
               qM14_c37 <= qM14_c36;
               qP13_c37 <= qP13_c36;
               qM13_c37 <= qM13_c36;
               qP12_c37 <= qP12_c36;
               qM12_c37 <= qM12_c36;
            end if;
            if ce_38 = '1' then
               expR0_c38 <= expR0_c37;
               sR_c38 <= sR_c37;
               exnR0_c38 <= exnR0_c37;
               D_c38 <= D_c37;
               betaw11_c38 <= betaw11_c37;
               q11_c38 <= q11_c37;
               absq11D_c38 <= absq11D_c37;
               qP28_c38 <= qP28_c37;
               qM28_c38 <= qM28_c37;
               qP27_c38 <= qP27_c37;
               qM27_c38 <= qM27_c37;
               qP26_c38 <= qP26_c37;
               qM26_c38 <= qM26_c37;
               qP25_c38 <= qP25_c37;
               qM25_c38 <= qM25_c37;
               qP24_c38 <= qP24_c37;
               qM24_c38 <= qM24_c37;
               qP23_c38 <= qP23_c37;
               qM23_c38 <= qM23_c37;
               qP22_c38 <= qP22_c37;
               qM22_c38 <= qM22_c37;
               qP21_c38 <= qP21_c37;
               qM21_c38 <= qM21_c37;
               qP20_c38 <= qP20_c37;
               qM20_c38 <= qM20_c37;
               qP19_c38 <= qP19_c37;
               qM19_c38 <= qM19_c37;
               qP18_c38 <= qP18_c37;
               qM18_c38 <= qM18_c37;
               qP17_c38 <= qP17_c37;
               qM17_c38 <= qM17_c37;
               qP16_c38 <= qP16_c37;
               qM16_c38 <= qM16_c37;
               qP15_c38 <= qP15_c37;
               qM15_c38 <= qM15_c37;
               qP14_c38 <= qP14_c37;
               qM14_c38 <= qM14_c37;
               qP13_c38 <= qP13_c37;
               qM13_c38 <= qM13_c37;
               qP12_c38 <= qP12_c37;
               qM12_c38 <= qM12_c37;
               qP11_c38 <= qP11_c37;
               qM11_c38 <= qM11_c37;
            end if;
            if ce_39 = '1' then
               expR0_c39 <= expR0_c38;
               sR_c39 <= sR_c38;
               exnR0_c39 <= exnR0_c38;
               D_c39 <= D_c38;
               betaw10_c39 <= betaw10_c38;
               q10_copy23_c39 <= q10_copy23_c38;
               qP28_c39 <= qP28_c38;
               qM28_c39 <= qM28_c38;
               qP27_c39 <= qP27_c38;
               qM27_c39 <= qM27_c38;
               qP26_c39 <= qP26_c38;
               qM26_c39 <= qM26_c38;
               qP25_c39 <= qP25_c38;
               qM25_c39 <= qM25_c38;
               qP24_c39 <= qP24_c38;
               qM24_c39 <= qM24_c38;
               qP23_c39 <= qP23_c38;
               qM23_c39 <= qM23_c38;
               qP22_c39 <= qP22_c38;
               qM22_c39 <= qM22_c38;
               qP21_c39 <= qP21_c38;
               qM21_c39 <= qM21_c38;
               qP20_c39 <= qP20_c38;
               qM20_c39 <= qM20_c38;
               qP19_c39 <= qP19_c38;
               qM19_c39 <= qM19_c38;
               qP18_c39 <= qP18_c38;
               qM18_c39 <= qM18_c38;
               qP17_c39 <= qP17_c38;
               qM17_c39 <= qM17_c38;
               qP16_c39 <= qP16_c38;
               qM16_c39 <= qM16_c38;
               qP15_c39 <= qP15_c38;
               qM15_c39 <= qM15_c38;
               qP14_c39 <= qP14_c38;
               qM14_c39 <= qM14_c38;
               qP13_c39 <= qP13_c38;
               qM13_c39 <= qM13_c38;
               qP12_c39 <= qP12_c38;
               qM12_c39 <= qM12_c38;
               qP11_c39 <= qP11_c38;
               qM11_c39 <= qM11_c38;
            end if;
            if ce_40 = '1' then
               expR0_c40 <= expR0_c39;
               sR_c40 <= sR_c39;
               exnR0_c40 <= exnR0_c39;
               D_c40 <= D_c39;
               betaw10_c40 <= betaw10_c39;
               q10_c40 <= q10_c39;
               absq10D_c40 <= absq10D_c39;
               qP28_c40 <= qP28_c39;
               qM28_c40 <= qM28_c39;
               qP27_c40 <= qP27_c39;
               qM27_c40 <= qM27_c39;
               qP26_c40 <= qP26_c39;
               qM26_c40 <= qM26_c39;
               qP25_c40 <= qP25_c39;
               qM25_c40 <= qM25_c39;
               qP24_c40 <= qP24_c39;
               qM24_c40 <= qM24_c39;
               qP23_c40 <= qP23_c39;
               qM23_c40 <= qM23_c39;
               qP22_c40 <= qP22_c39;
               qM22_c40 <= qM22_c39;
               qP21_c40 <= qP21_c39;
               qM21_c40 <= qM21_c39;
               qP20_c40 <= qP20_c39;
               qM20_c40 <= qM20_c39;
               qP19_c40 <= qP19_c39;
               qM19_c40 <= qM19_c39;
               qP18_c40 <= qP18_c39;
               qM18_c40 <= qM18_c39;
               qP17_c40 <= qP17_c39;
               qM17_c40 <= qM17_c39;
               qP16_c40 <= qP16_c39;
               qM16_c40 <= qM16_c39;
               qP15_c40 <= qP15_c39;
               qM15_c40 <= qM15_c39;
               qP14_c40 <= qP14_c39;
               qM14_c40 <= qM14_c39;
               qP13_c40 <= qP13_c39;
               qM13_c40 <= qM13_c39;
               qP12_c40 <= qP12_c39;
               qM12_c40 <= qM12_c39;
               qP11_c40 <= qP11_c39;
               qM11_c40 <= qM11_c39;
               qP10_c40 <= qP10_c39;
               qM10_c40 <= qM10_c39;
            end if;
            if ce_41 = '1' then
               expR0_c41 <= expR0_c40;
               sR_c41 <= sR_c40;
               exnR0_c41 <= exnR0_c40;
               D_c41 <= D_c40;
               betaw9_c41 <= betaw9_c40;
               q9_copy24_c41 <= q9_copy24_c40;
               qP28_c41 <= qP28_c40;
               qM28_c41 <= qM28_c40;
               qP27_c41 <= qP27_c40;
               qM27_c41 <= qM27_c40;
               qP26_c41 <= qP26_c40;
               qM26_c41 <= qM26_c40;
               qP25_c41 <= qP25_c40;
               qM25_c41 <= qM25_c40;
               qP24_c41 <= qP24_c40;
               qM24_c41 <= qM24_c40;
               qP23_c41 <= qP23_c40;
               qM23_c41 <= qM23_c40;
               qP22_c41 <= qP22_c40;
               qM22_c41 <= qM22_c40;
               qP21_c41 <= qP21_c40;
               qM21_c41 <= qM21_c40;
               qP20_c41 <= qP20_c40;
               qM20_c41 <= qM20_c40;
               qP19_c41 <= qP19_c40;
               qM19_c41 <= qM19_c40;
               qP18_c41 <= qP18_c40;
               qM18_c41 <= qM18_c40;
               qP17_c41 <= qP17_c40;
               qM17_c41 <= qM17_c40;
               qP16_c41 <= qP16_c40;
               qM16_c41 <= qM16_c40;
               qP15_c41 <= qP15_c40;
               qM15_c41 <= qM15_c40;
               qP14_c41 <= qP14_c40;
               qM14_c41 <= qM14_c40;
               qP13_c41 <= qP13_c40;
               qM13_c41 <= qM13_c40;
               qP12_c41 <= qP12_c40;
               qM12_c41 <= qM12_c40;
               qP11_c41 <= qP11_c40;
               qM11_c41 <= qM11_c40;
               qP10_c41 <= qP10_c40;
               qM10_c41 <= qM10_c40;
            end if;
            if ce_42 = '1' then
               expR0_c42 <= expR0_c41;
               sR_c42 <= sR_c41;
               exnR0_c42 <= exnR0_c41;
               D_c42 <= D_c41;
               betaw9_c42 <= betaw9_c41;
               q9_c42 <= q9_c41;
               absq9D_c42 <= absq9D_c41;
               qP28_c42 <= qP28_c41;
               qM28_c42 <= qM28_c41;
               qP27_c42 <= qP27_c41;
               qM27_c42 <= qM27_c41;
               qP26_c42 <= qP26_c41;
               qM26_c42 <= qM26_c41;
               qP25_c42 <= qP25_c41;
               qM25_c42 <= qM25_c41;
               qP24_c42 <= qP24_c41;
               qM24_c42 <= qM24_c41;
               qP23_c42 <= qP23_c41;
               qM23_c42 <= qM23_c41;
               qP22_c42 <= qP22_c41;
               qM22_c42 <= qM22_c41;
               qP21_c42 <= qP21_c41;
               qM21_c42 <= qM21_c41;
               qP20_c42 <= qP20_c41;
               qM20_c42 <= qM20_c41;
               qP19_c42 <= qP19_c41;
               qM19_c42 <= qM19_c41;
               qP18_c42 <= qP18_c41;
               qM18_c42 <= qM18_c41;
               qP17_c42 <= qP17_c41;
               qM17_c42 <= qM17_c41;
               qP16_c42 <= qP16_c41;
               qM16_c42 <= qM16_c41;
               qP15_c42 <= qP15_c41;
               qM15_c42 <= qM15_c41;
               qP14_c42 <= qP14_c41;
               qM14_c42 <= qM14_c41;
               qP13_c42 <= qP13_c41;
               qM13_c42 <= qM13_c41;
               qP12_c42 <= qP12_c41;
               qM12_c42 <= qM12_c41;
               qP11_c42 <= qP11_c41;
               qM11_c42 <= qM11_c41;
               qP10_c42 <= qP10_c41;
               qM10_c42 <= qM10_c41;
               qP9_c42 <= qP9_c41;
               qM9_c42 <= qM9_c41;
            end if;
            if ce_43 = '1' then
               expR0_c43 <= expR0_c42;
               sR_c43 <= sR_c42;
               exnR0_c43 <= exnR0_c42;
               D_c43 <= D_c42;
               betaw8_c43 <= betaw8_c42;
               q8_copy25_c43 <= q8_copy25_c42;
               qP28_c43 <= qP28_c42;
               qM28_c43 <= qM28_c42;
               qP27_c43 <= qP27_c42;
               qM27_c43 <= qM27_c42;
               qP26_c43 <= qP26_c42;
               qM26_c43 <= qM26_c42;
               qP25_c43 <= qP25_c42;
               qM25_c43 <= qM25_c42;
               qP24_c43 <= qP24_c42;
               qM24_c43 <= qM24_c42;
               qP23_c43 <= qP23_c42;
               qM23_c43 <= qM23_c42;
               qP22_c43 <= qP22_c42;
               qM22_c43 <= qM22_c42;
               qP21_c43 <= qP21_c42;
               qM21_c43 <= qM21_c42;
               qP20_c43 <= qP20_c42;
               qM20_c43 <= qM20_c42;
               qP19_c43 <= qP19_c42;
               qM19_c43 <= qM19_c42;
               qP18_c43 <= qP18_c42;
               qM18_c43 <= qM18_c42;
               qP17_c43 <= qP17_c42;
               qM17_c43 <= qM17_c42;
               qP16_c43 <= qP16_c42;
               qM16_c43 <= qM16_c42;
               qP15_c43 <= qP15_c42;
               qM15_c43 <= qM15_c42;
               qP14_c43 <= qP14_c42;
               qM14_c43 <= qM14_c42;
               qP13_c43 <= qP13_c42;
               qM13_c43 <= qM13_c42;
               qP12_c43 <= qP12_c42;
               qM12_c43 <= qM12_c42;
               qP11_c43 <= qP11_c42;
               qM11_c43 <= qM11_c42;
               qP10_c43 <= qP10_c42;
               qM10_c43 <= qM10_c42;
               qP9_c43 <= qP9_c42;
               qM9_c43 <= qM9_c42;
            end if;
            if ce_44 = '1' then
               expR0_c44 <= expR0_c43;
               sR_c44 <= sR_c43;
               exnR0_c44 <= exnR0_c43;
               D_c44 <= D_c43;
               betaw8_c44 <= betaw8_c43;
               q8_c44 <= q8_c43;
               absq8D_c44 <= absq8D_c43;
               qP28_c44 <= qP28_c43;
               qM28_c44 <= qM28_c43;
               qP27_c44 <= qP27_c43;
               qM27_c44 <= qM27_c43;
               qP26_c44 <= qP26_c43;
               qM26_c44 <= qM26_c43;
               qP25_c44 <= qP25_c43;
               qM25_c44 <= qM25_c43;
               qP24_c44 <= qP24_c43;
               qM24_c44 <= qM24_c43;
               qP23_c44 <= qP23_c43;
               qM23_c44 <= qM23_c43;
               qP22_c44 <= qP22_c43;
               qM22_c44 <= qM22_c43;
               qP21_c44 <= qP21_c43;
               qM21_c44 <= qM21_c43;
               qP20_c44 <= qP20_c43;
               qM20_c44 <= qM20_c43;
               qP19_c44 <= qP19_c43;
               qM19_c44 <= qM19_c43;
               qP18_c44 <= qP18_c43;
               qM18_c44 <= qM18_c43;
               qP17_c44 <= qP17_c43;
               qM17_c44 <= qM17_c43;
               qP16_c44 <= qP16_c43;
               qM16_c44 <= qM16_c43;
               qP15_c44 <= qP15_c43;
               qM15_c44 <= qM15_c43;
               qP14_c44 <= qP14_c43;
               qM14_c44 <= qM14_c43;
               qP13_c44 <= qP13_c43;
               qM13_c44 <= qM13_c43;
               qP12_c44 <= qP12_c43;
               qM12_c44 <= qM12_c43;
               qP11_c44 <= qP11_c43;
               qM11_c44 <= qM11_c43;
               qP10_c44 <= qP10_c43;
               qM10_c44 <= qM10_c43;
               qP9_c44 <= qP9_c43;
               qM9_c44 <= qM9_c43;
               qP8_c44 <= qP8_c43;
               qM8_c44 <= qM8_c43;
            end if;
            if ce_45 = '1' then
               expR0_c45 <= expR0_c44;
               sR_c45 <= sR_c44;
               exnR0_c45 <= exnR0_c44;
               D_c45 <= D_c44;
               betaw8_c45 <= betaw8_c44;
               q8_c45 <= q8_c44;
               absq8D_c45 <= absq8D_c44;
               qP28_c45 <= qP28_c44;
               qM28_c45 <= qM28_c44;
               qP27_c45 <= qP27_c44;
               qM27_c45 <= qM27_c44;
               qP26_c45 <= qP26_c44;
               qM26_c45 <= qM26_c44;
               qP25_c45 <= qP25_c44;
               qM25_c45 <= qM25_c44;
               qP24_c45 <= qP24_c44;
               qM24_c45 <= qM24_c44;
               qP23_c45 <= qP23_c44;
               qM23_c45 <= qM23_c44;
               qP22_c45 <= qP22_c44;
               qM22_c45 <= qM22_c44;
               qP21_c45 <= qP21_c44;
               qM21_c45 <= qM21_c44;
               qP20_c45 <= qP20_c44;
               qM20_c45 <= qM20_c44;
               qP19_c45 <= qP19_c44;
               qM19_c45 <= qM19_c44;
               qP18_c45 <= qP18_c44;
               qM18_c45 <= qM18_c44;
               qP17_c45 <= qP17_c44;
               qM17_c45 <= qM17_c44;
               qP16_c45 <= qP16_c44;
               qM16_c45 <= qM16_c44;
               qP15_c45 <= qP15_c44;
               qM15_c45 <= qM15_c44;
               qP14_c45 <= qP14_c44;
               qM14_c45 <= qM14_c44;
               qP13_c45 <= qP13_c44;
               qM13_c45 <= qM13_c44;
               qP12_c45 <= qP12_c44;
               qM12_c45 <= qM12_c44;
               qP11_c45 <= qP11_c44;
               qM11_c45 <= qM11_c44;
               qP10_c45 <= qP10_c44;
               qM10_c45 <= qM10_c44;
               qP9_c45 <= qP9_c44;
               qM9_c45 <= qM9_c44;
               qP8_c45 <= qP8_c44;
               qM8_c45 <= qM8_c44;
            end if;
            if ce_46 = '1' then
               expR0_c46 <= expR0_c45;
               sR_c46 <= sR_c45;
               exnR0_c46 <= exnR0_c45;
               D_c46 <= D_c45;
               betaw7_c46 <= betaw7_c45;
               q7_c46 <= q7_c45;
               absq7D_c46 <= absq7D_c45;
               qP28_c46 <= qP28_c45;
               qM28_c46 <= qM28_c45;
               qP27_c46 <= qP27_c45;
               qM27_c46 <= qM27_c45;
               qP26_c46 <= qP26_c45;
               qM26_c46 <= qM26_c45;
               qP25_c46 <= qP25_c45;
               qM25_c46 <= qM25_c45;
               qP24_c46 <= qP24_c45;
               qM24_c46 <= qM24_c45;
               qP23_c46 <= qP23_c45;
               qM23_c46 <= qM23_c45;
               qP22_c46 <= qP22_c45;
               qM22_c46 <= qM22_c45;
               qP21_c46 <= qP21_c45;
               qM21_c46 <= qM21_c45;
               qP20_c46 <= qP20_c45;
               qM20_c46 <= qM20_c45;
               qP19_c46 <= qP19_c45;
               qM19_c46 <= qM19_c45;
               qP18_c46 <= qP18_c45;
               qM18_c46 <= qM18_c45;
               qP17_c46 <= qP17_c45;
               qM17_c46 <= qM17_c45;
               qP16_c46 <= qP16_c45;
               qM16_c46 <= qM16_c45;
               qP15_c46 <= qP15_c45;
               qM15_c46 <= qM15_c45;
               qP14_c46 <= qP14_c45;
               qM14_c46 <= qM14_c45;
               qP13_c46 <= qP13_c45;
               qM13_c46 <= qM13_c45;
               qP12_c46 <= qP12_c45;
               qM12_c46 <= qM12_c45;
               qP11_c46 <= qP11_c45;
               qM11_c46 <= qM11_c45;
               qP10_c46 <= qP10_c45;
               qM10_c46 <= qM10_c45;
               qP9_c46 <= qP9_c45;
               qM9_c46 <= qM9_c45;
               qP8_c46 <= qP8_c45;
               qM8_c46 <= qM8_c45;
               qP7_c46 <= qP7_c45;
               qM7_c46 <= qM7_c45;
            end if;
            if ce_47 = '1' then
               expR0_c47 <= expR0_c46;
               sR_c47 <= sR_c46;
               exnR0_c47 <= exnR0_c46;
               D_c47 <= D_c46;
               betaw7_c47 <= betaw7_c46;
               q7_c47 <= q7_c46;
               absq7D_c47 <= absq7D_c46;
               qP28_c47 <= qP28_c46;
               qM28_c47 <= qM28_c46;
               qP27_c47 <= qP27_c46;
               qM27_c47 <= qM27_c46;
               qP26_c47 <= qP26_c46;
               qM26_c47 <= qM26_c46;
               qP25_c47 <= qP25_c46;
               qM25_c47 <= qM25_c46;
               qP24_c47 <= qP24_c46;
               qM24_c47 <= qM24_c46;
               qP23_c47 <= qP23_c46;
               qM23_c47 <= qM23_c46;
               qP22_c47 <= qP22_c46;
               qM22_c47 <= qM22_c46;
               qP21_c47 <= qP21_c46;
               qM21_c47 <= qM21_c46;
               qP20_c47 <= qP20_c46;
               qM20_c47 <= qM20_c46;
               qP19_c47 <= qP19_c46;
               qM19_c47 <= qM19_c46;
               qP18_c47 <= qP18_c46;
               qM18_c47 <= qM18_c46;
               qP17_c47 <= qP17_c46;
               qM17_c47 <= qM17_c46;
               qP16_c47 <= qP16_c46;
               qM16_c47 <= qM16_c46;
               qP15_c47 <= qP15_c46;
               qM15_c47 <= qM15_c46;
               qP14_c47 <= qP14_c46;
               qM14_c47 <= qM14_c46;
               qP13_c47 <= qP13_c46;
               qM13_c47 <= qM13_c46;
               qP12_c47 <= qP12_c46;
               qM12_c47 <= qM12_c46;
               qP11_c47 <= qP11_c46;
               qM11_c47 <= qM11_c46;
               qP10_c47 <= qP10_c46;
               qM10_c47 <= qM10_c46;
               qP9_c47 <= qP9_c46;
               qM9_c47 <= qM9_c46;
               qP8_c47 <= qP8_c46;
               qM8_c47 <= qM8_c46;
               qP7_c47 <= qP7_c46;
               qM7_c47 <= qM7_c46;
            end if;
            if ce_48 = '1' then
               expR0_c48 <= expR0_c47;
               sR_c48 <= sR_c47;
               exnR0_c48 <= exnR0_c47;
               D_c48 <= D_c47;
               betaw6_c48 <= betaw6_c47;
               q6_c48 <= q6_c47;
               absq6D_c48 <= absq6D_c47;
               qP28_c48 <= qP28_c47;
               qM28_c48 <= qM28_c47;
               qP27_c48 <= qP27_c47;
               qM27_c48 <= qM27_c47;
               qP26_c48 <= qP26_c47;
               qM26_c48 <= qM26_c47;
               qP25_c48 <= qP25_c47;
               qM25_c48 <= qM25_c47;
               qP24_c48 <= qP24_c47;
               qM24_c48 <= qM24_c47;
               qP23_c48 <= qP23_c47;
               qM23_c48 <= qM23_c47;
               qP22_c48 <= qP22_c47;
               qM22_c48 <= qM22_c47;
               qP21_c48 <= qP21_c47;
               qM21_c48 <= qM21_c47;
               qP20_c48 <= qP20_c47;
               qM20_c48 <= qM20_c47;
               qP19_c48 <= qP19_c47;
               qM19_c48 <= qM19_c47;
               qP18_c48 <= qP18_c47;
               qM18_c48 <= qM18_c47;
               qP17_c48 <= qP17_c47;
               qM17_c48 <= qM17_c47;
               qP16_c48 <= qP16_c47;
               qM16_c48 <= qM16_c47;
               qP15_c48 <= qP15_c47;
               qM15_c48 <= qM15_c47;
               qP14_c48 <= qP14_c47;
               qM14_c48 <= qM14_c47;
               qP13_c48 <= qP13_c47;
               qM13_c48 <= qM13_c47;
               qP12_c48 <= qP12_c47;
               qM12_c48 <= qM12_c47;
               qP11_c48 <= qP11_c47;
               qM11_c48 <= qM11_c47;
               qP10_c48 <= qP10_c47;
               qM10_c48 <= qM10_c47;
               qP9_c48 <= qP9_c47;
               qM9_c48 <= qM9_c47;
               qP8_c48 <= qP8_c47;
               qM8_c48 <= qM8_c47;
               qP7_c48 <= qP7_c47;
               qM7_c48 <= qM7_c47;
               qP6_c48 <= qP6_c47;
               qM6_c48 <= qM6_c47;
            end if;
            if ce_49 = '1' then
               expR0_c49 <= expR0_c48;
               sR_c49 <= sR_c48;
               exnR0_c49 <= exnR0_c48;
               D_c49 <= D_c48;
               betaw6_c49 <= betaw6_c48;
               q6_c49 <= q6_c48;
               absq6D_c49 <= absq6D_c48;
               qP28_c49 <= qP28_c48;
               qM28_c49 <= qM28_c48;
               qP27_c49 <= qP27_c48;
               qM27_c49 <= qM27_c48;
               qP26_c49 <= qP26_c48;
               qM26_c49 <= qM26_c48;
               qP25_c49 <= qP25_c48;
               qM25_c49 <= qM25_c48;
               qP24_c49 <= qP24_c48;
               qM24_c49 <= qM24_c48;
               qP23_c49 <= qP23_c48;
               qM23_c49 <= qM23_c48;
               qP22_c49 <= qP22_c48;
               qM22_c49 <= qM22_c48;
               qP21_c49 <= qP21_c48;
               qM21_c49 <= qM21_c48;
               qP20_c49 <= qP20_c48;
               qM20_c49 <= qM20_c48;
               qP19_c49 <= qP19_c48;
               qM19_c49 <= qM19_c48;
               qP18_c49 <= qP18_c48;
               qM18_c49 <= qM18_c48;
               qP17_c49 <= qP17_c48;
               qM17_c49 <= qM17_c48;
               qP16_c49 <= qP16_c48;
               qM16_c49 <= qM16_c48;
               qP15_c49 <= qP15_c48;
               qM15_c49 <= qM15_c48;
               qP14_c49 <= qP14_c48;
               qM14_c49 <= qM14_c48;
               qP13_c49 <= qP13_c48;
               qM13_c49 <= qM13_c48;
               qP12_c49 <= qP12_c48;
               qM12_c49 <= qM12_c48;
               qP11_c49 <= qP11_c48;
               qM11_c49 <= qM11_c48;
               qP10_c49 <= qP10_c48;
               qM10_c49 <= qM10_c48;
               qP9_c49 <= qP9_c48;
               qM9_c49 <= qM9_c48;
               qP8_c49 <= qP8_c48;
               qM8_c49 <= qM8_c48;
               qP7_c49 <= qP7_c48;
               qM7_c49 <= qM7_c48;
               qP6_c49 <= qP6_c48;
               qM6_c49 <= qM6_c48;
            end if;
            if ce_50 = '1' then
               expR0_c50 <= expR0_c49;
               sR_c50 <= sR_c49;
               exnR0_c50 <= exnR0_c49;
               D_c50 <= D_c49;
               betaw5_c50 <= betaw5_c49;
               q5_c50 <= q5_c49;
               absq5D_c50 <= absq5D_c49;
               qP28_c50 <= qP28_c49;
               qM28_c50 <= qM28_c49;
               qP27_c50 <= qP27_c49;
               qM27_c50 <= qM27_c49;
               qP26_c50 <= qP26_c49;
               qM26_c50 <= qM26_c49;
               qP25_c50 <= qP25_c49;
               qM25_c50 <= qM25_c49;
               qP24_c50 <= qP24_c49;
               qM24_c50 <= qM24_c49;
               qP23_c50 <= qP23_c49;
               qM23_c50 <= qM23_c49;
               qP22_c50 <= qP22_c49;
               qM22_c50 <= qM22_c49;
               qP21_c50 <= qP21_c49;
               qM21_c50 <= qM21_c49;
               qP20_c50 <= qP20_c49;
               qM20_c50 <= qM20_c49;
               qP19_c50 <= qP19_c49;
               qM19_c50 <= qM19_c49;
               qP18_c50 <= qP18_c49;
               qM18_c50 <= qM18_c49;
               qP17_c50 <= qP17_c49;
               qM17_c50 <= qM17_c49;
               qP16_c50 <= qP16_c49;
               qM16_c50 <= qM16_c49;
               qP15_c50 <= qP15_c49;
               qM15_c50 <= qM15_c49;
               qP14_c50 <= qP14_c49;
               qM14_c50 <= qM14_c49;
               qP13_c50 <= qP13_c49;
               qM13_c50 <= qM13_c49;
               qP12_c50 <= qP12_c49;
               qM12_c50 <= qM12_c49;
               qP11_c50 <= qP11_c49;
               qM11_c50 <= qM11_c49;
               qP10_c50 <= qP10_c49;
               qM10_c50 <= qM10_c49;
               qP9_c50 <= qP9_c49;
               qM9_c50 <= qM9_c49;
               qP8_c50 <= qP8_c49;
               qM8_c50 <= qM8_c49;
               qP7_c50 <= qP7_c49;
               qM7_c50 <= qM7_c49;
               qP6_c50 <= qP6_c49;
               qM6_c50 <= qM6_c49;
               qP5_c50 <= qP5_c49;
               qM5_c50 <= qM5_c49;
            end if;
            if ce_51 = '1' then
               expR0_c51 <= expR0_c50;
               sR_c51 <= sR_c50;
               exnR0_c51 <= exnR0_c50;
               D_c51 <= D_c50;
               betaw5_c51 <= betaw5_c50;
               q5_c51 <= q5_c50;
               absq5D_c51 <= absq5D_c50;
               qP28_c51 <= qP28_c50;
               qM28_c51 <= qM28_c50;
               qP27_c51 <= qP27_c50;
               qM27_c51 <= qM27_c50;
               qP26_c51 <= qP26_c50;
               qM26_c51 <= qM26_c50;
               qP25_c51 <= qP25_c50;
               qM25_c51 <= qM25_c50;
               qP24_c51 <= qP24_c50;
               qM24_c51 <= qM24_c50;
               qP23_c51 <= qP23_c50;
               qM23_c51 <= qM23_c50;
               qP22_c51 <= qP22_c50;
               qM22_c51 <= qM22_c50;
               qP21_c51 <= qP21_c50;
               qM21_c51 <= qM21_c50;
               qP20_c51 <= qP20_c50;
               qM20_c51 <= qM20_c50;
               qP19_c51 <= qP19_c50;
               qM19_c51 <= qM19_c50;
               qP18_c51 <= qP18_c50;
               qM18_c51 <= qM18_c50;
               qP17_c51 <= qP17_c50;
               qM17_c51 <= qM17_c50;
               qP16_c51 <= qP16_c50;
               qM16_c51 <= qM16_c50;
               qP15_c51 <= qP15_c50;
               qM15_c51 <= qM15_c50;
               qP14_c51 <= qP14_c50;
               qM14_c51 <= qM14_c50;
               qP13_c51 <= qP13_c50;
               qM13_c51 <= qM13_c50;
               qP12_c51 <= qP12_c50;
               qM12_c51 <= qM12_c50;
               qP11_c51 <= qP11_c50;
               qM11_c51 <= qM11_c50;
               qP10_c51 <= qP10_c50;
               qM10_c51 <= qM10_c50;
               qP9_c51 <= qP9_c50;
               qM9_c51 <= qM9_c50;
               qP8_c51 <= qP8_c50;
               qM8_c51 <= qM8_c50;
               qP7_c51 <= qP7_c50;
               qM7_c51 <= qM7_c50;
               qP6_c51 <= qP6_c50;
               qM6_c51 <= qM6_c50;
               qP5_c51 <= qP5_c50;
               qM5_c51 <= qM5_c50;
            end if;
            if ce_52 = '1' then
               expR0_c52 <= expR0_c51;
               sR_c52 <= sR_c51;
               exnR0_c52 <= exnR0_c51;
               D_c52 <= D_c51;
               betaw4_c52 <= betaw4_c51;
               q4_copy29_c52 <= q4_copy29_c51;
               qP28_c52 <= qP28_c51;
               qM28_c52 <= qM28_c51;
               qP27_c52 <= qP27_c51;
               qM27_c52 <= qM27_c51;
               qP26_c52 <= qP26_c51;
               qM26_c52 <= qM26_c51;
               qP25_c52 <= qP25_c51;
               qM25_c52 <= qM25_c51;
               qP24_c52 <= qP24_c51;
               qM24_c52 <= qM24_c51;
               qP23_c52 <= qP23_c51;
               qM23_c52 <= qM23_c51;
               qP22_c52 <= qP22_c51;
               qM22_c52 <= qM22_c51;
               qP21_c52 <= qP21_c51;
               qM21_c52 <= qM21_c51;
               qP20_c52 <= qP20_c51;
               qM20_c52 <= qM20_c51;
               qP19_c52 <= qP19_c51;
               qM19_c52 <= qM19_c51;
               qP18_c52 <= qP18_c51;
               qM18_c52 <= qM18_c51;
               qP17_c52 <= qP17_c51;
               qM17_c52 <= qM17_c51;
               qP16_c52 <= qP16_c51;
               qM16_c52 <= qM16_c51;
               qP15_c52 <= qP15_c51;
               qM15_c52 <= qM15_c51;
               qP14_c52 <= qP14_c51;
               qM14_c52 <= qM14_c51;
               qP13_c52 <= qP13_c51;
               qM13_c52 <= qM13_c51;
               qP12_c52 <= qP12_c51;
               qM12_c52 <= qM12_c51;
               qP11_c52 <= qP11_c51;
               qM11_c52 <= qM11_c51;
               qP10_c52 <= qP10_c51;
               qM10_c52 <= qM10_c51;
               qP9_c52 <= qP9_c51;
               qM9_c52 <= qM9_c51;
               qP8_c52 <= qP8_c51;
               qM8_c52 <= qM8_c51;
               qP7_c52 <= qP7_c51;
               qM7_c52 <= qM7_c51;
               qP6_c52 <= qP6_c51;
               qM6_c52 <= qM6_c51;
               qP5_c52 <= qP5_c51;
               qM5_c52 <= qM5_c51;
            end if;
            if ce_53 = '1' then
               expR0_c53 <= expR0_c52;
               sR_c53 <= sR_c52;
               exnR0_c53 <= exnR0_c52;
               D_c53 <= D_c52;
               betaw4_c53 <= betaw4_c52;
               q4_c53 <= q4_c52;
               absq4D_c53 <= absq4D_c52;
               qP28_c53 <= qP28_c52;
               qM28_c53 <= qM28_c52;
               qP27_c53 <= qP27_c52;
               qM27_c53 <= qM27_c52;
               qP26_c53 <= qP26_c52;
               qM26_c53 <= qM26_c52;
               qP25_c53 <= qP25_c52;
               qM25_c53 <= qM25_c52;
               qP24_c53 <= qP24_c52;
               qM24_c53 <= qM24_c52;
               qP23_c53 <= qP23_c52;
               qM23_c53 <= qM23_c52;
               qP22_c53 <= qP22_c52;
               qM22_c53 <= qM22_c52;
               qP21_c53 <= qP21_c52;
               qM21_c53 <= qM21_c52;
               qP20_c53 <= qP20_c52;
               qM20_c53 <= qM20_c52;
               qP19_c53 <= qP19_c52;
               qM19_c53 <= qM19_c52;
               qP18_c53 <= qP18_c52;
               qM18_c53 <= qM18_c52;
               qP17_c53 <= qP17_c52;
               qM17_c53 <= qM17_c52;
               qP16_c53 <= qP16_c52;
               qM16_c53 <= qM16_c52;
               qP15_c53 <= qP15_c52;
               qM15_c53 <= qM15_c52;
               qP14_c53 <= qP14_c52;
               qM14_c53 <= qM14_c52;
               qP13_c53 <= qP13_c52;
               qM13_c53 <= qM13_c52;
               qP12_c53 <= qP12_c52;
               qM12_c53 <= qM12_c52;
               qP11_c53 <= qP11_c52;
               qM11_c53 <= qM11_c52;
               qP10_c53 <= qP10_c52;
               qM10_c53 <= qM10_c52;
               qP9_c53 <= qP9_c52;
               qM9_c53 <= qM9_c52;
               qP8_c53 <= qP8_c52;
               qM8_c53 <= qM8_c52;
               qP7_c53 <= qP7_c52;
               qM7_c53 <= qM7_c52;
               qP6_c53 <= qP6_c52;
               qM6_c53 <= qM6_c52;
               qP5_c53 <= qP5_c52;
               qM5_c53 <= qM5_c52;
               qP4_c53 <= qP4_c52;
               qM4_c53 <= qM4_c52;
            end if;
            if ce_54 = '1' then
               expR0_c54 <= expR0_c53;
               sR_c54 <= sR_c53;
               exnR0_c54 <= exnR0_c53;
               D_c54 <= D_c53;
               betaw3_c54 <= betaw3_c53;
               q3_copy30_c54 <= q3_copy30_c53;
               qP28_c54 <= qP28_c53;
               qM28_c54 <= qM28_c53;
               qP27_c54 <= qP27_c53;
               qM27_c54 <= qM27_c53;
               qP26_c54 <= qP26_c53;
               qM26_c54 <= qM26_c53;
               qP25_c54 <= qP25_c53;
               qM25_c54 <= qM25_c53;
               qP24_c54 <= qP24_c53;
               qM24_c54 <= qM24_c53;
               qP23_c54 <= qP23_c53;
               qM23_c54 <= qM23_c53;
               qP22_c54 <= qP22_c53;
               qM22_c54 <= qM22_c53;
               qP21_c54 <= qP21_c53;
               qM21_c54 <= qM21_c53;
               qP20_c54 <= qP20_c53;
               qM20_c54 <= qM20_c53;
               qP19_c54 <= qP19_c53;
               qM19_c54 <= qM19_c53;
               qP18_c54 <= qP18_c53;
               qM18_c54 <= qM18_c53;
               qP17_c54 <= qP17_c53;
               qM17_c54 <= qM17_c53;
               qP16_c54 <= qP16_c53;
               qM16_c54 <= qM16_c53;
               qP15_c54 <= qP15_c53;
               qM15_c54 <= qM15_c53;
               qP14_c54 <= qP14_c53;
               qM14_c54 <= qM14_c53;
               qP13_c54 <= qP13_c53;
               qM13_c54 <= qM13_c53;
               qP12_c54 <= qP12_c53;
               qM12_c54 <= qM12_c53;
               qP11_c54 <= qP11_c53;
               qM11_c54 <= qM11_c53;
               qP10_c54 <= qP10_c53;
               qM10_c54 <= qM10_c53;
               qP9_c54 <= qP9_c53;
               qM9_c54 <= qM9_c53;
               qP8_c54 <= qP8_c53;
               qM8_c54 <= qM8_c53;
               qP7_c54 <= qP7_c53;
               qM7_c54 <= qM7_c53;
               qP6_c54 <= qP6_c53;
               qM6_c54 <= qM6_c53;
               qP5_c54 <= qP5_c53;
               qM5_c54 <= qM5_c53;
               qP4_c54 <= qP4_c53;
               qM4_c54 <= qM4_c53;
            end if;
            if ce_55 = '1' then
               expR0_c55 <= expR0_c54;
               sR_c55 <= sR_c54;
               exnR0_c55 <= exnR0_c54;
               D_c55 <= D_c54;
               betaw3_c55 <= betaw3_c54;
               q3_c55 <= q3_c54;
               absq3D_c55 <= absq3D_c54;
               qP28_c55 <= qP28_c54;
               qM28_c55 <= qM28_c54;
               qP27_c55 <= qP27_c54;
               qM27_c55 <= qM27_c54;
               qP26_c55 <= qP26_c54;
               qM26_c55 <= qM26_c54;
               qP25_c55 <= qP25_c54;
               qM25_c55 <= qM25_c54;
               qP24_c55 <= qP24_c54;
               qM24_c55 <= qM24_c54;
               qP23_c55 <= qP23_c54;
               qM23_c55 <= qM23_c54;
               qP22_c55 <= qP22_c54;
               qM22_c55 <= qM22_c54;
               qP21_c55 <= qP21_c54;
               qM21_c55 <= qM21_c54;
               qP20_c55 <= qP20_c54;
               qM20_c55 <= qM20_c54;
               qP19_c55 <= qP19_c54;
               qM19_c55 <= qM19_c54;
               qP18_c55 <= qP18_c54;
               qM18_c55 <= qM18_c54;
               qP17_c55 <= qP17_c54;
               qM17_c55 <= qM17_c54;
               qP16_c55 <= qP16_c54;
               qM16_c55 <= qM16_c54;
               qP15_c55 <= qP15_c54;
               qM15_c55 <= qM15_c54;
               qP14_c55 <= qP14_c54;
               qM14_c55 <= qM14_c54;
               qP13_c55 <= qP13_c54;
               qM13_c55 <= qM13_c54;
               qP12_c55 <= qP12_c54;
               qM12_c55 <= qM12_c54;
               qP11_c55 <= qP11_c54;
               qM11_c55 <= qM11_c54;
               qP10_c55 <= qP10_c54;
               qM10_c55 <= qM10_c54;
               qP9_c55 <= qP9_c54;
               qM9_c55 <= qM9_c54;
               qP8_c55 <= qP8_c54;
               qM8_c55 <= qM8_c54;
               qP7_c55 <= qP7_c54;
               qM7_c55 <= qM7_c54;
               qP6_c55 <= qP6_c54;
               qM6_c55 <= qM6_c54;
               qP5_c55 <= qP5_c54;
               qM5_c55 <= qM5_c54;
               qP4_c55 <= qP4_c54;
               qM4_c55 <= qM4_c54;
               qP3_c55 <= qP3_c54;
               qM3_c55 <= qM3_c54;
            end if;
            if ce_56 = '1' then
               expR0_c56 <= expR0_c55;
               sR_c56 <= sR_c55;
               exnR0_c56 <= exnR0_c55;
               D_c56 <= D_c55;
               betaw2_c56 <= betaw2_c55;
               q2_copy31_c56 <= q2_copy31_c55;
               qP28_c56 <= qP28_c55;
               qM28_c56 <= qM28_c55;
               qP27_c56 <= qP27_c55;
               qM27_c56 <= qM27_c55;
               qP26_c56 <= qP26_c55;
               qM26_c56 <= qM26_c55;
               qP25_c56 <= qP25_c55;
               qM25_c56 <= qM25_c55;
               qP24_c56 <= qP24_c55;
               qM24_c56 <= qM24_c55;
               qP23_c56 <= qP23_c55;
               qM23_c56 <= qM23_c55;
               qP22_c56 <= qP22_c55;
               qM22_c56 <= qM22_c55;
               qP21_c56 <= qP21_c55;
               qM21_c56 <= qM21_c55;
               qP20_c56 <= qP20_c55;
               qM20_c56 <= qM20_c55;
               qP19_c56 <= qP19_c55;
               qM19_c56 <= qM19_c55;
               qP18_c56 <= qP18_c55;
               qM18_c56 <= qM18_c55;
               qP17_c56 <= qP17_c55;
               qM17_c56 <= qM17_c55;
               qP16_c56 <= qP16_c55;
               qM16_c56 <= qM16_c55;
               qP15_c56 <= qP15_c55;
               qM15_c56 <= qM15_c55;
               qP14_c56 <= qP14_c55;
               qM14_c56 <= qM14_c55;
               qP13_c56 <= qP13_c55;
               qM13_c56 <= qM13_c55;
               qP12_c56 <= qP12_c55;
               qM12_c56 <= qM12_c55;
               qP11_c56 <= qP11_c55;
               qM11_c56 <= qM11_c55;
               qP10_c56 <= qP10_c55;
               qM10_c56 <= qM10_c55;
               qP9_c56 <= qP9_c55;
               qM9_c56 <= qM9_c55;
               qP8_c56 <= qP8_c55;
               qM8_c56 <= qM8_c55;
               qP7_c56 <= qP7_c55;
               qM7_c56 <= qM7_c55;
               qP6_c56 <= qP6_c55;
               qM6_c56 <= qM6_c55;
               qP5_c56 <= qP5_c55;
               qM5_c56 <= qM5_c55;
               qP4_c56 <= qP4_c55;
               qM4_c56 <= qM4_c55;
               qP3_c56 <= qP3_c55;
               qM3_c56 <= qM3_c55;
            end if;
            if ce_57 = '1' then
               expR0_c57 <= expR0_c56;
               sR_c57 <= sR_c56;
               exnR0_c57 <= exnR0_c56;
               D_c57 <= D_c56;
               betaw2_c57 <= betaw2_c56;
               q2_c57 <= q2_c56;
               absq2D_c57 <= absq2D_c56;
               qP28_c57 <= qP28_c56;
               qM28_c57 <= qM28_c56;
               qP27_c57 <= qP27_c56;
               qM27_c57 <= qM27_c56;
               qP26_c57 <= qP26_c56;
               qM26_c57 <= qM26_c56;
               qP25_c57 <= qP25_c56;
               qM25_c57 <= qM25_c56;
               qP24_c57 <= qP24_c56;
               qM24_c57 <= qM24_c56;
               qP23_c57 <= qP23_c56;
               qM23_c57 <= qM23_c56;
               qP22_c57 <= qP22_c56;
               qM22_c57 <= qM22_c56;
               qP21_c57 <= qP21_c56;
               qM21_c57 <= qM21_c56;
               qP20_c57 <= qP20_c56;
               qM20_c57 <= qM20_c56;
               qP19_c57 <= qP19_c56;
               qM19_c57 <= qM19_c56;
               qP18_c57 <= qP18_c56;
               qM18_c57 <= qM18_c56;
               qP17_c57 <= qP17_c56;
               qM17_c57 <= qM17_c56;
               qP16_c57 <= qP16_c56;
               qM16_c57 <= qM16_c56;
               qP15_c57 <= qP15_c56;
               qM15_c57 <= qM15_c56;
               qP14_c57 <= qP14_c56;
               qM14_c57 <= qM14_c56;
               qP13_c57 <= qP13_c56;
               qM13_c57 <= qM13_c56;
               qP12_c57 <= qP12_c56;
               qM12_c57 <= qM12_c56;
               qP11_c57 <= qP11_c56;
               qM11_c57 <= qM11_c56;
               qP10_c57 <= qP10_c56;
               qM10_c57 <= qM10_c56;
               qP9_c57 <= qP9_c56;
               qM9_c57 <= qM9_c56;
               qP8_c57 <= qP8_c56;
               qM8_c57 <= qM8_c56;
               qP7_c57 <= qP7_c56;
               qM7_c57 <= qM7_c56;
               qP6_c57 <= qP6_c56;
               qM6_c57 <= qM6_c56;
               qP5_c57 <= qP5_c56;
               qM5_c57 <= qM5_c56;
               qP4_c57 <= qP4_c56;
               qM4_c57 <= qM4_c56;
               qP3_c57 <= qP3_c56;
               qM3_c57 <= qM3_c56;
               qP2_c57 <= qP2_c56;
               qM2_c57 <= qM2_c56;
            end if;
            if ce_58 = '1' then
               expR0_c58 <= expR0_c57;
               sR_c58 <= sR_c57;
               exnR0_c58 <= exnR0_c57;
               D_c58 <= D_c57;
               betaw2_c58 <= betaw2_c57;
               q2_c58 <= q2_c57;
               absq2D_c58 <= absq2D_c57;
               qP28_c58 <= qP28_c57;
               qM28_c58 <= qM28_c57;
               qP27_c58 <= qP27_c57;
               qM27_c58 <= qM27_c57;
               qP26_c58 <= qP26_c57;
               qM26_c58 <= qM26_c57;
               qP25_c58 <= qP25_c57;
               qM25_c58 <= qM25_c57;
               qP24_c58 <= qP24_c57;
               qM24_c58 <= qM24_c57;
               qP23_c58 <= qP23_c57;
               qM23_c58 <= qM23_c57;
               qP22_c58 <= qP22_c57;
               qM22_c58 <= qM22_c57;
               qP21_c58 <= qP21_c57;
               qM21_c58 <= qM21_c57;
               qP20_c58 <= qP20_c57;
               qM20_c58 <= qM20_c57;
               qP19_c58 <= qP19_c57;
               qM19_c58 <= qM19_c57;
               qP18_c58 <= qP18_c57;
               qM18_c58 <= qM18_c57;
               qP17_c58 <= qP17_c57;
               qM17_c58 <= qM17_c57;
               qP16_c58 <= qP16_c57;
               qM16_c58 <= qM16_c57;
               qP15_c58 <= qP15_c57;
               qM15_c58 <= qM15_c57;
               qP14_c58 <= qP14_c57;
               qM14_c58 <= qM14_c57;
               qP13_c58 <= qP13_c57;
               qM13_c58 <= qM13_c57;
               qP12_c58 <= qP12_c57;
               qM12_c58 <= qM12_c57;
               qP11_c58 <= qP11_c57;
               qM11_c58 <= qM11_c57;
               qP10_c58 <= qP10_c57;
               qM10_c58 <= qM10_c57;
               qP9_c58 <= qP9_c57;
               qM9_c58 <= qM9_c57;
               qP8_c58 <= qP8_c57;
               qM8_c58 <= qM8_c57;
               qP7_c58 <= qP7_c57;
               qM7_c58 <= qM7_c57;
               qP6_c58 <= qP6_c57;
               qM6_c58 <= qM6_c57;
               qP5_c58 <= qP5_c57;
               qM5_c58 <= qM5_c57;
               qP4_c58 <= qP4_c57;
               qM4_c58 <= qM4_c57;
               qP3_c58 <= qP3_c57;
               qM3_c58 <= qM3_c57;
               qP2_c58 <= qP2_c57;
               qM2_c58 <= qM2_c57;
            end if;
            if ce_59 = '1' then
               expR0_c59 <= expR0_c58;
               sR_c59 <= sR_c58;
               exnR0_c59 <= exnR0_c58;
               betaw1_c59 <= betaw1_c58;
               q1_c59 <= q1_c58;
               absq1D_c59 <= absq1D_c58;
               qM28_c59 <= qM28_c58;
               qM27_c59 <= qM27_c58;
               qM26_c59 <= qM26_c58;
               qM25_c59 <= qM25_c58;
               qM24_c59 <= qM24_c58;
               qM23_c59 <= qM23_c58;
               qM22_c59 <= qM22_c58;
               qM21_c59 <= qM21_c58;
               qM20_c59 <= qM20_c58;
               qM19_c59 <= qM19_c58;
               qM18_c59 <= qM18_c58;
               qM17_c59 <= qM17_c58;
               qM16_c59 <= qM16_c58;
               qM15_c59 <= qM15_c58;
               qM14_c59 <= qM14_c58;
               qM13_c59 <= qM13_c58;
               qM12_c59 <= qM12_c58;
               qM11_c59 <= qM11_c58;
               qM10_c59 <= qM10_c58;
               qM9_c59 <= qM9_c58;
               qM8_c59 <= qM8_c58;
               qM7_c59 <= qM7_c58;
               qM6_c59 <= qM6_c58;
               qM5_c59 <= qM5_c58;
               qM4_c59 <= qM4_c58;
               qM3_c59 <= qM3_c58;
               qM2_c59 <= qM2_c58;
               qM1_c59 <= qM1_c58;
               qP_c59 <= qP_c58;
            end if;
            if ce_60 = '1' then
               expR0_c60 <= expR0_c59;
               sR_c60 <= sR_c59;
               exnR0_c60 <= exnR0_c59;
               betaw1_c60 <= betaw1_c59;
               q1_c60 <= q1_c59;
               absq1D_c60 <= absq1D_c59;
               qM28_c60 <= qM28_c59;
               qM27_c60 <= qM27_c59;
               qM26_c60 <= qM26_c59;
               qM25_c60 <= qM25_c59;
               qM24_c60 <= qM24_c59;
               qM23_c60 <= qM23_c59;
               qM22_c60 <= qM22_c59;
               qM21_c60 <= qM21_c59;
               qM20_c60 <= qM20_c59;
               qM19_c60 <= qM19_c59;
               qM18_c60 <= qM18_c59;
               qM17_c60 <= qM17_c59;
               qM16_c60 <= qM16_c59;
               qM15_c60 <= qM15_c59;
               qM14_c60 <= qM14_c59;
               qM13_c60 <= qM13_c59;
               qM12_c60 <= qM12_c59;
               qM11_c60 <= qM11_c59;
               qM10_c60 <= qM10_c59;
               qM9_c60 <= qM9_c59;
               qM8_c60 <= qM8_c59;
               qM7_c60 <= qM7_c59;
               qM6_c60 <= qM6_c59;
               qM5_c60 <= qM5_c59;
               qM4_c60 <= qM4_c59;
               qM3_c60 <= qM3_c59;
               qM2_c60 <= qM2_c59;
               qM1_c60 <= qM1_c59;
               qP_c60 <= qP_c59;
            end if;
            if ce_61 = '1' then
               expR0_c61 <= expR0_c60;
               sR_c61 <= sR_c60;
               exnR0_c61 <= exnR0_c60;
               qP_c61 <= qP_c60;
               qM_c61 <= qM_c60;
            end if;
            if ce_62 = '1' then
               expR0_c62 <= expR0_c61;
               sR_c62 <= sR_c61;
               exnR0_c62 <= exnR0_c61;
               mR_c62 <= mR_c61;
               fRnorm_c62 <= fRnorm_c61;
               round_c62 <= round_c61;
            end if;
            if ce_63 = '1' then
               sR_c63 <= sR_c62;
               exnR0_c63 <= exnR0_c62;
               expfracR_c63 <= expfracR_c62;
            end if;
         end if;
      end process;
   fX_c0 <= "1" & X(51 downto 0);
   fY_c0 <= "1" & Y(51 downto 0);
   -- exponent difference, sign and exception combination computed early, to have fewer bits to pipeline
   expR0_c0 <= ("00" & X(62 downto 52)) - ("00" & Y(62 downto 52));
   sR_c0 <= X(63) xor Y(63);
   -- early exception handling 
   exnXY_c0 <= X(65 downto 64) & Y(65 downto 64);
   with exnXY_c0  select 
      exnR0_c0 <= 
         "01"	 when "0101",										-- normal
         "00"	 when "0001" | "0010" | "0110", -- zero
         "10"	 when "0100" | "1000" | "1001", -- overflow
         "11"	 when others;										-- NaN
   D_c0 <= fY_c0 ;
   psX_c0 <= "0" & fX_c0 ;
   betaw28_c0 <=  "00" & psX_c0;
   sel28_c0 <= betaw28_c0(55 downto 50) & D_c0(51 downto 49);
   SelFunctionTable28: selFunction_Freq800_uid4
      port map ( X => sel28_c0,
                 Y => q28_copy5_c0);
   q28_c0 <= q28_copy5_c0; -- output copy to hold a pipeline register if needed

   with q28_c0  select 
      absq28D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q28_c2(2)  select 
   w27_c2<= betaw28_c2 - absq28D_c2 when '0',
         betaw28_c2 + absq28D_c2 when others;

   betaw27_c2 <= w27_c2(53 downto 0) & "00"; -- multiplication by the radix
   sel27_c2 <= betaw27_c2(55 downto 50) & D_c2(51 downto 49);
   SelFunctionTable27: selFunction_Freq800_uid4
      port map ( X => sel27_c2,
                 Y => q27_copy6_c2);
   q27_c2 <= q27_copy6_c2; -- output copy to hold a pipeline register if needed

   with q27_c2  select 
      absq27D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q27_c4(2)  select 
   w26_c4<= betaw27_c4 - absq27D_c4 when '0',
         betaw27_c4 + absq27D_c4 when others;

   betaw26_c4 <= w26_c4(53 downto 0) & "00"; -- multiplication by the radix
   sel26_c4 <= betaw26_c4(55 downto 50) & D_c4(51 downto 49);
   SelFunctionTable26: selFunction_Freq800_uid4
      port map ( X => sel26_c4,
                 Y => q26_copy7_c4);
   q26_c4 <= q26_copy7_c4; -- output copy to hold a pipeline register if needed

   with q26_c4  select 
      absq26D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q26_c6(2)  select 
   w25_c6<= betaw26_c6 - absq26D_c6 when '0',
         betaw26_c6 + absq26D_c6 when others;

   betaw25_c6 <= w25_c6(53 downto 0) & "00"; -- multiplication by the radix
   sel25_c6 <= betaw25_c6(55 downto 50) & D_c6(51 downto 49);
   SelFunctionTable25: selFunction_Freq800_uid4
      port map ( X => sel25_c6,
                 Y => q25_copy8_c6);
   q25_c6 <= q25_copy8_c6; -- output copy to hold a pipeline register if needed

   with q25_c6  select 
      absq25D_c6 <= 
         "000" & D_c6						 when "001" | "111", -- mult by 1
         "00" & D_c6 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q25_c8(2)  select 
   w24_c8<= betaw25_c8 - absq25D_c8 when '0',
         betaw25_c8 + absq25D_c8 when others;

   betaw24_c8 <= w24_c8(53 downto 0) & "00"; -- multiplication by the radix
   sel24_c8 <= betaw24_c8(55 downto 50) & D_c8(51 downto 49);
   SelFunctionTable24: selFunction_Freq800_uid4
      port map ( X => sel24_c8,
                 Y => q24_copy9_c8);
   q24_c9 <= q24_copy9_c9; -- output copy to hold a pipeline register if needed

   with q24_c9  select 
      absq24D_c9 <= 
         "000" & D_c9						 when "001" | "111", -- mult by 1
         "00" & D_c9 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q24_c10(2)  select 
   w23_c10<= betaw24_c10 - absq24D_c10 when '0',
         betaw24_c10 + absq24D_c10 when others;

   betaw23_c10 <= w23_c10(53 downto 0) & "00"; -- multiplication by the radix
   sel23_c10 <= betaw23_c10(55 downto 50) & D_c10(51 downto 49);
   SelFunctionTable23: selFunction_Freq800_uid4
      port map ( X => sel23_c10,
                 Y => q23_copy10_c10);
   q23_c11 <= q23_copy10_c11; -- output copy to hold a pipeline register if needed

   with q23_c11  select 
      absq23D_c11 <= 
         "000" & D_c11						 when "001" | "111", -- mult by 1
         "00" & D_c11 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q23_c12(2)  select 
   w22_c12<= betaw23_c12 - absq23D_c12 when '0',
         betaw23_c12 + absq23D_c12 when others;

   betaw22_c12 <= w22_c12(53 downto 0) & "00"; -- multiplication by the radix
   sel22_c12 <= betaw22_c12(55 downto 50) & D_c12(51 downto 49);
   SelFunctionTable22: selFunction_Freq800_uid4
      port map ( X => sel22_c12,
                 Y => q22_copy11_c12);
   q22_c13 <= q22_copy11_c13; -- output copy to hold a pipeline register if needed

   with q22_c13  select 
      absq22D_c13 <= 
         "000" & D_c13						 when "001" | "111", -- mult by 1
         "00" & D_c13 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q22_c15(2)  select 
   w21_c15<= betaw22_c15 - absq22D_c15 when '0',
         betaw22_c15 + absq22D_c15 when others;

   betaw21_c15 <= w21_c15(53 downto 0) & "00"; -- multiplication by the radix
   sel21_c15 <= betaw21_c15(55 downto 50) & D_c15(51 downto 49);
   SelFunctionTable21: selFunction_Freq800_uid4
      port map ( X => sel21_c15,
                 Y => q21_copy12_c15);
   q21_c15 <= q21_copy12_c15; -- output copy to hold a pipeline register if needed

   with q21_c15  select 
      absq21D_c15 <= 
         "000" & D_c15						 when "001" | "111", -- mult by 1
         "00" & D_c15 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q21_c17(2)  select 
   w20_c17<= betaw21_c17 - absq21D_c17 when '0',
         betaw21_c17 + absq21D_c17 when others;

   betaw20_c17 <= w20_c17(53 downto 0) & "00"; -- multiplication by the radix
   sel20_c17 <= betaw20_c17(55 downto 50) & D_c17(51 downto 49);
   SelFunctionTable20: selFunction_Freq800_uid4
      port map ( X => sel20_c17,
                 Y => q20_copy13_c17);
   q20_c17 <= q20_copy13_c17; -- output copy to hold a pipeline register if needed

   with q20_c17  select 
      absq20D_c17 <= 
         "000" & D_c17						 when "001" | "111", -- mult by 1
         "00" & D_c17 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q20_c19(2)  select 
   w19_c19<= betaw20_c19 - absq20D_c19 when '0',
         betaw20_c19 + absq20D_c19 when others;

   betaw19_c19 <= w19_c19(53 downto 0) & "00"; -- multiplication by the radix
   sel19_c19 <= betaw19_c19(55 downto 50) & D_c19(51 downto 49);
   SelFunctionTable19: selFunction_Freq800_uid4
      port map ( X => sel19_c19,
                 Y => q19_copy14_c19);
   q19_c19 <= q19_copy14_c19; -- output copy to hold a pipeline register if needed

   with q19_c19  select 
      absq19D_c19 <= 
         "000" & D_c19						 when "001" | "111", -- mult by 1
         "00" & D_c19 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q19_c21(2)  select 
   w18_c21<= betaw19_c21 - absq19D_c21 when '0',
         betaw19_c21 + absq19D_c21 when others;

   betaw18_c21 <= w18_c21(53 downto 0) & "00"; -- multiplication by the radix
   sel18_c21 <= betaw18_c21(55 downto 50) & D_c21(51 downto 49);
   SelFunctionTable18: selFunction_Freq800_uid4
      port map ( X => sel18_c21,
                 Y => q18_copy15_c21);
   q18_c22 <= q18_copy15_c22; -- output copy to hold a pipeline register if needed

   with q18_c22  select 
      absq18D_c22 <= 
         "000" & D_c22						 when "001" | "111", -- mult by 1
         "00" & D_c22 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q18_c23(2)  select 
   w17_c23<= betaw18_c23 - absq18D_c23 when '0',
         betaw18_c23 + absq18D_c23 when others;

   betaw17_c23 <= w17_c23(53 downto 0) & "00"; -- multiplication by the radix
   sel17_c23 <= betaw17_c23(55 downto 50) & D_c23(51 downto 49);
   SelFunctionTable17: selFunction_Freq800_uid4
      port map ( X => sel17_c23,
                 Y => q17_copy16_c23);
   q17_c24 <= q17_copy16_c24; -- output copy to hold a pipeline register if needed

   with q17_c24  select 
      absq17D_c24 <= 
         "000" & D_c24						 when "001" | "111", -- mult by 1
         "00" & D_c24 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q17_c25(2)  select 
   w16_c25<= betaw17_c25 - absq17D_c25 when '0',
         betaw17_c25 + absq17D_c25 when others;

   betaw16_c25 <= w16_c25(53 downto 0) & "00"; -- multiplication by the radix
   sel16_c25 <= betaw16_c25(55 downto 50) & D_c25(51 downto 49);
   SelFunctionTable16: selFunction_Freq800_uid4
      port map ( X => sel16_c25,
                 Y => q16_copy17_c25);
   q16_c26 <= q16_copy17_c26; -- output copy to hold a pipeline register if needed

   with q16_c26  select 
      absq16D_c26 <= 
         "000" & D_c26						 when "001" | "111", -- mult by 1
         "00" & D_c26 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q16_c27(2)  select 
   w15_c27<= betaw16_c27 - absq16D_c27 when '0',
         betaw16_c27 + absq16D_c27 when others;

   betaw15_c27 <= w15_c27(53 downto 0) & "00"; -- multiplication by the radix
   sel15_c27 <= betaw15_c27(55 downto 50) & D_c27(51 downto 49);
   SelFunctionTable15: selFunction_Freq800_uid4
      port map ( X => sel15_c27,
                 Y => q15_copy18_c27);
   q15_c28 <= q15_copy18_c28; -- output copy to hold a pipeline register if needed

   with q15_c28  select 
      absq15D_c28 <= 
         "000" & D_c28						 when "001" | "111", -- mult by 1
         "00" & D_c28 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q15_c30(2)  select 
   w14_c30<= betaw15_c30 - absq15D_c30 when '0',
         betaw15_c30 + absq15D_c30 when others;

   betaw14_c30 <= w14_c30(53 downto 0) & "00"; -- multiplication by the radix
   sel14_c30 <= betaw14_c30(55 downto 50) & D_c30(51 downto 49);
   SelFunctionTable14: selFunction_Freq800_uid4
      port map ( X => sel14_c30,
                 Y => q14_copy19_c30);
   q14_c30 <= q14_copy19_c30; -- output copy to hold a pipeline register if needed

   with q14_c30  select 
      absq14D_c30 <= 
         "000" & D_c30						 when "001" | "111", -- mult by 1
         "00" & D_c30 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q14_c32(2)  select 
   w13_c32<= betaw14_c32 - absq14D_c32 when '0',
         betaw14_c32 + absq14D_c32 when others;

   betaw13_c32 <= w13_c32(53 downto 0) & "00"; -- multiplication by the radix
   sel13_c32 <= betaw13_c32(55 downto 50) & D_c32(51 downto 49);
   SelFunctionTable13: selFunction_Freq800_uid4
      port map ( X => sel13_c32,
                 Y => q13_copy20_c32);
   q13_c32 <= q13_copy20_c32; -- output copy to hold a pipeline register if needed

   with q13_c32  select 
      absq13D_c32 <= 
         "000" & D_c32						 when "001" | "111", -- mult by 1
         "00" & D_c32 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q13_c34(2)  select 
   w12_c34<= betaw13_c34 - absq13D_c34 when '0',
         betaw13_c34 + absq13D_c34 when others;

   betaw12_c34 <= w12_c34(53 downto 0) & "00"; -- multiplication by the radix
   sel12_c34 <= betaw12_c34(55 downto 50) & D_c34(51 downto 49);
   SelFunctionTable12: selFunction_Freq800_uid4
      port map ( X => sel12_c34,
                 Y => q12_copy21_c34);
   q12_c34 <= q12_copy21_c34; -- output copy to hold a pipeline register if needed

   with q12_c34  select 
      absq12D_c34 <= 
         "000" & D_c34						 when "001" | "111", -- mult by 1
         "00" & D_c34 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q12_c36(2)  select 
   w11_c36<= betaw12_c36 - absq12D_c36 when '0',
         betaw12_c36 + absq12D_c36 when others;

   betaw11_c36 <= w11_c36(53 downto 0) & "00"; -- multiplication by the radix
   sel11_c36 <= betaw11_c36(55 downto 50) & D_c36(51 downto 49);
   SelFunctionTable11: selFunction_Freq800_uid4
      port map ( X => sel11_c36,
                 Y => q11_copy22_c36);
   q11_c37 <= q11_copy22_c37; -- output copy to hold a pipeline register if needed

   with q11_c37  select 
      absq11D_c37 <= 
         "000" & D_c37						 when "001" | "111", -- mult by 1
         "00" & D_c37 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q11_c38(2)  select 
   w10_c38<= betaw11_c38 - absq11D_c38 when '0',
         betaw11_c38 + absq11D_c38 when others;

   betaw10_c38 <= w10_c38(53 downto 0) & "00"; -- multiplication by the radix
   sel10_c38 <= betaw10_c38(55 downto 50) & D_c38(51 downto 49);
   SelFunctionTable10: selFunction_Freq800_uid4
      port map ( X => sel10_c38,
                 Y => q10_copy23_c38);
   q10_c39 <= q10_copy23_c39; -- output copy to hold a pipeline register if needed

   with q10_c39  select 
      absq10D_c39 <= 
         "000" & D_c39						 when "001" | "111", -- mult by 1
         "00" & D_c39 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q10_c40(2)  select 
   w9_c40<= betaw10_c40 - absq10D_c40 when '0',
         betaw10_c40 + absq10D_c40 when others;

   betaw9_c40 <= w9_c40(53 downto 0) & "00"; -- multiplication by the radix
   sel9_c40 <= betaw9_c40(55 downto 50) & D_c40(51 downto 49);
   SelFunctionTable9: selFunction_Freq800_uid4
      port map ( X => sel9_c40,
                 Y => q9_copy24_c40);
   q9_c41 <= q9_copy24_c41; -- output copy to hold a pipeline register if needed

   with q9_c41  select 
      absq9D_c41 <= 
         "000" & D_c41						 when "001" | "111", -- mult by 1
         "00" & D_c41 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q9_c42(2)  select 
   w8_c42<= betaw9_c42 - absq9D_c42 when '0',
         betaw9_c42 + absq9D_c42 when others;

   betaw8_c42 <= w8_c42(53 downto 0) & "00"; -- multiplication by the radix
   sel8_c42 <= betaw8_c42(55 downto 50) & D_c42(51 downto 49);
   SelFunctionTable8: selFunction_Freq800_uid4
      port map ( X => sel8_c42,
                 Y => q8_copy25_c42);
   q8_c43 <= q8_copy25_c43; -- output copy to hold a pipeline register if needed

   with q8_c43  select 
      absq8D_c43 <= 
         "000" & D_c43						 when "001" | "111", -- mult by 1
         "00" & D_c43 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q8_c45(2)  select 
   w7_c45<= betaw8_c45 - absq8D_c45 when '0',
         betaw8_c45 + absq8D_c45 when others;

   betaw7_c45 <= w7_c45(53 downto 0) & "00"; -- multiplication by the radix
   sel7_c45 <= betaw7_c45(55 downto 50) & D_c45(51 downto 49);
   SelFunctionTable7: selFunction_Freq800_uid4
      port map ( X => sel7_c45,
                 Y => q7_copy26_c45);
   q7_c45 <= q7_copy26_c45; -- output copy to hold a pipeline register if needed

   with q7_c45  select 
      absq7D_c45 <= 
         "000" & D_c45						 when "001" | "111", -- mult by 1
         "00" & D_c45 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q7_c47(2)  select 
   w6_c47<= betaw7_c47 - absq7D_c47 when '0',
         betaw7_c47 + absq7D_c47 when others;

   betaw6_c47 <= w6_c47(53 downto 0) & "00"; -- multiplication by the radix
   sel6_c47 <= betaw6_c47(55 downto 50) & D_c47(51 downto 49);
   SelFunctionTable6: selFunction_Freq800_uid4
      port map ( X => sel6_c47,
                 Y => q6_copy27_c47);
   q6_c47 <= q6_copy27_c47; -- output copy to hold a pipeline register if needed

   with q6_c47  select 
      absq6D_c47 <= 
         "000" & D_c47						 when "001" | "111", -- mult by 1
         "00" & D_c47 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q6_c49(2)  select 
   w5_c49<= betaw6_c49 - absq6D_c49 when '0',
         betaw6_c49 + absq6D_c49 when others;

   betaw5_c49 <= w5_c49(53 downto 0) & "00"; -- multiplication by the radix
   sel5_c49 <= betaw5_c49(55 downto 50) & D_c49(51 downto 49);
   SelFunctionTable5: selFunction_Freq800_uid4
      port map ( X => sel5_c49,
                 Y => q5_copy28_c49);
   q5_c49 <= q5_copy28_c49; -- output copy to hold a pipeline register if needed

   with q5_c49  select 
      absq5D_c49 <= 
         "000" & D_c49						 when "001" | "111", -- mult by 1
         "00" & D_c49 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q5_c51(2)  select 
   w4_c51<= betaw5_c51 - absq5D_c51 when '0',
         betaw5_c51 + absq5D_c51 when others;

   betaw4_c51 <= w4_c51(53 downto 0) & "00"; -- multiplication by the radix
   sel4_c51 <= betaw4_c51(55 downto 50) & D_c51(51 downto 49);
   SelFunctionTable4: selFunction_Freq800_uid4
      port map ( X => sel4_c51,
                 Y => q4_copy29_c51);
   q4_c52 <= q4_copy29_c52; -- output copy to hold a pipeline register if needed

   with q4_c52  select 
      absq4D_c52 <= 
         "000" & D_c52						 when "001" | "111", -- mult by 1
         "00" & D_c52 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q4_c53(2)  select 
   w3_c53<= betaw4_c53 - absq4D_c53 when '0',
         betaw4_c53 + absq4D_c53 when others;

   betaw3_c53 <= w3_c53(53 downto 0) & "00"; -- multiplication by the radix
   sel3_c53 <= betaw3_c53(55 downto 50) & D_c53(51 downto 49);
   SelFunctionTable3: selFunction_Freq800_uid4
      port map ( X => sel3_c53,
                 Y => q3_copy30_c53);
   q3_c54 <= q3_copy30_c54; -- output copy to hold a pipeline register if needed

   with q3_c54  select 
      absq3D_c54 <= 
         "000" & D_c54						 when "001" | "111", -- mult by 1
         "00" & D_c54 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q3_c55(2)  select 
   w2_c55<= betaw3_c55 - absq3D_c55 when '0',
         betaw3_c55 + absq3D_c55 when others;

   betaw2_c55 <= w2_c55(53 downto 0) & "00"; -- multiplication by the radix
   sel2_c55 <= betaw2_c55(55 downto 50) & D_c55(51 downto 49);
   SelFunctionTable2: selFunction_Freq800_uid4
      port map ( X => sel2_c55,
                 Y => q2_copy31_c55);
   q2_c56 <= q2_copy31_c56; -- output copy to hold a pipeline register if needed

   with q2_c56  select 
      absq2D_c56 <= 
         "000" & D_c56						 when "001" | "111", -- mult by 1
         "00" & D_c56 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q2_c58(2)  select 
   w1_c58<= betaw2_c58 - absq2D_c58 when '0',
         betaw2_c58 + absq2D_c58 when others;

   betaw1_c58 <= w1_c58(53 downto 0) & "00"; -- multiplication by the radix
   sel1_c58 <= betaw1_c58(55 downto 50) & D_c58(51 downto 49);
   SelFunctionTable1: selFunction_Freq800_uid4
      port map ( X => sel1_c58,
                 Y => q1_copy32_c58);
   q1_c58 <= q1_copy32_c58; -- output copy to hold a pipeline register if needed

   with q1_c58  select 
      absq1D_c58 <= 
         "000" & D_c58						 when "001" | "111", -- mult by 1
         "00" & D_c58 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q1_c60(2)  select 
   w0_c60<= betaw1_c60 - absq1D_c60 when '0',
         betaw1_c60 + absq1D_c60 when others;

   wfinal_c60 <= w0_c60(53 downto 0);
   qM0_c60 <= wfinal_c60(53); -- rounding bit is the sign of the remainder
   qP28_c0 <=      q28_c0(1 downto 0);
   qM28_c0 <=      q28_c0(2) & "0";
   qP27_c2 <=      q27_c2(1 downto 0);
   qM27_c2 <=      q27_c2(2) & "0";
   qP26_c4 <=      q26_c4(1 downto 0);
   qM26_c4 <=      q26_c4(2) & "0";
   qP25_c6 <=      q25_c6(1 downto 0);
   qM25_c6 <=      q25_c6(2) & "0";
   qP24_c9 <=      q24_c9(1 downto 0);
   qM24_c9 <=      q24_c9(2) & "0";
   qP23_c11 <=      q23_c11(1 downto 0);
   qM23_c11 <=      q23_c11(2) & "0";
   qP22_c13 <=      q22_c13(1 downto 0);
   qM22_c13 <=      q22_c13(2) & "0";
   qP21_c15 <=      q21_c15(1 downto 0);
   qM21_c15 <=      q21_c15(2) & "0";
   qP20_c17 <=      q20_c17(1 downto 0);
   qM20_c17 <=      q20_c17(2) & "0";
   qP19_c19 <=      q19_c19(1 downto 0);
   qM19_c19 <=      q19_c19(2) & "0";
   qP18_c22 <=      q18_c22(1 downto 0);
   qM18_c22 <=      q18_c22(2) & "0";
   qP17_c24 <=      q17_c24(1 downto 0);
   qM17_c24 <=      q17_c24(2) & "0";
   qP16_c26 <=      q16_c26(1 downto 0);
   qM16_c26 <=      q16_c26(2) & "0";
   qP15_c28 <=      q15_c28(1 downto 0);
   qM15_c28 <=      q15_c28(2) & "0";
   qP14_c30 <=      q14_c30(1 downto 0);
   qM14_c30 <=      q14_c30(2) & "0";
   qP13_c32 <=      q13_c32(1 downto 0);
   qM13_c32 <=      q13_c32(2) & "0";
   qP12_c34 <=      q12_c34(1 downto 0);
   qM12_c34 <=      q12_c34(2) & "0";
   qP11_c37 <=      q11_c37(1 downto 0);
   qM11_c37 <=      q11_c37(2) & "0";
   qP10_c39 <=      q10_c39(1 downto 0);
   qM10_c39 <=      q10_c39(2) & "0";
   qP9_c41 <=      q9_c41(1 downto 0);
   qM9_c41 <=      q9_c41(2) & "0";
   qP8_c43 <=      q8_c43(1 downto 0);
   qM8_c43 <=      q8_c43(2) & "0";
   qP7_c45 <=      q7_c45(1 downto 0);
   qM7_c45 <=      q7_c45(2) & "0";
   qP6_c47 <=      q6_c47(1 downto 0);
   qM6_c47 <=      q6_c47(2) & "0";
   qP5_c49 <=      q5_c49(1 downto 0);
   qM5_c49 <=      q5_c49(2) & "0";
   qP4_c52 <=      q4_c52(1 downto 0);
   qM4_c52 <=      q4_c52(2) & "0";
   qP3_c54 <=      q3_c54(1 downto 0);
   qM3_c54 <=      q3_c54(2) & "0";
   qP2_c56 <=      q2_c56(1 downto 0);
   qM2_c56 <=      q2_c56(2) & "0";
   qP1_c58 <=      q1_c58(1 downto 0);
   qM1_c58 <=      q1_c58(2) & "0";
   qP_c58 <= qP28_c58 & qP27_c58 & qP26_c58 & qP25_c58 & qP24_c58 & qP23_c58 & qP22_c58 & qP21_c58 & qP20_c58 & qP19_c58 & qP18_c58 & qP17_c58 & qP16_c58 & qP15_c58 & qP14_c58 & qP13_c58 & qP12_c58 & qP11_c58 & qP10_c58 & qP9_c58 & qP8_c58 & qP7_c58 & qP6_c58 & qP5_c58 & qP4_c58 & qP3_c58 & qP2_c58 & qP1_c58;
   qM_c60 <= qM28_c60(0) & qM27_c60 & qM26_c60 & qM25_c60 & qM24_c60 & qM23_c60 & qM22_c60 & qM21_c60 & qM20_c60 & qM19_c60 & qM18_c60 & qM17_c60 & qM16_c60 & qM15_c60 & qM14_c60 & qM13_c60 & qM12_c60 & qM11_c60 & qM10_c60 & qM9_c60 & qM8_c60 & qM7_c60 & qM6_c60 & qM5_c60 & qM4_c60 & qM3_c60 & qM2_c60 & qM1_c60 & qM0_c60;
   quotient_c61 <= qP_c61 - qM_c61;
   -- We need a mR in (0, -wf-2) format: 1+wF fraction bits, 1 round bit, and 1 guard bit for the normalisation,
   -- quotient is the truncation of the exact quotient to at least 2^(-wF-2) bits
   -- now discarding its possible known MSB zeroes, and dropping the possible extra LSB bit (due to radix 4) 
   mR_c61 <= quotient_c61(54 downto 0); 
   -- normalisation
   fRnorm_c61 <=    mR_c61(53 downto 1)  when mR_c61(54)= '1'
           else mR_c61(52 downto 0);  -- now fRnorm is a (-1, -wF-1) fraction
   round_c61 <= fRnorm_c61(0); 
   expR1_c62 <= expR0_c62 + ("000" & (9 downto 1 => '1') & mR_c62(54)); -- add back bias
   -- final rounding
   expfrac_c62 <= expR1_c62 & fRnorm_c62(52 downto 1) ;
   expfracR_c62 <= expfrac_c62 + ((64 downto 1 => '0') & round_c62);
   exnR_c63 <=      "00"  when expfracR_c63(64) = '1'   -- underflow
           else "10"  when  expfracR_c63(64 downto 63) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_c63  select 
      exnRfinal_c63 <= 
         exnR_c63   when "01", -- normal
         exnR0_c63  when others;
   R <= exnRfinal_c63 & sR_c63 & expfracR_c63(62 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          selFunction_Freq500_uid4
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity selFunction_Freq500_uid4 is
    port (X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of selFunction_Freq500_uid4 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000000000",
      "000" when "000000001",
      "000" when "000000010",
      "000" when "000000011",
      "000" when "000000100",
      "000" when "000000101",
      "000" when "000000110",
      "000" when "000000111",
      "000" when "000001000",
      "000" when "000001001",
      "000" when "000001010",
      "000" when "000001011",
      "000" when "000001100",
      "000" when "000001101",
      "000" when "000001110",
      "000" when "000001111",
      "001" when "000010000",
      "000" when "000010001",
      "000" when "000010010",
      "000" when "000010011",
      "000" when "000010100",
      "000" when "000010101",
      "000" when "000010110",
      "000" when "000010111",
      "001" when "000011000",
      "001" when "000011001",
      "001" when "000011010",
      "001" when "000011011",
      "000" when "000011100",
      "000" when "000011101",
      "000" when "000011110",
      "000" when "000011111",
      "001" when "000100000",
      "001" when "000100001",
      "001" when "000100010",
      "001" when "000100011",
      "001" when "000100100",
      "001" when "000100101",
      "001" when "000100110",
      "000" when "000100111",
      "001" when "000101000",
      "001" when "000101001",
      "001" when "000101010",
      "001" when "000101011",
      "001" when "000101100",
      "001" when "000101101",
      "001" when "000101110",
      "001" when "000101111",
      "010" when "000110000",
      "001" when "000110001",
      "001" when "000110010",
      "001" when "000110011",
      "001" when "000110100",
      "001" when "000110101",
      "001" when "000110110",
      "001" when "000110111",
      "010" when "000111000",
      "010" when "000111001",
      "001" when "000111010",
      "001" when "000111011",
      "001" when "000111100",
      "001" when "000111101",
      "001" when "000111110",
      "001" when "000111111",
      "010" when "001000000",
      "010" when "001000001",
      "010" when "001000010",
      "001" when "001000011",
      "001" when "001000100",
      "001" when "001000101",
      "001" when "001000110",
      "001" when "001000111",
      "010" when "001001000",
      "010" when "001001001",
      "010" when "001001010",
      "010" when "001001011",
      "001" when "001001100",
      "001" when "001001101",
      "001" when "001001110",
      "001" when "001001111",
      "010" when "001010000",
      "010" when "001010001",
      "010" when "001010010",
      "010" when "001010011",
      "010" when "001010100",
      "010" when "001010101",
      "001" when "001010110",
      "001" when "001010111",
      "010" when "001011000",
      "010" when "001011001",
      "010" when "001011010",
      "010" when "001011011",
      "010" when "001011100",
      "010" when "001011101",
      "010" when "001011110",
      "001" when "001011111",
      "010" when "001100000",
      "010" when "001100001",
      "010" when "001100010",
      "010" when "001100011",
      "010" when "001100100",
      "010" when "001100101",
      "010" when "001100110",
      "010" when "001100111",
      "010" when "001101000",
      "010" when "001101001",
      "010" when "001101010",
      "010" when "001101011",
      "010" when "001101100",
      "010" when "001101101",
      "010" when "001101110",
      "010" when "001101111",
      "010" when "001110000",
      "010" when "001110001",
      "010" when "001110010",
      "010" when "001110011",
      "010" when "001110100",
      "010" when "001110101",
      "010" when "001110110",
      "010" when "001110111",
      "010" when "001111000",
      "010" when "001111001",
      "010" when "001111010",
      "010" when "001111011",
      "010" when "001111100",
      "010" when "001111101",
      "010" when "001111110",
      "010" when "001111111",
      "010" when "010000000",
      "010" when "010000001",
      "010" when "010000010",
      "010" when "010000011",
      "010" when "010000100",
      "010" when "010000101",
      "010" when "010000110",
      "010" when "010000111",
      "010" when "010001000",
      "010" when "010001001",
      "010" when "010001010",
      "010" when "010001011",
      "010" when "010001100",
      "010" when "010001101",
      "010" when "010001110",
      "010" when "010001111",
      "010" when "010010000",
      "010" when "010010001",
      "010" when "010010010",
      "010" when "010010011",
      "010" when "010010100",
      "010" when "010010101",
      "010" when "010010110",
      "010" when "010010111",
      "010" when "010011000",
      "010" when "010011001",
      "010" when "010011010",
      "010" when "010011011",
      "010" when "010011100",
      "010" when "010011101",
      "010" when "010011110",
      "010" when "010011111",
      "010" when "010100000",
      "010" when "010100001",
      "010" when "010100010",
      "010" when "010100011",
      "010" when "010100100",
      "010" when "010100101",
      "010" when "010100110",
      "010" when "010100111",
      "010" when "010101000",
      "010" when "010101001",
      "010" when "010101010",
      "010" when "010101011",
      "010" when "010101100",
      "010" when "010101101",
      "010" when "010101110",
      "010" when "010101111",
      "010" when "010110000",
      "010" when "010110001",
      "010" when "010110010",
      "010" when "010110011",
      "010" when "010110100",
      "010" when "010110101",
      "010" when "010110110",
      "010" when "010110111",
      "010" when "010111000",
      "010" when "010111001",
      "010" when "010111010",
      "010" when "010111011",
      "010" when "010111100",
      "010" when "010111101",
      "010" when "010111110",
      "010" when "010111111",
      "010" when "011000000",
      "010" when "011000001",
      "010" when "011000010",
      "010" when "011000011",
      "010" when "011000100",
      "010" when "011000101",
      "010" when "011000110",
      "010" when "011000111",
      "010" when "011001000",
      "010" when "011001001",
      "010" when "011001010",
      "010" when "011001011",
      "010" when "011001100",
      "010" when "011001101",
      "010" when "011001110",
      "010" when "011001111",
      "010" when "011010000",
      "010" when "011010001",
      "010" when "011010010",
      "010" when "011010011",
      "010" when "011010100",
      "010" when "011010101",
      "010" when "011010110",
      "010" when "011010111",
      "010" when "011011000",
      "010" when "011011001",
      "010" when "011011010",
      "010" when "011011011",
      "010" when "011011100",
      "010" when "011011101",
      "010" when "011011110",
      "010" when "011011111",
      "010" when "011100000",
      "010" when "011100001",
      "010" when "011100010",
      "010" when "011100011",
      "010" when "011100100",
      "010" when "011100101",
      "010" when "011100110",
      "010" when "011100111",
      "010" when "011101000",
      "010" when "011101001",
      "010" when "011101010",
      "010" when "011101011",
      "010" when "011101100",
      "010" when "011101101",
      "010" when "011101110",
      "010" when "011101111",
      "010" when "011110000",
      "010" when "011110001",
      "010" when "011110010",
      "010" when "011110011",
      "010" when "011110100",
      "010" when "011110101",
      "010" when "011110110",
      "010" when "011110111",
      "010" when "011111000",
      "010" when "011111001",
      "010" when "011111010",
      "010" when "011111011",
      "010" when "011111100",
      "010" when "011111101",
      "010" when "011111110",
      "010" when "011111111",
      "110" when "100000000",
      "110" when "100000001",
      "110" when "100000010",
      "110" when "100000011",
      "110" when "100000100",
      "110" when "100000101",
      "110" when "100000110",
      "110" when "100000111",
      "110" when "100001000",
      "110" when "100001001",
      "110" when "100001010",
      "110" when "100001011",
      "110" when "100001100",
      "110" when "100001101",
      "110" when "100001110",
      "110" when "100001111",
      "110" when "100010000",
      "110" when "100010001",
      "110" when "100010010",
      "110" when "100010011",
      "110" when "100010100",
      "110" when "100010101",
      "110" when "100010110",
      "110" when "100010111",
      "110" when "100011000",
      "110" when "100011001",
      "110" when "100011010",
      "110" when "100011011",
      "110" when "100011100",
      "110" when "100011101",
      "110" when "100011110",
      "110" when "100011111",
      "110" when "100100000",
      "110" when "100100001",
      "110" when "100100010",
      "110" when "100100011",
      "110" when "100100100",
      "110" when "100100101",
      "110" when "100100110",
      "110" when "100100111",
      "110" when "100101000",
      "110" when "100101001",
      "110" when "100101010",
      "110" when "100101011",
      "110" when "100101100",
      "110" when "100101101",
      "110" when "100101110",
      "110" when "100101111",
      "110" when "100110000",
      "110" when "100110001",
      "110" when "100110010",
      "110" when "100110011",
      "110" when "100110100",
      "110" when "100110101",
      "110" when "100110110",
      "110" when "100110111",
      "110" when "100111000",
      "110" when "100111001",
      "110" when "100111010",
      "110" when "100111011",
      "110" when "100111100",
      "110" when "100111101",
      "110" when "100111110",
      "110" when "100111111",
      "110" when "101000000",
      "110" when "101000001",
      "110" when "101000010",
      "110" when "101000011",
      "110" when "101000100",
      "110" when "101000101",
      "110" when "101000110",
      "110" when "101000111",
      "110" when "101001000",
      "110" when "101001001",
      "110" when "101001010",
      "110" when "101001011",
      "110" when "101001100",
      "110" when "101001101",
      "110" when "101001110",
      "110" when "101001111",
      "110" when "101010000",
      "110" when "101010001",
      "110" when "101010010",
      "110" when "101010011",
      "110" when "101010100",
      "110" when "101010101",
      "110" when "101010110",
      "110" when "101010111",
      "110" when "101011000",
      "110" when "101011001",
      "110" when "101011010",
      "110" when "101011011",
      "110" when "101011100",
      "110" when "101011101",
      "110" when "101011110",
      "110" when "101011111",
      "110" when "101100000",
      "110" when "101100001",
      "110" when "101100010",
      "110" when "101100011",
      "110" when "101100100",
      "110" when "101100101",
      "110" when "101100110",
      "110" when "101100111",
      "110" when "101101000",
      "110" when "101101001",
      "110" when "101101010",
      "110" when "101101011",
      "110" when "101101100",
      "110" when "101101101",
      "110" when "101101110",
      "110" when "101101111",
      "110" when "101110000",
      "110" when "101110001",
      "110" when "101110010",
      "110" when "101110011",
      "110" when "101110100",
      "110" when "101110101",
      "110" when "101110110",
      "110" when "101110111",
      "110" when "101111000",
      "110" when "101111001",
      "110" when "101111010",
      "110" when "101111011",
      "110" when "101111100",
      "110" when "101111101",
      "110" when "101111110",
      "110" when "101111111",
      "110" when "110000000",
      "110" when "110000001",
      "110" when "110000010",
      "110" when "110000011",
      "110" when "110000100",
      "110" when "110000101",
      "110" when "110000110",
      "110" when "110000111",
      "110" when "110001000",
      "110" when "110001001",
      "110" when "110001010",
      "110" when "110001011",
      "110" when "110001100",
      "110" when "110001101",
      "110" when "110001110",
      "110" when "110001111",
      "110" when "110010000",
      "110" when "110010001",
      "110" when "110010010",
      "110" when "110010011",
      "110" when "110010100",
      "110" when "110010101",
      "110" when "110010110",
      "110" when "110010111",
      "110" when "110011000",
      "110" when "110011001",
      "110" when "110011010",
      "110" when "110011011",
      "110" when "110011100",
      "110" when "110011101",
      "110" when "110011110",
      "110" when "110011111",
      "110" when "110100000",
      "110" when "110100001",
      "110" when "110100010",
      "110" when "110100011",
      "110" when "110100100",
      "110" when "110100101",
      "110" when "110100110",
      "110" when "110100111",
      "110" when "110101000",
      "110" when "110101001",
      "110" when "110101010",
      "110" when "110101011",
      "110" when "110101100",
      "110" when "110101101",
      "110" when "110101110",
      "111" when "110101111",
      "110" when "110110000",
      "110" when "110110001",
      "110" when "110110010",
      "110" when "110110011",
      "110" when "110110100",
      "111" when "110110101",
      "111" when "110110110",
      "111" when "110110111",
      "110" when "110111000",
      "110" when "110111001",
      "110" when "110111010",
      "110" when "110111011",
      "111" when "110111100",
      "111" when "110111101",
      "111" when "110111110",
      "111" when "110111111",
      "110" when "111000000",
      "110" when "111000001",
      "111" when "111000010",
      "111" when "111000011",
      "111" when "111000100",
      "111" when "111000101",
      "111" when "111000110",
      "111" when "111000111",
      "110" when "111001000",
      "111" when "111001001",
      "111" when "111001010",
      "111" when "111001011",
      "111" when "111001100",
      "111" when "111001101",
      "111" when "111001110",
      "111" when "111001111",
      "111" when "111010000",
      "111" when "111010001",
      "111" when "111010010",
      "111" when "111010011",
      "111" when "111010100",
      "111" when "111010101",
      "111" when "111010110",
      "111" when "111010111",
      "111" when "111011000",
      "111" when "111011001",
      "111" when "111011010",
      "111" when "111011011",
      "111" when "111011100",
      "111" when "111011101",
      "111" when "111011110",
      "111" when "111011111",
      "111" when "111100000",
      "111" when "111100001",
      "111" when "111100010",
      "111" when "111100011",
      "111" when "111100100",
      "111" when "111100101",
      "111" when "111100110",
      "111" when "111100111",
      "111" when "111101000",
      "111" when "111101001",
      "111" when "111101010",
      "111" when "111101011",
      "000" when "111101100",
      "000" when "111101101",
      "000" when "111101110",
      "000" when "111101111",
      "000" when "111110000",
      "000" when "111110001",
      "000" when "111110010",
      "000" when "111110011",
      "000" when "111110100",
      "000" when "111110101",
      "000" when "111110110",
      "000" when "111110111",
      "000" when "111111000",
      "000" when "111111001",
      "000" when "111111010",
      "000" when "111111011",
      "000" when "111111100",
      "000" when "111111101",
      "000" when "111111110",
      "000" when "111111111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            FloatingPointDivider
--                         (FPDiv_11_52_Freq500_uid2)
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 36 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointDivider_64_4_398000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20, ce_21, ce_22, ce_23, ce_24, ce_25, ce_26, ce_27, ce_28, ce_29, ce_30, ce_31, ce_32, ce_33, ce_34, ce_35, ce_36 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointDivider_64_4_398000 is
   component selFunction_Freq500_uid4 is
      port ( X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal fX_c0 :  std_logic_vector(52 downto 0);
signal fY_c0 :  std_logic_vector(52 downto 0);
signal expR0_c0, expR0_c1, expR0_c2, expR0_c3, expR0_c4, expR0_c5, expR0_c6, expR0_c7, expR0_c8, expR0_c9, expR0_c10, expR0_c11, expR0_c12, expR0_c13, expR0_c14, expR0_c15, expR0_c16, expR0_c17, expR0_c18, expR0_c19, expR0_c20, expR0_c21, expR0_c22, expR0_c23, expR0_c24, expR0_c25, expR0_c26, expR0_c27, expR0_c28, expR0_c29, expR0_c30, expR0_c31, expR0_c32, expR0_c33, expR0_c34, expR0_c35, expR0_c36 :  std_logic_vector(12 downto 0);
signal sR_c0, sR_c1, sR_c2, sR_c3, sR_c4, sR_c5, sR_c6, sR_c7, sR_c8, sR_c9, sR_c10, sR_c11, sR_c12, sR_c13, sR_c14, sR_c15, sR_c16, sR_c17, sR_c18, sR_c19, sR_c20, sR_c21, sR_c22, sR_c23, sR_c24, sR_c25, sR_c26, sR_c27, sR_c28, sR_c29, sR_c30, sR_c31, sR_c32, sR_c33, sR_c34, sR_c35, sR_c36 :  std_logic;
signal exnXY_c0 :  std_logic_vector(3 downto 0);
signal exnR0_c0, exnR0_c1, exnR0_c2, exnR0_c3, exnR0_c4, exnR0_c5, exnR0_c6, exnR0_c7, exnR0_c8, exnR0_c9, exnR0_c10, exnR0_c11, exnR0_c12, exnR0_c13, exnR0_c14, exnR0_c15, exnR0_c16, exnR0_c17, exnR0_c18, exnR0_c19, exnR0_c20, exnR0_c21, exnR0_c22, exnR0_c23, exnR0_c24, exnR0_c25, exnR0_c26, exnR0_c27, exnR0_c28, exnR0_c29, exnR0_c30, exnR0_c31, exnR0_c32, exnR0_c33, exnR0_c34, exnR0_c35, exnR0_c36 :  std_logic_vector(1 downto 0);
signal D_c0, D_c1, D_c2, D_c3, D_c4, D_c5, D_c6, D_c7, D_c8, D_c9, D_c10, D_c11, D_c12, D_c13, D_c14, D_c15, D_c16, D_c17, D_c18, D_c19, D_c20, D_c21, D_c22, D_c23, D_c24, D_c25, D_c26, D_c27, D_c28, D_c29, D_c30, D_c31, D_c32, D_c33 :  std_logic_vector(52 downto 0);
signal psX_c0 :  std_logic_vector(53 downto 0);
signal betaw28_c0, betaw28_c1 :  std_logic_vector(55 downto 0);
signal sel28_c0 :  std_logic_vector(8 downto 0);
signal q28_c0, q28_c1 :  std_logic_vector(2 downto 0);
signal q28_copy5_c0 :  std_logic_vector(2 downto 0);
signal absq28D_c0, absq28D_c1 :  std_logic_vector(55 downto 0);
signal w27_c1 :  std_logic_vector(55 downto 0);
signal betaw27_c1, betaw27_c2 :  std_logic_vector(55 downto 0);
signal sel27_c1 :  std_logic_vector(8 downto 0);
signal q27_c1, q27_c2 :  std_logic_vector(2 downto 0);
signal q27_copy6_c1 :  std_logic_vector(2 downto 0);
signal absq27D_c1, absq27D_c2 :  std_logic_vector(55 downto 0);
signal w26_c2 :  std_logic_vector(55 downto 0);
signal betaw26_c2, betaw26_c3 :  std_logic_vector(55 downto 0);
signal sel26_c2 :  std_logic_vector(8 downto 0);
signal q26_c2, q26_c3 :  std_logic_vector(2 downto 0);
signal q26_copy7_c2 :  std_logic_vector(2 downto 0);
signal absq26D_c2, absq26D_c3 :  std_logic_vector(55 downto 0);
signal w25_c3 :  std_logic_vector(55 downto 0);
signal betaw25_c3, betaw25_c4 :  std_logic_vector(55 downto 0);
signal sel25_c3 :  std_logic_vector(8 downto 0);
signal q25_c4 :  std_logic_vector(2 downto 0);
signal q25_copy8_c3, q25_copy8_c4 :  std_logic_vector(2 downto 0);
signal absq25D_c4 :  std_logic_vector(55 downto 0);
signal w24_c4 :  std_logic_vector(55 downto 0);
signal betaw24_c4, betaw24_c5, betaw24_c6 :  std_logic_vector(55 downto 0);
signal sel24_c4 :  std_logic_vector(8 downto 0);
signal q24_c5, q24_c6 :  std_logic_vector(2 downto 0);
signal q24_copy9_c4, q24_copy9_c5 :  std_logic_vector(2 downto 0);
signal absq24D_c5, absq24D_c6 :  std_logic_vector(55 downto 0);
signal w23_c6 :  std_logic_vector(55 downto 0);
signal betaw23_c6, betaw23_c7 :  std_logic_vector(55 downto 0);
signal sel23_c6 :  std_logic_vector(8 downto 0);
signal q23_c6, q23_c7 :  std_logic_vector(2 downto 0);
signal q23_copy10_c6 :  std_logic_vector(2 downto 0);
signal absq23D_c6, absq23D_c7 :  std_logic_vector(55 downto 0);
signal w22_c7 :  std_logic_vector(55 downto 0);
signal betaw22_c7, betaw22_c8 :  std_logic_vector(55 downto 0);
signal sel22_c7 :  std_logic_vector(8 downto 0);
signal q22_c7, q22_c8 :  std_logic_vector(2 downto 0);
signal q22_copy11_c7 :  std_logic_vector(2 downto 0);
signal absq22D_c7, absq22D_c8 :  std_logic_vector(55 downto 0);
signal w21_c8 :  std_logic_vector(55 downto 0);
signal betaw21_c8, betaw21_c9 :  std_logic_vector(55 downto 0);
signal sel21_c8 :  std_logic_vector(8 downto 0);
signal q21_c9 :  std_logic_vector(2 downto 0);
signal q21_copy12_c8, q21_copy12_c9 :  std_logic_vector(2 downto 0);
signal absq21D_c9 :  std_logic_vector(55 downto 0);
signal w20_c9 :  std_logic_vector(55 downto 0);
signal betaw20_c9, betaw20_c10, betaw20_c11 :  std_logic_vector(55 downto 0);
signal sel20_c9 :  std_logic_vector(8 downto 0);
signal q20_c10, q20_c11 :  std_logic_vector(2 downto 0);
signal q20_copy13_c9, q20_copy13_c10 :  std_logic_vector(2 downto 0);
signal absq20D_c10, absq20D_c11 :  std_logic_vector(55 downto 0);
signal w19_c11 :  std_logic_vector(55 downto 0);
signal betaw19_c11, betaw19_c12 :  std_logic_vector(55 downto 0);
signal sel19_c11 :  std_logic_vector(8 downto 0);
signal q19_c11, q19_c12 :  std_logic_vector(2 downto 0);
signal q19_copy14_c11 :  std_logic_vector(2 downto 0);
signal absq19D_c11, absq19D_c12 :  std_logic_vector(55 downto 0);
signal w18_c12 :  std_logic_vector(55 downto 0);
signal betaw18_c12, betaw18_c13 :  std_logic_vector(55 downto 0);
signal sel18_c12 :  std_logic_vector(8 downto 0);
signal q18_c12, q18_c13 :  std_logic_vector(2 downto 0);
signal q18_copy15_c12 :  std_logic_vector(2 downto 0);
signal absq18D_c12, absq18D_c13 :  std_logic_vector(55 downto 0);
signal w17_c13 :  std_logic_vector(55 downto 0);
signal betaw17_c13, betaw17_c14 :  std_logic_vector(55 downto 0);
signal sel17_c13 :  std_logic_vector(8 downto 0);
signal q17_c14 :  std_logic_vector(2 downto 0);
signal q17_copy16_c13, q17_copy16_c14 :  std_logic_vector(2 downto 0);
signal absq17D_c14 :  std_logic_vector(55 downto 0);
signal w16_c14 :  std_logic_vector(55 downto 0);
signal betaw16_c14, betaw16_c15, betaw16_c16 :  std_logic_vector(55 downto 0);
signal sel16_c14 :  std_logic_vector(8 downto 0);
signal q16_c15, q16_c16 :  std_logic_vector(2 downto 0);
signal q16_copy17_c14, q16_copy17_c15 :  std_logic_vector(2 downto 0);
signal absq16D_c15, absq16D_c16 :  std_logic_vector(55 downto 0);
signal w15_c16 :  std_logic_vector(55 downto 0);
signal betaw15_c16, betaw15_c17 :  std_logic_vector(55 downto 0);
signal sel15_c16 :  std_logic_vector(8 downto 0);
signal q15_c16, q15_c17 :  std_logic_vector(2 downto 0);
signal q15_copy18_c16 :  std_logic_vector(2 downto 0);
signal absq15D_c16, absq15D_c17 :  std_logic_vector(55 downto 0);
signal w14_c17 :  std_logic_vector(55 downto 0);
signal betaw14_c17, betaw14_c18 :  std_logic_vector(55 downto 0);
signal sel14_c17 :  std_logic_vector(8 downto 0);
signal q14_c17, q14_c18 :  std_logic_vector(2 downto 0);
signal q14_copy19_c17 :  std_logic_vector(2 downto 0);
signal absq14D_c17, absq14D_c18 :  std_logic_vector(55 downto 0);
signal w13_c18 :  std_logic_vector(55 downto 0);
signal betaw13_c18, betaw13_c19 :  std_logic_vector(55 downto 0);
signal sel13_c18 :  std_logic_vector(8 downto 0);
signal q13_c18, q13_c19 :  std_logic_vector(2 downto 0);
signal q13_copy20_c18 :  std_logic_vector(2 downto 0);
signal absq13D_c18, absq13D_c19 :  std_logic_vector(55 downto 0);
signal w12_c19 :  std_logic_vector(55 downto 0);
signal betaw12_c19, betaw12_c20, betaw12_c21 :  std_logic_vector(55 downto 0);
signal sel12_c19 :  std_logic_vector(8 downto 0);
signal q12_c20, q12_c21 :  std_logic_vector(2 downto 0);
signal q12_copy21_c19, q12_copy21_c20 :  std_logic_vector(2 downto 0);
signal absq12D_c20, absq12D_c21 :  std_logic_vector(55 downto 0);
signal w11_c21 :  std_logic_vector(55 downto 0);
signal betaw11_c21, betaw11_c22 :  std_logic_vector(55 downto 0);
signal sel11_c21 :  std_logic_vector(8 downto 0);
signal q11_c21, q11_c22 :  std_logic_vector(2 downto 0);
signal q11_copy22_c21 :  std_logic_vector(2 downto 0);
signal absq11D_c21, absq11D_c22 :  std_logic_vector(55 downto 0);
signal w10_c22 :  std_logic_vector(55 downto 0);
signal betaw10_c22, betaw10_c23 :  std_logic_vector(55 downto 0);
signal sel10_c22 :  std_logic_vector(8 downto 0);
signal q10_c22, q10_c23 :  std_logic_vector(2 downto 0);
signal q10_copy23_c22 :  std_logic_vector(2 downto 0);
signal absq10D_c22, absq10D_c23 :  std_logic_vector(55 downto 0);
signal w9_c23 :  std_logic_vector(55 downto 0);
signal betaw9_c23, betaw9_c24 :  std_logic_vector(55 downto 0);
signal sel9_c23 :  std_logic_vector(8 downto 0);
signal q9_c23, q9_c24 :  std_logic_vector(2 downto 0);
signal q9_copy24_c23 :  std_logic_vector(2 downto 0);
signal absq9D_c23, absq9D_c24 :  std_logic_vector(55 downto 0);
signal w8_c24 :  std_logic_vector(55 downto 0);
signal betaw8_c24, betaw8_c25, betaw8_c26 :  std_logic_vector(55 downto 0);
signal sel8_c24 :  std_logic_vector(8 downto 0);
signal q8_c25, q8_c26 :  std_logic_vector(2 downto 0);
signal q8_copy25_c24, q8_copy25_c25 :  std_logic_vector(2 downto 0);
signal absq8D_c25, absq8D_c26 :  std_logic_vector(55 downto 0);
signal w7_c26 :  std_logic_vector(55 downto 0);
signal betaw7_c26, betaw7_c27 :  std_logic_vector(55 downto 0);
signal sel7_c26 :  std_logic_vector(8 downto 0);
signal q7_c26, q7_c27 :  std_logic_vector(2 downto 0);
signal q7_copy26_c26 :  std_logic_vector(2 downto 0);
signal absq7D_c26, absq7D_c27 :  std_logic_vector(55 downto 0);
signal w6_c27 :  std_logic_vector(55 downto 0);
signal betaw6_c27, betaw6_c28 :  std_logic_vector(55 downto 0);
signal sel6_c27 :  std_logic_vector(8 downto 0);
signal q6_c27, q6_c28 :  std_logic_vector(2 downto 0);
signal q6_copy27_c27 :  std_logic_vector(2 downto 0);
signal absq6D_c27, absq6D_c28 :  std_logic_vector(55 downto 0);
signal w5_c28 :  std_logic_vector(55 downto 0);
signal betaw5_c28, betaw5_c29 :  std_logic_vector(55 downto 0);
signal sel5_c28 :  std_logic_vector(8 downto 0);
signal q5_c28, q5_c29 :  std_logic_vector(2 downto 0);
signal q5_copy28_c28 :  std_logic_vector(2 downto 0);
signal absq5D_c28, absq5D_c29 :  std_logic_vector(55 downto 0);
signal w4_c29 :  std_logic_vector(55 downto 0);
signal betaw4_c29, betaw4_c30, betaw4_c31 :  std_logic_vector(55 downto 0);
signal sel4_c29 :  std_logic_vector(8 downto 0);
signal q4_c30, q4_c31 :  std_logic_vector(2 downto 0);
signal q4_copy29_c29, q4_copy29_c30 :  std_logic_vector(2 downto 0);
signal absq4D_c30, absq4D_c31 :  std_logic_vector(55 downto 0);
signal w3_c31 :  std_logic_vector(55 downto 0);
signal betaw3_c31, betaw3_c32 :  std_logic_vector(55 downto 0);
signal sel3_c31 :  std_logic_vector(8 downto 0);
signal q3_c31, q3_c32 :  std_logic_vector(2 downto 0);
signal q3_copy30_c31 :  std_logic_vector(2 downto 0);
signal absq3D_c31, absq3D_c32 :  std_logic_vector(55 downto 0);
signal w2_c32 :  std_logic_vector(55 downto 0);
signal betaw2_c32, betaw2_c33 :  std_logic_vector(55 downto 0);
signal sel2_c32 :  std_logic_vector(8 downto 0);
signal q2_c32, q2_c33 :  std_logic_vector(2 downto 0);
signal q2_copy31_c32 :  std_logic_vector(2 downto 0);
signal absq2D_c32, absq2D_c33 :  std_logic_vector(55 downto 0);
signal w1_c33 :  std_logic_vector(55 downto 0);
signal betaw1_c33, betaw1_c34 :  std_logic_vector(55 downto 0);
signal sel1_c33 :  std_logic_vector(8 downto 0);
signal q1_c33, q1_c34 :  std_logic_vector(2 downto 0);
signal q1_copy32_c33 :  std_logic_vector(2 downto 0);
signal absq1D_c33, absq1D_c34 :  std_logic_vector(55 downto 0);
signal w0_c34 :  std_logic_vector(55 downto 0);
signal wfinal_c34 :  std_logic_vector(53 downto 0);
signal qM0_c34 :  std_logic;
signal qP28_c0, qP28_c1, qP28_c2, qP28_c3, qP28_c4, qP28_c5, qP28_c6, qP28_c7, qP28_c8, qP28_c9, qP28_c10, qP28_c11, qP28_c12, qP28_c13, qP28_c14, qP28_c15, qP28_c16, qP28_c17, qP28_c18, qP28_c19, qP28_c20, qP28_c21, qP28_c22, qP28_c23, qP28_c24, qP28_c25, qP28_c26, qP28_c27, qP28_c28, qP28_c29, qP28_c30, qP28_c31, qP28_c32, qP28_c33 :  std_logic_vector(1 downto 0);
signal qM28_c0, qM28_c1, qM28_c2, qM28_c3, qM28_c4, qM28_c5, qM28_c6, qM28_c7, qM28_c8, qM28_c9, qM28_c10, qM28_c11, qM28_c12, qM28_c13, qM28_c14, qM28_c15, qM28_c16, qM28_c17, qM28_c18, qM28_c19, qM28_c20, qM28_c21, qM28_c22, qM28_c23, qM28_c24, qM28_c25, qM28_c26, qM28_c27, qM28_c28, qM28_c29, qM28_c30, qM28_c31, qM28_c32, qM28_c33, qM28_c34 :  std_logic_vector(1 downto 0);
signal qP27_c1, qP27_c2, qP27_c3, qP27_c4, qP27_c5, qP27_c6, qP27_c7, qP27_c8, qP27_c9, qP27_c10, qP27_c11, qP27_c12, qP27_c13, qP27_c14, qP27_c15, qP27_c16, qP27_c17, qP27_c18, qP27_c19, qP27_c20, qP27_c21, qP27_c22, qP27_c23, qP27_c24, qP27_c25, qP27_c26, qP27_c27, qP27_c28, qP27_c29, qP27_c30, qP27_c31, qP27_c32, qP27_c33 :  std_logic_vector(1 downto 0);
signal qM27_c1, qM27_c2, qM27_c3, qM27_c4, qM27_c5, qM27_c6, qM27_c7, qM27_c8, qM27_c9, qM27_c10, qM27_c11, qM27_c12, qM27_c13, qM27_c14, qM27_c15, qM27_c16, qM27_c17, qM27_c18, qM27_c19, qM27_c20, qM27_c21, qM27_c22, qM27_c23, qM27_c24, qM27_c25, qM27_c26, qM27_c27, qM27_c28, qM27_c29, qM27_c30, qM27_c31, qM27_c32, qM27_c33, qM27_c34 :  std_logic_vector(1 downto 0);
signal qP26_c2, qP26_c3, qP26_c4, qP26_c5, qP26_c6, qP26_c7, qP26_c8, qP26_c9, qP26_c10, qP26_c11, qP26_c12, qP26_c13, qP26_c14, qP26_c15, qP26_c16, qP26_c17, qP26_c18, qP26_c19, qP26_c20, qP26_c21, qP26_c22, qP26_c23, qP26_c24, qP26_c25, qP26_c26, qP26_c27, qP26_c28, qP26_c29, qP26_c30, qP26_c31, qP26_c32, qP26_c33 :  std_logic_vector(1 downto 0);
signal qM26_c2, qM26_c3, qM26_c4, qM26_c5, qM26_c6, qM26_c7, qM26_c8, qM26_c9, qM26_c10, qM26_c11, qM26_c12, qM26_c13, qM26_c14, qM26_c15, qM26_c16, qM26_c17, qM26_c18, qM26_c19, qM26_c20, qM26_c21, qM26_c22, qM26_c23, qM26_c24, qM26_c25, qM26_c26, qM26_c27, qM26_c28, qM26_c29, qM26_c30, qM26_c31, qM26_c32, qM26_c33, qM26_c34 :  std_logic_vector(1 downto 0);
signal qP25_c4, qP25_c5, qP25_c6, qP25_c7, qP25_c8, qP25_c9, qP25_c10, qP25_c11, qP25_c12, qP25_c13, qP25_c14, qP25_c15, qP25_c16, qP25_c17, qP25_c18, qP25_c19, qP25_c20, qP25_c21, qP25_c22, qP25_c23, qP25_c24, qP25_c25, qP25_c26, qP25_c27, qP25_c28, qP25_c29, qP25_c30, qP25_c31, qP25_c32, qP25_c33 :  std_logic_vector(1 downto 0);
signal qM25_c4, qM25_c5, qM25_c6, qM25_c7, qM25_c8, qM25_c9, qM25_c10, qM25_c11, qM25_c12, qM25_c13, qM25_c14, qM25_c15, qM25_c16, qM25_c17, qM25_c18, qM25_c19, qM25_c20, qM25_c21, qM25_c22, qM25_c23, qM25_c24, qM25_c25, qM25_c26, qM25_c27, qM25_c28, qM25_c29, qM25_c30, qM25_c31, qM25_c32, qM25_c33, qM25_c34 :  std_logic_vector(1 downto 0);
signal qP24_c5, qP24_c6, qP24_c7, qP24_c8, qP24_c9, qP24_c10, qP24_c11, qP24_c12, qP24_c13, qP24_c14, qP24_c15, qP24_c16, qP24_c17, qP24_c18, qP24_c19, qP24_c20, qP24_c21, qP24_c22, qP24_c23, qP24_c24, qP24_c25, qP24_c26, qP24_c27, qP24_c28, qP24_c29, qP24_c30, qP24_c31, qP24_c32, qP24_c33 :  std_logic_vector(1 downto 0);
signal qM24_c5, qM24_c6, qM24_c7, qM24_c8, qM24_c9, qM24_c10, qM24_c11, qM24_c12, qM24_c13, qM24_c14, qM24_c15, qM24_c16, qM24_c17, qM24_c18, qM24_c19, qM24_c20, qM24_c21, qM24_c22, qM24_c23, qM24_c24, qM24_c25, qM24_c26, qM24_c27, qM24_c28, qM24_c29, qM24_c30, qM24_c31, qM24_c32, qM24_c33, qM24_c34 :  std_logic_vector(1 downto 0);
signal qP23_c6, qP23_c7, qP23_c8, qP23_c9, qP23_c10, qP23_c11, qP23_c12, qP23_c13, qP23_c14, qP23_c15, qP23_c16, qP23_c17, qP23_c18, qP23_c19, qP23_c20, qP23_c21, qP23_c22, qP23_c23, qP23_c24, qP23_c25, qP23_c26, qP23_c27, qP23_c28, qP23_c29, qP23_c30, qP23_c31, qP23_c32, qP23_c33 :  std_logic_vector(1 downto 0);
signal qM23_c6, qM23_c7, qM23_c8, qM23_c9, qM23_c10, qM23_c11, qM23_c12, qM23_c13, qM23_c14, qM23_c15, qM23_c16, qM23_c17, qM23_c18, qM23_c19, qM23_c20, qM23_c21, qM23_c22, qM23_c23, qM23_c24, qM23_c25, qM23_c26, qM23_c27, qM23_c28, qM23_c29, qM23_c30, qM23_c31, qM23_c32, qM23_c33, qM23_c34 :  std_logic_vector(1 downto 0);
signal qP22_c7, qP22_c8, qP22_c9, qP22_c10, qP22_c11, qP22_c12, qP22_c13, qP22_c14, qP22_c15, qP22_c16, qP22_c17, qP22_c18, qP22_c19, qP22_c20, qP22_c21, qP22_c22, qP22_c23, qP22_c24, qP22_c25, qP22_c26, qP22_c27, qP22_c28, qP22_c29, qP22_c30, qP22_c31, qP22_c32, qP22_c33 :  std_logic_vector(1 downto 0);
signal qM22_c7, qM22_c8, qM22_c9, qM22_c10, qM22_c11, qM22_c12, qM22_c13, qM22_c14, qM22_c15, qM22_c16, qM22_c17, qM22_c18, qM22_c19, qM22_c20, qM22_c21, qM22_c22, qM22_c23, qM22_c24, qM22_c25, qM22_c26, qM22_c27, qM22_c28, qM22_c29, qM22_c30, qM22_c31, qM22_c32, qM22_c33, qM22_c34 :  std_logic_vector(1 downto 0);
signal qP21_c9, qP21_c10, qP21_c11, qP21_c12, qP21_c13, qP21_c14, qP21_c15, qP21_c16, qP21_c17, qP21_c18, qP21_c19, qP21_c20, qP21_c21, qP21_c22, qP21_c23, qP21_c24, qP21_c25, qP21_c26, qP21_c27, qP21_c28, qP21_c29, qP21_c30, qP21_c31, qP21_c32, qP21_c33 :  std_logic_vector(1 downto 0);
signal qM21_c9, qM21_c10, qM21_c11, qM21_c12, qM21_c13, qM21_c14, qM21_c15, qM21_c16, qM21_c17, qM21_c18, qM21_c19, qM21_c20, qM21_c21, qM21_c22, qM21_c23, qM21_c24, qM21_c25, qM21_c26, qM21_c27, qM21_c28, qM21_c29, qM21_c30, qM21_c31, qM21_c32, qM21_c33, qM21_c34 :  std_logic_vector(1 downto 0);
signal qP20_c10, qP20_c11, qP20_c12, qP20_c13, qP20_c14, qP20_c15, qP20_c16, qP20_c17, qP20_c18, qP20_c19, qP20_c20, qP20_c21, qP20_c22, qP20_c23, qP20_c24, qP20_c25, qP20_c26, qP20_c27, qP20_c28, qP20_c29, qP20_c30, qP20_c31, qP20_c32, qP20_c33 :  std_logic_vector(1 downto 0);
signal qM20_c10, qM20_c11, qM20_c12, qM20_c13, qM20_c14, qM20_c15, qM20_c16, qM20_c17, qM20_c18, qM20_c19, qM20_c20, qM20_c21, qM20_c22, qM20_c23, qM20_c24, qM20_c25, qM20_c26, qM20_c27, qM20_c28, qM20_c29, qM20_c30, qM20_c31, qM20_c32, qM20_c33, qM20_c34 :  std_logic_vector(1 downto 0);
signal qP19_c11, qP19_c12, qP19_c13, qP19_c14, qP19_c15, qP19_c16, qP19_c17, qP19_c18, qP19_c19, qP19_c20, qP19_c21, qP19_c22, qP19_c23, qP19_c24, qP19_c25, qP19_c26, qP19_c27, qP19_c28, qP19_c29, qP19_c30, qP19_c31, qP19_c32, qP19_c33 :  std_logic_vector(1 downto 0);
signal qM19_c11, qM19_c12, qM19_c13, qM19_c14, qM19_c15, qM19_c16, qM19_c17, qM19_c18, qM19_c19, qM19_c20, qM19_c21, qM19_c22, qM19_c23, qM19_c24, qM19_c25, qM19_c26, qM19_c27, qM19_c28, qM19_c29, qM19_c30, qM19_c31, qM19_c32, qM19_c33, qM19_c34 :  std_logic_vector(1 downto 0);
signal qP18_c12, qP18_c13, qP18_c14, qP18_c15, qP18_c16, qP18_c17, qP18_c18, qP18_c19, qP18_c20, qP18_c21, qP18_c22, qP18_c23, qP18_c24, qP18_c25, qP18_c26, qP18_c27, qP18_c28, qP18_c29, qP18_c30, qP18_c31, qP18_c32, qP18_c33 :  std_logic_vector(1 downto 0);
signal qM18_c12, qM18_c13, qM18_c14, qM18_c15, qM18_c16, qM18_c17, qM18_c18, qM18_c19, qM18_c20, qM18_c21, qM18_c22, qM18_c23, qM18_c24, qM18_c25, qM18_c26, qM18_c27, qM18_c28, qM18_c29, qM18_c30, qM18_c31, qM18_c32, qM18_c33, qM18_c34 :  std_logic_vector(1 downto 0);
signal qP17_c14, qP17_c15, qP17_c16, qP17_c17, qP17_c18, qP17_c19, qP17_c20, qP17_c21, qP17_c22, qP17_c23, qP17_c24, qP17_c25, qP17_c26, qP17_c27, qP17_c28, qP17_c29, qP17_c30, qP17_c31, qP17_c32, qP17_c33 :  std_logic_vector(1 downto 0);
signal qM17_c14, qM17_c15, qM17_c16, qM17_c17, qM17_c18, qM17_c19, qM17_c20, qM17_c21, qM17_c22, qM17_c23, qM17_c24, qM17_c25, qM17_c26, qM17_c27, qM17_c28, qM17_c29, qM17_c30, qM17_c31, qM17_c32, qM17_c33, qM17_c34 :  std_logic_vector(1 downto 0);
signal qP16_c15, qP16_c16, qP16_c17, qP16_c18, qP16_c19, qP16_c20, qP16_c21, qP16_c22, qP16_c23, qP16_c24, qP16_c25, qP16_c26, qP16_c27, qP16_c28, qP16_c29, qP16_c30, qP16_c31, qP16_c32, qP16_c33 :  std_logic_vector(1 downto 0);
signal qM16_c15, qM16_c16, qM16_c17, qM16_c18, qM16_c19, qM16_c20, qM16_c21, qM16_c22, qM16_c23, qM16_c24, qM16_c25, qM16_c26, qM16_c27, qM16_c28, qM16_c29, qM16_c30, qM16_c31, qM16_c32, qM16_c33, qM16_c34 :  std_logic_vector(1 downto 0);
signal qP15_c16, qP15_c17, qP15_c18, qP15_c19, qP15_c20, qP15_c21, qP15_c22, qP15_c23, qP15_c24, qP15_c25, qP15_c26, qP15_c27, qP15_c28, qP15_c29, qP15_c30, qP15_c31, qP15_c32, qP15_c33 :  std_logic_vector(1 downto 0);
signal qM15_c16, qM15_c17, qM15_c18, qM15_c19, qM15_c20, qM15_c21, qM15_c22, qM15_c23, qM15_c24, qM15_c25, qM15_c26, qM15_c27, qM15_c28, qM15_c29, qM15_c30, qM15_c31, qM15_c32, qM15_c33, qM15_c34 :  std_logic_vector(1 downto 0);
signal qP14_c17, qP14_c18, qP14_c19, qP14_c20, qP14_c21, qP14_c22, qP14_c23, qP14_c24, qP14_c25, qP14_c26, qP14_c27, qP14_c28, qP14_c29, qP14_c30, qP14_c31, qP14_c32, qP14_c33 :  std_logic_vector(1 downto 0);
signal qM14_c17, qM14_c18, qM14_c19, qM14_c20, qM14_c21, qM14_c22, qM14_c23, qM14_c24, qM14_c25, qM14_c26, qM14_c27, qM14_c28, qM14_c29, qM14_c30, qM14_c31, qM14_c32, qM14_c33, qM14_c34 :  std_logic_vector(1 downto 0);
signal qP13_c18, qP13_c19, qP13_c20, qP13_c21, qP13_c22, qP13_c23, qP13_c24, qP13_c25, qP13_c26, qP13_c27, qP13_c28, qP13_c29, qP13_c30, qP13_c31, qP13_c32, qP13_c33 :  std_logic_vector(1 downto 0);
signal qM13_c18, qM13_c19, qM13_c20, qM13_c21, qM13_c22, qM13_c23, qM13_c24, qM13_c25, qM13_c26, qM13_c27, qM13_c28, qM13_c29, qM13_c30, qM13_c31, qM13_c32, qM13_c33, qM13_c34 :  std_logic_vector(1 downto 0);
signal qP12_c20, qP12_c21, qP12_c22, qP12_c23, qP12_c24, qP12_c25, qP12_c26, qP12_c27, qP12_c28, qP12_c29, qP12_c30, qP12_c31, qP12_c32, qP12_c33 :  std_logic_vector(1 downto 0);
signal qM12_c20, qM12_c21, qM12_c22, qM12_c23, qM12_c24, qM12_c25, qM12_c26, qM12_c27, qM12_c28, qM12_c29, qM12_c30, qM12_c31, qM12_c32, qM12_c33, qM12_c34 :  std_logic_vector(1 downto 0);
signal qP11_c21, qP11_c22, qP11_c23, qP11_c24, qP11_c25, qP11_c26, qP11_c27, qP11_c28, qP11_c29, qP11_c30, qP11_c31, qP11_c32, qP11_c33 :  std_logic_vector(1 downto 0);
signal qM11_c21, qM11_c22, qM11_c23, qM11_c24, qM11_c25, qM11_c26, qM11_c27, qM11_c28, qM11_c29, qM11_c30, qM11_c31, qM11_c32, qM11_c33, qM11_c34 :  std_logic_vector(1 downto 0);
signal qP10_c22, qP10_c23, qP10_c24, qP10_c25, qP10_c26, qP10_c27, qP10_c28, qP10_c29, qP10_c30, qP10_c31, qP10_c32, qP10_c33 :  std_logic_vector(1 downto 0);
signal qM10_c22, qM10_c23, qM10_c24, qM10_c25, qM10_c26, qM10_c27, qM10_c28, qM10_c29, qM10_c30, qM10_c31, qM10_c32, qM10_c33, qM10_c34 :  std_logic_vector(1 downto 0);
signal qP9_c23, qP9_c24, qP9_c25, qP9_c26, qP9_c27, qP9_c28, qP9_c29, qP9_c30, qP9_c31, qP9_c32, qP9_c33 :  std_logic_vector(1 downto 0);
signal qM9_c23, qM9_c24, qM9_c25, qM9_c26, qM9_c27, qM9_c28, qM9_c29, qM9_c30, qM9_c31, qM9_c32, qM9_c33, qM9_c34 :  std_logic_vector(1 downto 0);
signal qP8_c25, qP8_c26, qP8_c27, qP8_c28, qP8_c29, qP8_c30, qP8_c31, qP8_c32, qP8_c33 :  std_logic_vector(1 downto 0);
signal qM8_c25, qM8_c26, qM8_c27, qM8_c28, qM8_c29, qM8_c30, qM8_c31, qM8_c32, qM8_c33, qM8_c34 :  std_logic_vector(1 downto 0);
signal qP7_c26, qP7_c27, qP7_c28, qP7_c29, qP7_c30, qP7_c31, qP7_c32, qP7_c33 :  std_logic_vector(1 downto 0);
signal qM7_c26, qM7_c27, qM7_c28, qM7_c29, qM7_c30, qM7_c31, qM7_c32, qM7_c33, qM7_c34 :  std_logic_vector(1 downto 0);
signal qP6_c27, qP6_c28, qP6_c29, qP6_c30, qP6_c31, qP6_c32, qP6_c33 :  std_logic_vector(1 downto 0);
signal qM6_c27, qM6_c28, qM6_c29, qM6_c30, qM6_c31, qM6_c32, qM6_c33, qM6_c34 :  std_logic_vector(1 downto 0);
signal qP5_c28, qP5_c29, qP5_c30, qP5_c31, qP5_c32, qP5_c33 :  std_logic_vector(1 downto 0);
signal qM5_c28, qM5_c29, qM5_c30, qM5_c31, qM5_c32, qM5_c33, qM5_c34 :  std_logic_vector(1 downto 0);
signal qP4_c30, qP4_c31, qP4_c32, qP4_c33 :  std_logic_vector(1 downto 0);
signal qM4_c30, qM4_c31, qM4_c32, qM4_c33, qM4_c34 :  std_logic_vector(1 downto 0);
signal qP3_c31, qP3_c32, qP3_c33 :  std_logic_vector(1 downto 0);
signal qM3_c31, qM3_c32, qM3_c33, qM3_c34 :  std_logic_vector(1 downto 0);
signal qP2_c32, qP2_c33 :  std_logic_vector(1 downto 0);
signal qM2_c32, qM2_c33, qM2_c34 :  std_logic_vector(1 downto 0);
signal qP1_c33 :  std_logic_vector(1 downto 0);
signal qM1_c33, qM1_c34 :  std_logic_vector(1 downto 0);
signal qP_c33, qP_c34, qP_c35 :  std_logic_vector(55 downto 0);
signal qM_c34, qM_c35 :  std_logic_vector(55 downto 0);
signal quotient_c35 :  std_logic_vector(55 downto 0);
signal mR_c35, mR_c36 :  std_logic_vector(54 downto 0);
signal fRnorm_c35, fRnorm_c36 :  std_logic_vector(52 downto 0);
signal round_c35, round_c36 :  std_logic;
signal expR1_c36 :  std_logic_vector(12 downto 0);
signal expfrac_c36 :  std_logic_vector(64 downto 0);
signal expfracR_c36 :  std_logic_vector(64 downto 0);
signal exnR_c36 :  std_logic_vector(1 downto 0);
signal exnRfinal_c36 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               expR0_c1 <= expR0_c0;
               sR_c1 <= sR_c0;
               exnR0_c1 <= exnR0_c0;
               D_c1 <= D_c0;
               betaw28_c1 <= betaw28_c0;
               q28_c1 <= q28_c0;
               absq28D_c1 <= absq28D_c0;
               qP28_c1 <= qP28_c0;
               qM28_c1 <= qM28_c0;
            end if;
            if ce_2 = '1' then
               expR0_c2 <= expR0_c1;
               sR_c2 <= sR_c1;
               exnR0_c2 <= exnR0_c1;
               D_c2 <= D_c1;
               betaw27_c2 <= betaw27_c1;
               q27_c2 <= q27_c1;
               absq27D_c2 <= absq27D_c1;
               qP28_c2 <= qP28_c1;
               qM28_c2 <= qM28_c1;
               qP27_c2 <= qP27_c1;
               qM27_c2 <= qM27_c1;
            end if;
            if ce_3 = '1' then
               expR0_c3 <= expR0_c2;
               sR_c3 <= sR_c2;
               exnR0_c3 <= exnR0_c2;
               D_c3 <= D_c2;
               betaw26_c3 <= betaw26_c2;
               q26_c3 <= q26_c2;
               absq26D_c3 <= absq26D_c2;
               qP28_c3 <= qP28_c2;
               qM28_c3 <= qM28_c2;
               qP27_c3 <= qP27_c2;
               qM27_c3 <= qM27_c2;
               qP26_c3 <= qP26_c2;
               qM26_c3 <= qM26_c2;
            end if;
            if ce_4 = '1' then
               expR0_c4 <= expR0_c3;
               sR_c4 <= sR_c3;
               exnR0_c4 <= exnR0_c3;
               D_c4 <= D_c3;
               betaw25_c4 <= betaw25_c3;
               q25_copy8_c4 <= q25_copy8_c3;
               qP28_c4 <= qP28_c3;
               qM28_c4 <= qM28_c3;
               qP27_c4 <= qP27_c3;
               qM27_c4 <= qM27_c3;
               qP26_c4 <= qP26_c3;
               qM26_c4 <= qM26_c3;
            end if;
            if ce_5 = '1' then
               expR0_c5 <= expR0_c4;
               sR_c5 <= sR_c4;
               exnR0_c5 <= exnR0_c4;
               D_c5 <= D_c4;
               betaw24_c5 <= betaw24_c4;
               q24_copy9_c5 <= q24_copy9_c4;
               qP28_c5 <= qP28_c4;
               qM28_c5 <= qM28_c4;
               qP27_c5 <= qP27_c4;
               qM27_c5 <= qM27_c4;
               qP26_c5 <= qP26_c4;
               qM26_c5 <= qM26_c4;
               qP25_c5 <= qP25_c4;
               qM25_c5 <= qM25_c4;
            end if;
            if ce_6 = '1' then
               expR0_c6 <= expR0_c5;
               sR_c6 <= sR_c5;
               exnR0_c6 <= exnR0_c5;
               D_c6 <= D_c5;
               betaw24_c6 <= betaw24_c5;
               q24_c6 <= q24_c5;
               absq24D_c6 <= absq24D_c5;
               qP28_c6 <= qP28_c5;
               qM28_c6 <= qM28_c5;
               qP27_c6 <= qP27_c5;
               qM27_c6 <= qM27_c5;
               qP26_c6 <= qP26_c5;
               qM26_c6 <= qM26_c5;
               qP25_c6 <= qP25_c5;
               qM25_c6 <= qM25_c5;
               qP24_c6 <= qP24_c5;
               qM24_c6 <= qM24_c5;
            end if;
            if ce_7 = '1' then
               expR0_c7 <= expR0_c6;
               sR_c7 <= sR_c6;
               exnR0_c7 <= exnR0_c6;
               D_c7 <= D_c6;
               betaw23_c7 <= betaw23_c6;
               q23_c7 <= q23_c6;
               absq23D_c7 <= absq23D_c6;
               qP28_c7 <= qP28_c6;
               qM28_c7 <= qM28_c6;
               qP27_c7 <= qP27_c6;
               qM27_c7 <= qM27_c6;
               qP26_c7 <= qP26_c6;
               qM26_c7 <= qM26_c6;
               qP25_c7 <= qP25_c6;
               qM25_c7 <= qM25_c6;
               qP24_c7 <= qP24_c6;
               qM24_c7 <= qM24_c6;
               qP23_c7 <= qP23_c6;
               qM23_c7 <= qM23_c6;
            end if;
            if ce_8 = '1' then
               expR0_c8 <= expR0_c7;
               sR_c8 <= sR_c7;
               exnR0_c8 <= exnR0_c7;
               D_c8 <= D_c7;
               betaw22_c8 <= betaw22_c7;
               q22_c8 <= q22_c7;
               absq22D_c8 <= absq22D_c7;
               qP28_c8 <= qP28_c7;
               qM28_c8 <= qM28_c7;
               qP27_c8 <= qP27_c7;
               qM27_c8 <= qM27_c7;
               qP26_c8 <= qP26_c7;
               qM26_c8 <= qM26_c7;
               qP25_c8 <= qP25_c7;
               qM25_c8 <= qM25_c7;
               qP24_c8 <= qP24_c7;
               qM24_c8 <= qM24_c7;
               qP23_c8 <= qP23_c7;
               qM23_c8 <= qM23_c7;
               qP22_c8 <= qP22_c7;
               qM22_c8 <= qM22_c7;
            end if;
            if ce_9 = '1' then
               expR0_c9 <= expR0_c8;
               sR_c9 <= sR_c8;
               exnR0_c9 <= exnR0_c8;
               D_c9 <= D_c8;
               betaw21_c9 <= betaw21_c8;
               q21_copy12_c9 <= q21_copy12_c8;
               qP28_c9 <= qP28_c8;
               qM28_c9 <= qM28_c8;
               qP27_c9 <= qP27_c8;
               qM27_c9 <= qM27_c8;
               qP26_c9 <= qP26_c8;
               qM26_c9 <= qM26_c8;
               qP25_c9 <= qP25_c8;
               qM25_c9 <= qM25_c8;
               qP24_c9 <= qP24_c8;
               qM24_c9 <= qM24_c8;
               qP23_c9 <= qP23_c8;
               qM23_c9 <= qM23_c8;
               qP22_c9 <= qP22_c8;
               qM22_c9 <= qM22_c8;
            end if;
            if ce_10 = '1' then
               expR0_c10 <= expR0_c9;
               sR_c10 <= sR_c9;
               exnR0_c10 <= exnR0_c9;
               D_c10 <= D_c9;
               betaw20_c10 <= betaw20_c9;
               q20_copy13_c10 <= q20_copy13_c9;
               qP28_c10 <= qP28_c9;
               qM28_c10 <= qM28_c9;
               qP27_c10 <= qP27_c9;
               qM27_c10 <= qM27_c9;
               qP26_c10 <= qP26_c9;
               qM26_c10 <= qM26_c9;
               qP25_c10 <= qP25_c9;
               qM25_c10 <= qM25_c9;
               qP24_c10 <= qP24_c9;
               qM24_c10 <= qM24_c9;
               qP23_c10 <= qP23_c9;
               qM23_c10 <= qM23_c9;
               qP22_c10 <= qP22_c9;
               qM22_c10 <= qM22_c9;
               qP21_c10 <= qP21_c9;
               qM21_c10 <= qM21_c9;
            end if;
            if ce_11 = '1' then
               expR0_c11 <= expR0_c10;
               sR_c11 <= sR_c10;
               exnR0_c11 <= exnR0_c10;
               D_c11 <= D_c10;
               betaw20_c11 <= betaw20_c10;
               q20_c11 <= q20_c10;
               absq20D_c11 <= absq20D_c10;
               qP28_c11 <= qP28_c10;
               qM28_c11 <= qM28_c10;
               qP27_c11 <= qP27_c10;
               qM27_c11 <= qM27_c10;
               qP26_c11 <= qP26_c10;
               qM26_c11 <= qM26_c10;
               qP25_c11 <= qP25_c10;
               qM25_c11 <= qM25_c10;
               qP24_c11 <= qP24_c10;
               qM24_c11 <= qM24_c10;
               qP23_c11 <= qP23_c10;
               qM23_c11 <= qM23_c10;
               qP22_c11 <= qP22_c10;
               qM22_c11 <= qM22_c10;
               qP21_c11 <= qP21_c10;
               qM21_c11 <= qM21_c10;
               qP20_c11 <= qP20_c10;
               qM20_c11 <= qM20_c10;
            end if;
            if ce_12 = '1' then
               expR0_c12 <= expR0_c11;
               sR_c12 <= sR_c11;
               exnR0_c12 <= exnR0_c11;
               D_c12 <= D_c11;
               betaw19_c12 <= betaw19_c11;
               q19_c12 <= q19_c11;
               absq19D_c12 <= absq19D_c11;
               qP28_c12 <= qP28_c11;
               qM28_c12 <= qM28_c11;
               qP27_c12 <= qP27_c11;
               qM27_c12 <= qM27_c11;
               qP26_c12 <= qP26_c11;
               qM26_c12 <= qM26_c11;
               qP25_c12 <= qP25_c11;
               qM25_c12 <= qM25_c11;
               qP24_c12 <= qP24_c11;
               qM24_c12 <= qM24_c11;
               qP23_c12 <= qP23_c11;
               qM23_c12 <= qM23_c11;
               qP22_c12 <= qP22_c11;
               qM22_c12 <= qM22_c11;
               qP21_c12 <= qP21_c11;
               qM21_c12 <= qM21_c11;
               qP20_c12 <= qP20_c11;
               qM20_c12 <= qM20_c11;
               qP19_c12 <= qP19_c11;
               qM19_c12 <= qM19_c11;
            end if;
            if ce_13 = '1' then
               expR0_c13 <= expR0_c12;
               sR_c13 <= sR_c12;
               exnR0_c13 <= exnR0_c12;
               D_c13 <= D_c12;
               betaw18_c13 <= betaw18_c12;
               q18_c13 <= q18_c12;
               absq18D_c13 <= absq18D_c12;
               qP28_c13 <= qP28_c12;
               qM28_c13 <= qM28_c12;
               qP27_c13 <= qP27_c12;
               qM27_c13 <= qM27_c12;
               qP26_c13 <= qP26_c12;
               qM26_c13 <= qM26_c12;
               qP25_c13 <= qP25_c12;
               qM25_c13 <= qM25_c12;
               qP24_c13 <= qP24_c12;
               qM24_c13 <= qM24_c12;
               qP23_c13 <= qP23_c12;
               qM23_c13 <= qM23_c12;
               qP22_c13 <= qP22_c12;
               qM22_c13 <= qM22_c12;
               qP21_c13 <= qP21_c12;
               qM21_c13 <= qM21_c12;
               qP20_c13 <= qP20_c12;
               qM20_c13 <= qM20_c12;
               qP19_c13 <= qP19_c12;
               qM19_c13 <= qM19_c12;
               qP18_c13 <= qP18_c12;
               qM18_c13 <= qM18_c12;
            end if;
            if ce_14 = '1' then
               expR0_c14 <= expR0_c13;
               sR_c14 <= sR_c13;
               exnR0_c14 <= exnR0_c13;
               D_c14 <= D_c13;
               betaw17_c14 <= betaw17_c13;
               q17_copy16_c14 <= q17_copy16_c13;
               qP28_c14 <= qP28_c13;
               qM28_c14 <= qM28_c13;
               qP27_c14 <= qP27_c13;
               qM27_c14 <= qM27_c13;
               qP26_c14 <= qP26_c13;
               qM26_c14 <= qM26_c13;
               qP25_c14 <= qP25_c13;
               qM25_c14 <= qM25_c13;
               qP24_c14 <= qP24_c13;
               qM24_c14 <= qM24_c13;
               qP23_c14 <= qP23_c13;
               qM23_c14 <= qM23_c13;
               qP22_c14 <= qP22_c13;
               qM22_c14 <= qM22_c13;
               qP21_c14 <= qP21_c13;
               qM21_c14 <= qM21_c13;
               qP20_c14 <= qP20_c13;
               qM20_c14 <= qM20_c13;
               qP19_c14 <= qP19_c13;
               qM19_c14 <= qM19_c13;
               qP18_c14 <= qP18_c13;
               qM18_c14 <= qM18_c13;
            end if;
            if ce_15 = '1' then
               expR0_c15 <= expR0_c14;
               sR_c15 <= sR_c14;
               exnR0_c15 <= exnR0_c14;
               D_c15 <= D_c14;
               betaw16_c15 <= betaw16_c14;
               q16_copy17_c15 <= q16_copy17_c14;
               qP28_c15 <= qP28_c14;
               qM28_c15 <= qM28_c14;
               qP27_c15 <= qP27_c14;
               qM27_c15 <= qM27_c14;
               qP26_c15 <= qP26_c14;
               qM26_c15 <= qM26_c14;
               qP25_c15 <= qP25_c14;
               qM25_c15 <= qM25_c14;
               qP24_c15 <= qP24_c14;
               qM24_c15 <= qM24_c14;
               qP23_c15 <= qP23_c14;
               qM23_c15 <= qM23_c14;
               qP22_c15 <= qP22_c14;
               qM22_c15 <= qM22_c14;
               qP21_c15 <= qP21_c14;
               qM21_c15 <= qM21_c14;
               qP20_c15 <= qP20_c14;
               qM20_c15 <= qM20_c14;
               qP19_c15 <= qP19_c14;
               qM19_c15 <= qM19_c14;
               qP18_c15 <= qP18_c14;
               qM18_c15 <= qM18_c14;
               qP17_c15 <= qP17_c14;
               qM17_c15 <= qM17_c14;
            end if;
            if ce_16 = '1' then
               expR0_c16 <= expR0_c15;
               sR_c16 <= sR_c15;
               exnR0_c16 <= exnR0_c15;
               D_c16 <= D_c15;
               betaw16_c16 <= betaw16_c15;
               q16_c16 <= q16_c15;
               absq16D_c16 <= absq16D_c15;
               qP28_c16 <= qP28_c15;
               qM28_c16 <= qM28_c15;
               qP27_c16 <= qP27_c15;
               qM27_c16 <= qM27_c15;
               qP26_c16 <= qP26_c15;
               qM26_c16 <= qM26_c15;
               qP25_c16 <= qP25_c15;
               qM25_c16 <= qM25_c15;
               qP24_c16 <= qP24_c15;
               qM24_c16 <= qM24_c15;
               qP23_c16 <= qP23_c15;
               qM23_c16 <= qM23_c15;
               qP22_c16 <= qP22_c15;
               qM22_c16 <= qM22_c15;
               qP21_c16 <= qP21_c15;
               qM21_c16 <= qM21_c15;
               qP20_c16 <= qP20_c15;
               qM20_c16 <= qM20_c15;
               qP19_c16 <= qP19_c15;
               qM19_c16 <= qM19_c15;
               qP18_c16 <= qP18_c15;
               qM18_c16 <= qM18_c15;
               qP17_c16 <= qP17_c15;
               qM17_c16 <= qM17_c15;
               qP16_c16 <= qP16_c15;
               qM16_c16 <= qM16_c15;
            end if;
            if ce_17 = '1' then
               expR0_c17 <= expR0_c16;
               sR_c17 <= sR_c16;
               exnR0_c17 <= exnR0_c16;
               D_c17 <= D_c16;
               betaw15_c17 <= betaw15_c16;
               q15_c17 <= q15_c16;
               absq15D_c17 <= absq15D_c16;
               qP28_c17 <= qP28_c16;
               qM28_c17 <= qM28_c16;
               qP27_c17 <= qP27_c16;
               qM27_c17 <= qM27_c16;
               qP26_c17 <= qP26_c16;
               qM26_c17 <= qM26_c16;
               qP25_c17 <= qP25_c16;
               qM25_c17 <= qM25_c16;
               qP24_c17 <= qP24_c16;
               qM24_c17 <= qM24_c16;
               qP23_c17 <= qP23_c16;
               qM23_c17 <= qM23_c16;
               qP22_c17 <= qP22_c16;
               qM22_c17 <= qM22_c16;
               qP21_c17 <= qP21_c16;
               qM21_c17 <= qM21_c16;
               qP20_c17 <= qP20_c16;
               qM20_c17 <= qM20_c16;
               qP19_c17 <= qP19_c16;
               qM19_c17 <= qM19_c16;
               qP18_c17 <= qP18_c16;
               qM18_c17 <= qM18_c16;
               qP17_c17 <= qP17_c16;
               qM17_c17 <= qM17_c16;
               qP16_c17 <= qP16_c16;
               qM16_c17 <= qM16_c16;
               qP15_c17 <= qP15_c16;
               qM15_c17 <= qM15_c16;
            end if;
            if ce_18 = '1' then
               expR0_c18 <= expR0_c17;
               sR_c18 <= sR_c17;
               exnR0_c18 <= exnR0_c17;
               D_c18 <= D_c17;
               betaw14_c18 <= betaw14_c17;
               q14_c18 <= q14_c17;
               absq14D_c18 <= absq14D_c17;
               qP28_c18 <= qP28_c17;
               qM28_c18 <= qM28_c17;
               qP27_c18 <= qP27_c17;
               qM27_c18 <= qM27_c17;
               qP26_c18 <= qP26_c17;
               qM26_c18 <= qM26_c17;
               qP25_c18 <= qP25_c17;
               qM25_c18 <= qM25_c17;
               qP24_c18 <= qP24_c17;
               qM24_c18 <= qM24_c17;
               qP23_c18 <= qP23_c17;
               qM23_c18 <= qM23_c17;
               qP22_c18 <= qP22_c17;
               qM22_c18 <= qM22_c17;
               qP21_c18 <= qP21_c17;
               qM21_c18 <= qM21_c17;
               qP20_c18 <= qP20_c17;
               qM20_c18 <= qM20_c17;
               qP19_c18 <= qP19_c17;
               qM19_c18 <= qM19_c17;
               qP18_c18 <= qP18_c17;
               qM18_c18 <= qM18_c17;
               qP17_c18 <= qP17_c17;
               qM17_c18 <= qM17_c17;
               qP16_c18 <= qP16_c17;
               qM16_c18 <= qM16_c17;
               qP15_c18 <= qP15_c17;
               qM15_c18 <= qM15_c17;
               qP14_c18 <= qP14_c17;
               qM14_c18 <= qM14_c17;
            end if;
            if ce_19 = '1' then
               expR0_c19 <= expR0_c18;
               sR_c19 <= sR_c18;
               exnR0_c19 <= exnR0_c18;
               D_c19 <= D_c18;
               betaw13_c19 <= betaw13_c18;
               q13_c19 <= q13_c18;
               absq13D_c19 <= absq13D_c18;
               qP28_c19 <= qP28_c18;
               qM28_c19 <= qM28_c18;
               qP27_c19 <= qP27_c18;
               qM27_c19 <= qM27_c18;
               qP26_c19 <= qP26_c18;
               qM26_c19 <= qM26_c18;
               qP25_c19 <= qP25_c18;
               qM25_c19 <= qM25_c18;
               qP24_c19 <= qP24_c18;
               qM24_c19 <= qM24_c18;
               qP23_c19 <= qP23_c18;
               qM23_c19 <= qM23_c18;
               qP22_c19 <= qP22_c18;
               qM22_c19 <= qM22_c18;
               qP21_c19 <= qP21_c18;
               qM21_c19 <= qM21_c18;
               qP20_c19 <= qP20_c18;
               qM20_c19 <= qM20_c18;
               qP19_c19 <= qP19_c18;
               qM19_c19 <= qM19_c18;
               qP18_c19 <= qP18_c18;
               qM18_c19 <= qM18_c18;
               qP17_c19 <= qP17_c18;
               qM17_c19 <= qM17_c18;
               qP16_c19 <= qP16_c18;
               qM16_c19 <= qM16_c18;
               qP15_c19 <= qP15_c18;
               qM15_c19 <= qM15_c18;
               qP14_c19 <= qP14_c18;
               qM14_c19 <= qM14_c18;
               qP13_c19 <= qP13_c18;
               qM13_c19 <= qM13_c18;
            end if;
            if ce_20 = '1' then
               expR0_c20 <= expR0_c19;
               sR_c20 <= sR_c19;
               exnR0_c20 <= exnR0_c19;
               D_c20 <= D_c19;
               betaw12_c20 <= betaw12_c19;
               q12_copy21_c20 <= q12_copy21_c19;
               qP28_c20 <= qP28_c19;
               qM28_c20 <= qM28_c19;
               qP27_c20 <= qP27_c19;
               qM27_c20 <= qM27_c19;
               qP26_c20 <= qP26_c19;
               qM26_c20 <= qM26_c19;
               qP25_c20 <= qP25_c19;
               qM25_c20 <= qM25_c19;
               qP24_c20 <= qP24_c19;
               qM24_c20 <= qM24_c19;
               qP23_c20 <= qP23_c19;
               qM23_c20 <= qM23_c19;
               qP22_c20 <= qP22_c19;
               qM22_c20 <= qM22_c19;
               qP21_c20 <= qP21_c19;
               qM21_c20 <= qM21_c19;
               qP20_c20 <= qP20_c19;
               qM20_c20 <= qM20_c19;
               qP19_c20 <= qP19_c19;
               qM19_c20 <= qM19_c19;
               qP18_c20 <= qP18_c19;
               qM18_c20 <= qM18_c19;
               qP17_c20 <= qP17_c19;
               qM17_c20 <= qM17_c19;
               qP16_c20 <= qP16_c19;
               qM16_c20 <= qM16_c19;
               qP15_c20 <= qP15_c19;
               qM15_c20 <= qM15_c19;
               qP14_c20 <= qP14_c19;
               qM14_c20 <= qM14_c19;
               qP13_c20 <= qP13_c19;
               qM13_c20 <= qM13_c19;
            end if;
            if ce_21 = '1' then
               expR0_c21 <= expR0_c20;
               sR_c21 <= sR_c20;
               exnR0_c21 <= exnR0_c20;
               D_c21 <= D_c20;
               betaw12_c21 <= betaw12_c20;
               q12_c21 <= q12_c20;
               absq12D_c21 <= absq12D_c20;
               qP28_c21 <= qP28_c20;
               qM28_c21 <= qM28_c20;
               qP27_c21 <= qP27_c20;
               qM27_c21 <= qM27_c20;
               qP26_c21 <= qP26_c20;
               qM26_c21 <= qM26_c20;
               qP25_c21 <= qP25_c20;
               qM25_c21 <= qM25_c20;
               qP24_c21 <= qP24_c20;
               qM24_c21 <= qM24_c20;
               qP23_c21 <= qP23_c20;
               qM23_c21 <= qM23_c20;
               qP22_c21 <= qP22_c20;
               qM22_c21 <= qM22_c20;
               qP21_c21 <= qP21_c20;
               qM21_c21 <= qM21_c20;
               qP20_c21 <= qP20_c20;
               qM20_c21 <= qM20_c20;
               qP19_c21 <= qP19_c20;
               qM19_c21 <= qM19_c20;
               qP18_c21 <= qP18_c20;
               qM18_c21 <= qM18_c20;
               qP17_c21 <= qP17_c20;
               qM17_c21 <= qM17_c20;
               qP16_c21 <= qP16_c20;
               qM16_c21 <= qM16_c20;
               qP15_c21 <= qP15_c20;
               qM15_c21 <= qM15_c20;
               qP14_c21 <= qP14_c20;
               qM14_c21 <= qM14_c20;
               qP13_c21 <= qP13_c20;
               qM13_c21 <= qM13_c20;
               qP12_c21 <= qP12_c20;
               qM12_c21 <= qM12_c20;
            end if;
            if ce_22 = '1' then
               expR0_c22 <= expR0_c21;
               sR_c22 <= sR_c21;
               exnR0_c22 <= exnR0_c21;
               D_c22 <= D_c21;
               betaw11_c22 <= betaw11_c21;
               q11_c22 <= q11_c21;
               absq11D_c22 <= absq11D_c21;
               qP28_c22 <= qP28_c21;
               qM28_c22 <= qM28_c21;
               qP27_c22 <= qP27_c21;
               qM27_c22 <= qM27_c21;
               qP26_c22 <= qP26_c21;
               qM26_c22 <= qM26_c21;
               qP25_c22 <= qP25_c21;
               qM25_c22 <= qM25_c21;
               qP24_c22 <= qP24_c21;
               qM24_c22 <= qM24_c21;
               qP23_c22 <= qP23_c21;
               qM23_c22 <= qM23_c21;
               qP22_c22 <= qP22_c21;
               qM22_c22 <= qM22_c21;
               qP21_c22 <= qP21_c21;
               qM21_c22 <= qM21_c21;
               qP20_c22 <= qP20_c21;
               qM20_c22 <= qM20_c21;
               qP19_c22 <= qP19_c21;
               qM19_c22 <= qM19_c21;
               qP18_c22 <= qP18_c21;
               qM18_c22 <= qM18_c21;
               qP17_c22 <= qP17_c21;
               qM17_c22 <= qM17_c21;
               qP16_c22 <= qP16_c21;
               qM16_c22 <= qM16_c21;
               qP15_c22 <= qP15_c21;
               qM15_c22 <= qM15_c21;
               qP14_c22 <= qP14_c21;
               qM14_c22 <= qM14_c21;
               qP13_c22 <= qP13_c21;
               qM13_c22 <= qM13_c21;
               qP12_c22 <= qP12_c21;
               qM12_c22 <= qM12_c21;
               qP11_c22 <= qP11_c21;
               qM11_c22 <= qM11_c21;
            end if;
            if ce_23 = '1' then
               expR0_c23 <= expR0_c22;
               sR_c23 <= sR_c22;
               exnR0_c23 <= exnR0_c22;
               D_c23 <= D_c22;
               betaw10_c23 <= betaw10_c22;
               q10_c23 <= q10_c22;
               absq10D_c23 <= absq10D_c22;
               qP28_c23 <= qP28_c22;
               qM28_c23 <= qM28_c22;
               qP27_c23 <= qP27_c22;
               qM27_c23 <= qM27_c22;
               qP26_c23 <= qP26_c22;
               qM26_c23 <= qM26_c22;
               qP25_c23 <= qP25_c22;
               qM25_c23 <= qM25_c22;
               qP24_c23 <= qP24_c22;
               qM24_c23 <= qM24_c22;
               qP23_c23 <= qP23_c22;
               qM23_c23 <= qM23_c22;
               qP22_c23 <= qP22_c22;
               qM22_c23 <= qM22_c22;
               qP21_c23 <= qP21_c22;
               qM21_c23 <= qM21_c22;
               qP20_c23 <= qP20_c22;
               qM20_c23 <= qM20_c22;
               qP19_c23 <= qP19_c22;
               qM19_c23 <= qM19_c22;
               qP18_c23 <= qP18_c22;
               qM18_c23 <= qM18_c22;
               qP17_c23 <= qP17_c22;
               qM17_c23 <= qM17_c22;
               qP16_c23 <= qP16_c22;
               qM16_c23 <= qM16_c22;
               qP15_c23 <= qP15_c22;
               qM15_c23 <= qM15_c22;
               qP14_c23 <= qP14_c22;
               qM14_c23 <= qM14_c22;
               qP13_c23 <= qP13_c22;
               qM13_c23 <= qM13_c22;
               qP12_c23 <= qP12_c22;
               qM12_c23 <= qM12_c22;
               qP11_c23 <= qP11_c22;
               qM11_c23 <= qM11_c22;
               qP10_c23 <= qP10_c22;
               qM10_c23 <= qM10_c22;
            end if;
            if ce_24 = '1' then
               expR0_c24 <= expR0_c23;
               sR_c24 <= sR_c23;
               exnR0_c24 <= exnR0_c23;
               D_c24 <= D_c23;
               betaw9_c24 <= betaw9_c23;
               q9_c24 <= q9_c23;
               absq9D_c24 <= absq9D_c23;
               qP28_c24 <= qP28_c23;
               qM28_c24 <= qM28_c23;
               qP27_c24 <= qP27_c23;
               qM27_c24 <= qM27_c23;
               qP26_c24 <= qP26_c23;
               qM26_c24 <= qM26_c23;
               qP25_c24 <= qP25_c23;
               qM25_c24 <= qM25_c23;
               qP24_c24 <= qP24_c23;
               qM24_c24 <= qM24_c23;
               qP23_c24 <= qP23_c23;
               qM23_c24 <= qM23_c23;
               qP22_c24 <= qP22_c23;
               qM22_c24 <= qM22_c23;
               qP21_c24 <= qP21_c23;
               qM21_c24 <= qM21_c23;
               qP20_c24 <= qP20_c23;
               qM20_c24 <= qM20_c23;
               qP19_c24 <= qP19_c23;
               qM19_c24 <= qM19_c23;
               qP18_c24 <= qP18_c23;
               qM18_c24 <= qM18_c23;
               qP17_c24 <= qP17_c23;
               qM17_c24 <= qM17_c23;
               qP16_c24 <= qP16_c23;
               qM16_c24 <= qM16_c23;
               qP15_c24 <= qP15_c23;
               qM15_c24 <= qM15_c23;
               qP14_c24 <= qP14_c23;
               qM14_c24 <= qM14_c23;
               qP13_c24 <= qP13_c23;
               qM13_c24 <= qM13_c23;
               qP12_c24 <= qP12_c23;
               qM12_c24 <= qM12_c23;
               qP11_c24 <= qP11_c23;
               qM11_c24 <= qM11_c23;
               qP10_c24 <= qP10_c23;
               qM10_c24 <= qM10_c23;
               qP9_c24 <= qP9_c23;
               qM9_c24 <= qM9_c23;
            end if;
            if ce_25 = '1' then
               expR0_c25 <= expR0_c24;
               sR_c25 <= sR_c24;
               exnR0_c25 <= exnR0_c24;
               D_c25 <= D_c24;
               betaw8_c25 <= betaw8_c24;
               q8_copy25_c25 <= q8_copy25_c24;
               qP28_c25 <= qP28_c24;
               qM28_c25 <= qM28_c24;
               qP27_c25 <= qP27_c24;
               qM27_c25 <= qM27_c24;
               qP26_c25 <= qP26_c24;
               qM26_c25 <= qM26_c24;
               qP25_c25 <= qP25_c24;
               qM25_c25 <= qM25_c24;
               qP24_c25 <= qP24_c24;
               qM24_c25 <= qM24_c24;
               qP23_c25 <= qP23_c24;
               qM23_c25 <= qM23_c24;
               qP22_c25 <= qP22_c24;
               qM22_c25 <= qM22_c24;
               qP21_c25 <= qP21_c24;
               qM21_c25 <= qM21_c24;
               qP20_c25 <= qP20_c24;
               qM20_c25 <= qM20_c24;
               qP19_c25 <= qP19_c24;
               qM19_c25 <= qM19_c24;
               qP18_c25 <= qP18_c24;
               qM18_c25 <= qM18_c24;
               qP17_c25 <= qP17_c24;
               qM17_c25 <= qM17_c24;
               qP16_c25 <= qP16_c24;
               qM16_c25 <= qM16_c24;
               qP15_c25 <= qP15_c24;
               qM15_c25 <= qM15_c24;
               qP14_c25 <= qP14_c24;
               qM14_c25 <= qM14_c24;
               qP13_c25 <= qP13_c24;
               qM13_c25 <= qM13_c24;
               qP12_c25 <= qP12_c24;
               qM12_c25 <= qM12_c24;
               qP11_c25 <= qP11_c24;
               qM11_c25 <= qM11_c24;
               qP10_c25 <= qP10_c24;
               qM10_c25 <= qM10_c24;
               qP9_c25 <= qP9_c24;
               qM9_c25 <= qM9_c24;
            end if;
            if ce_26 = '1' then
               expR0_c26 <= expR0_c25;
               sR_c26 <= sR_c25;
               exnR0_c26 <= exnR0_c25;
               D_c26 <= D_c25;
               betaw8_c26 <= betaw8_c25;
               q8_c26 <= q8_c25;
               absq8D_c26 <= absq8D_c25;
               qP28_c26 <= qP28_c25;
               qM28_c26 <= qM28_c25;
               qP27_c26 <= qP27_c25;
               qM27_c26 <= qM27_c25;
               qP26_c26 <= qP26_c25;
               qM26_c26 <= qM26_c25;
               qP25_c26 <= qP25_c25;
               qM25_c26 <= qM25_c25;
               qP24_c26 <= qP24_c25;
               qM24_c26 <= qM24_c25;
               qP23_c26 <= qP23_c25;
               qM23_c26 <= qM23_c25;
               qP22_c26 <= qP22_c25;
               qM22_c26 <= qM22_c25;
               qP21_c26 <= qP21_c25;
               qM21_c26 <= qM21_c25;
               qP20_c26 <= qP20_c25;
               qM20_c26 <= qM20_c25;
               qP19_c26 <= qP19_c25;
               qM19_c26 <= qM19_c25;
               qP18_c26 <= qP18_c25;
               qM18_c26 <= qM18_c25;
               qP17_c26 <= qP17_c25;
               qM17_c26 <= qM17_c25;
               qP16_c26 <= qP16_c25;
               qM16_c26 <= qM16_c25;
               qP15_c26 <= qP15_c25;
               qM15_c26 <= qM15_c25;
               qP14_c26 <= qP14_c25;
               qM14_c26 <= qM14_c25;
               qP13_c26 <= qP13_c25;
               qM13_c26 <= qM13_c25;
               qP12_c26 <= qP12_c25;
               qM12_c26 <= qM12_c25;
               qP11_c26 <= qP11_c25;
               qM11_c26 <= qM11_c25;
               qP10_c26 <= qP10_c25;
               qM10_c26 <= qM10_c25;
               qP9_c26 <= qP9_c25;
               qM9_c26 <= qM9_c25;
               qP8_c26 <= qP8_c25;
               qM8_c26 <= qM8_c25;
            end if;
            if ce_27 = '1' then
               expR0_c27 <= expR0_c26;
               sR_c27 <= sR_c26;
               exnR0_c27 <= exnR0_c26;
               D_c27 <= D_c26;
               betaw7_c27 <= betaw7_c26;
               q7_c27 <= q7_c26;
               absq7D_c27 <= absq7D_c26;
               qP28_c27 <= qP28_c26;
               qM28_c27 <= qM28_c26;
               qP27_c27 <= qP27_c26;
               qM27_c27 <= qM27_c26;
               qP26_c27 <= qP26_c26;
               qM26_c27 <= qM26_c26;
               qP25_c27 <= qP25_c26;
               qM25_c27 <= qM25_c26;
               qP24_c27 <= qP24_c26;
               qM24_c27 <= qM24_c26;
               qP23_c27 <= qP23_c26;
               qM23_c27 <= qM23_c26;
               qP22_c27 <= qP22_c26;
               qM22_c27 <= qM22_c26;
               qP21_c27 <= qP21_c26;
               qM21_c27 <= qM21_c26;
               qP20_c27 <= qP20_c26;
               qM20_c27 <= qM20_c26;
               qP19_c27 <= qP19_c26;
               qM19_c27 <= qM19_c26;
               qP18_c27 <= qP18_c26;
               qM18_c27 <= qM18_c26;
               qP17_c27 <= qP17_c26;
               qM17_c27 <= qM17_c26;
               qP16_c27 <= qP16_c26;
               qM16_c27 <= qM16_c26;
               qP15_c27 <= qP15_c26;
               qM15_c27 <= qM15_c26;
               qP14_c27 <= qP14_c26;
               qM14_c27 <= qM14_c26;
               qP13_c27 <= qP13_c26;
               qM13_c27 <= qM13_c26;
               qP12_c27 <= qP12_c26;
               qM12_c27 <= qM12_c26;
               qP11_c27 <= qP11_c26;
               qM11_c27 <= qM11_c26;
               qP10_c27 <= qP10_c26;
               qM10_c27 <= qM10_c26;
               qP9_c27 <= qP9_c26;
               qM9_c27 <= qM9_c26;
               qP8_c27 <= qP8_c26;
               qM8_c27 <= qM8_c26;
               qP7_c27 <= qP7_c26;
               qM7_c27 <= qM7_c26;
            end if;
            if ce_28 = '1' then
               expR0_c28 <= expR0_c27;
               sR_c28 <= sR_c27;
               exnR0_c28 <= exnR0_c27;
               D_c28 <= D_c27;
               betaw6_c28 <= betaw6_c27;
               q6_c28 <= q6_c27;
               absq6D_c28 <= absq6D_c27;
               qP28_c28 <= qP28_c27;
               qM28_c28 <= qM28_c27;
               qP27_c28 <= qP27_c27;
               qM27_c28 <= qM27_c27;
               qP26_c28 <= qP26_c27;
               qM26_c28 <= qM26_c27;
               qP25_c28 <= qP25_c27;
               qM25_c28 <= qM25_c27;
               qP24_c28 <= qP24_c27;
               qM24_c28 <= qM24_c27;
               qP23_c28 <= qP23_c27;
               qM23_c28 <= qM23_c27;
               qP22_c28 <= qP22_c27;
               qM22_c28 <= qM22_c27;
               qP21_c28 <= qP21_c27;
               qM21_c28 <= qM21_c27;
               qP20_c28 <= qP20_c27;
               qM20_c28 <= qM20_c27;
               qP19_c28 <= qP19_c27;
               qM19_c28 <= qM19_c27;
               qP18_c28 <= qP18_c27;
               qM18_c28 <= qM18_c27;
               qP17_c28 <= qP17_c27;
               qM17_c28 <= qM17_c27;
               qP16_c28 <= qP16_c27;
               qM16_c28 <= qM16_c27;
               qP15_c28 <= qP15_c27;
               qM15_c28 <= qM15_c27;
               qP14_c28 <= qP14_c27;
               qM14_c28 <= qM14_c27;
               qP13_c28 <= qP13_c27;
               qM13_c28 <= qM13_c27;
               qP12_c28 <= qP12_c27;
               qM12_c28 <= qM12_c27;
               qP11_c28 <= qP11_c27;
               qM11_c28 <= qM11_c27;
               qP10_c28 <= qP10_c27;
               qM10_c28 <= qM10_c27;
               qP9_c28 <= qP9_c27;
               qM9_c28 <= qM9_c27;
               qP8_c28 <= qP8_c27;
               qM8_c28 <= qM8_c27;
               qP7_c28 <= qP7_c27;
               qM7_c28 <= qM7_c27;
               qP6_c28 <= qP6_c27;
               qM6_c28 <= qM6_c27;
            end if;
            if ce_29 = '1' then
               expR0_c29 <= expR0_c28;
               sR_c29 <= sR_c28;
               exnR0_c29 <= exnR0_c28;
               D_c29 <= D_c28;
               betaw5_c29 <= betaw5_c28;
               q5_c29 <= q5_c28;
               absq5D_c29 <= absq5D_c28;
               qP28_c29 <= qP28_c28;
               qM28_c29 <= qM28_c28;
               qP27_c29 <= qP27_c28;
               qM27_c29 <= qM27_c28;
               qP26_c29 <= qP26_c28;
               qM26_c29 <= qM26_c28;
               qP25_c29 <= qP25_c28;
               qM25_c29 <= qM25_c28;
               qP24_c29 <= qP24_c28;
               qM24_c29 <= qM24_c28;
               qP23_c29 <= qP23_c28;
               qM23_c29 <= qM23_c28;
               qP22_c29 <= qP22_c28;
               qM22_c29 <= qM22_c28;
               qP21_c29 <= qP21_c28;
               qM21_c29 <= qM21_c28;
               qP20_c29 <= qP20_c28;
               qM20_c29 <= qM20_c28;
               qP19_c29 <= qP19_c28;
               qM19_c29 <= qM19_c28;
               qP18_c29 <= qP18_c28;
               qM18_c29 <= qM18_c28;
               qP17_c29 <= qP17_c28;
               qM17_c29 <= qM17_c28;
               qP16_c29 <= qP16_c28;
               qM16_c29 <= qM16_c28;
               qP15_c29 <= qP15_c28;
               qM15_c29 <= qM15_c28;
               qP14_c29 <= qP14_c28;
               qM14_c29 <= qM14_c28;
               qP13_c29 <= qP13_c28;
               qM13_c29 <= qM13_c28;
               qP12_c29 <= qP12_c28;
               qM12_c29 <= qM12_c28;
               qP11_c29 <= qP11_c28;
               qM11_c29 <= qM11_c28;
               qP10_c29 <= qP10_c28;
               qM10_c29 <= qM10_c28;
               qP9_c29 <= qP9_c28;
               qM9_c29 <= qM9_c28;
               qP8_c29 <= qP8_c28;
               qM8_c29 <= qM8_c28;
               qP7_c29 <= qP7_c28;
               qM7_c29 <= qM7_c28;
               qP6_c29 <= qP6_c28;
               qM6_c29 <= qM6_c28;
               qP5_c29 <= qP5_c28;
               qM5_c29 <= qM5_c28;
            end if;
            if ce_30 = '1' then
               expR0_c30 <= expR0_c29;
               sR_c30 <= sR_c29;
               exnR0_c30 <= exnR0_c29;
               D_c30 <= D_c29;
               betaw4_c30 <= betaw4_c29;
               q4_copy29_c30 <= q4_copy29_c29;
               qP28_c30 <= qP28_c29;
               qM28_c30 <= qM28_c29;
               qP27_c30 <= qP27_c29;
               qM27_c30 <= qM27_c29;
               qP26_c30 <= qP26_c29;
               qM26_c30 <= qM26_c29;
               qP25_c30 <= qP25_c29;
               qM25_c30 <= qM25_c29;
               qP24_c30 <= qP24_c29;
               qM24_c30 <= qM24_c29;
               qP23_c30 <= qP23_c29;
               qM23_c30 <= qM23_c29;
               qP22_c30 <= qP22_c29;
               qM22_c30 <= qM22_c29;
               qP21_c30 <= qP21_c29;
               qM21_c30 <= qM21_c29;
               qP20_c30 <= qP20_c29;
               qM20_c30 <= qM20_c29;
               qP19_c30 <= qP19_c29;
               qM19_c30 <= qM19_c29;
               qP18_c30 <= qP18_c29;
               qM18_c30 <= qM18_c29;
               qP17_c30 <= qP17_c29;
               qM17_c30 <= qM17_c29;
               qP16_c30 <= qP16_c29;
               qM16_c30 <= qM16_c29;
               qP15_c30 <= qP15_c29;
               qM15_c30 <= qM15_c29;
               qP14_c30 <= qP14_c29;
               qM14_c30 <= qM14_c29;
               qP13_c30 <= qP13_c29;
               qM13_c30 <= qM13_c29;
               qP12_c30 <= qP12_c29;
               qM12_c30 <= qM12_c29;
               qP11_c30 <= qP11_c29;
               qM11_c30 <= qM11_c29;
               qP10_c30 <= qP10_c29;
               qM10_c30 <= qM10_c29;
               qP9_c30 <= qP9_c29;
               qM9_c30 <= qM9_c29;
               qP8_c30 <= qP8_c29;
               qM8_c30 <= qM8_c29;
               qP7_c30 <= qP7_c29;
               qM7_c30 <= qM7_c29;
               qP6_c30 <= qP6_c29;
               qM6_c30 <= qM6_c29;
               qP5_c30 <= qP5_c29;
               qM5_c30 <= qM5_c29;
            end if;
            if ce_31 = '1' then
               expR0_c31 <= expR0_c30;
               sR_c31 <= sR_c30;
               exnR0_c31 <= exnR0_c30;
               D_c31 <= D_c30;
               betaw4_c31 <= betaw4_c30;
               q4_c31 <= q4_c30;
               absq4D_c31 <= absq4D_c30;
               qP28_c31 <= qP28_c30;
               qM28_c31 <= qM28_c30;
               qP27_c31 <= qP27_c30;
               qM27_c31 <= qM27_c30;
               qP26_c31 <= qP26_c30;
               qM26_c31 <= qM26_c30;
               qP25_c31 <= qP25_c30;
               qM25_c31 <= qM25_c30;
               qP24_c31 <= qP24_c30;
               qM24_c31 <= qM24_c30;
               qP23_c31 <= qP23_c30;
               qM23_c31 <= qM23_c30;
               qP22_c31 <= qP22_c30;
               qM22_c31 <= qM22_c30;
               qP21_c31 <= qP21_c30;
               qM21_c31 <= qM21_c30;
               qP20_c31 <= qP20_c30;
               qM20_c31 <= qM20_c30;
               qP19_c31 <= qP19_c30;
               qM19_c31 <= qM19_c30;
               qP18_c31 <= qP18_c30;
               qM18_c31 <= qM18_c30;
               qP17_c31 <= qP17_c30;
               qM17_c31 <= qM17_c30;
               qP16_c31 <= qP16_c30;
               qM16_c31 <= qM16_c30;
               qP15_c31 <= qP15_c30;
               qM15_c31 <= qM15_c30;
               qP14_c31 <= qP14_c30;
               qM14_c31 <= qM14_c30;
               qP13_c31 <= qP13_c30;
               qM13_c31 <= qM13_c30;
               qP12_c31 <= qP12_c30;
               qM12_c31 <= qM12_c30;
               qP11_c31 <= qP11_c30;
               qM11_c31 <= qM11_c30;
               qP10_c31 <= qP10_c30;
               qM10_c31 <= qM10_c30;
               qP9_c31 <= qP9_c30;
               qM9_c31 <= qM9_c30;
               qP8_c31 <= qP8_c30;
               qM8_c31 <= qM8_c30;
               qP7_c31 <= qP7_c30;
               qM7_c31 <= qM7_c30;
               qP6_c31 <= qP6_c30;
               qM6_c31 <= qM6_c30;
               qP5_c31 <= qP5_c30;
               qM5_c31 <= qM5_c30;
               qP4_c31 <= qP4_c30;
               qM4_c31 <= qM4_c30;
            end if;
            if ce_32 = '1' then
               expR0_c32 <= expR0_c31;
               sR_c32 <= sR_c31;
               exnR0_c32 <= exnR0_c31;
               D_c32 <= D_c31;
               betaw3_c32 <= betaw3_c31;
               q3_c32 <= q3_c31;
               absq3D_c32 <= absq3D_c31;
               qP28_c32 <= qP28_c31;
               qM28_c32 <= qM28_c31;
               qP27_c32 <= qP27_c31;
               qM27_c32 <= qM27_c31;
               qP26_c32 <= qP26_c31;
               qM26_c32 <= qM26_c31;
               qP25_c32 <= qP25_c31;
               qM25_c32 <= qM25_c31;
               qP24_c32 <= qP24_c31;
               qM24_c32 <= qM24_c31;
               qP23_c32 <= qP23_c31;
               qM23_c32 <= qM23_c31;
               qP22_c32 <= qP22_c31;
               qM22_c32 <= qM22_c31;
               qP21_c32 <= qP21_c31;
               qM21_c32 <= qM21_c31;
               qP20_c32 <= qP20_c31;
               qM20_c32 <= qM20_c31;
               qP19_c32 <= qP19_c31;
               qM19_c32 <= qM19_c31;
               qP18_c32 <= qP18_c31;
               qM18_c32 <= qM18_c31;
               qP17_c32 <= qP17_c31;
               qM17_c32 <= qM17_c31;
               qP16_c32 <= qP16_c31;
               qM16_c32 <= qM16_c31;
               qP15_c32 <= qP15_c31;
               qM15_c32 <= qM15_c31;
               qP14_c32 <= qP14_c31;
               qM14_c32 <= qM14_c31;
               qP13_c32 <= qP13_c31;
               qM13_c32 <= qM13_c31;
               qP12_c32 <= qP12_c31;
               qM12_c32 <= qM12_c31;
               qP11_c32 <= qP11_c31;
               qM11_c32 <= qM11_c31;
               qP10_c32 <= qP10_c31;
               qM10_c32 <= qM10_c31;
               qP9_c32 <= qP9_c31;
               qM9_c32 <= qM9_c31;
               qP8_c32 <= qP8_c31;
               qM8_c32 <= qM8_c31;
               qP7_c32 <= qP7_c31;
               qM7_c32 <= qM7_c31;
               qP6_c32 <= qP6_c31;
               qM6_c32 <= qM6_c31;
               qP5_c32 <= qP5_c31;
               qM5_c32 <= qM5_c31;
               qP4_c32 <= qP4_c31;
               qM4_c32 <= qM4_c31;
               qP3_c32 <= qP3_c31;
               qM3_c32 <= qM3_c31;
            end if;
            if ce_33 = '1' then
               expR0_c33 <= expR0_c32;
               sR_c33 <= sR_c32;
               exnR0_c33 <= exnR0_c32;
               D_c33 <= D_c32;
               betaw2_c33 <= betaw2_c32;
               q2_c33 <= q2_c32;
               absq2D_c33 <= absq2D_c32;
               qP28_c33 <= qP28_c32;
               qM28_c33 <= qM28_c32;
               qP27_c33 <= qP27_c32;
               qM27_c33 <= qM27_c32;
               qP26_c33 <= qP26_c32;
               qM26_c33 <= qM26_c32;
               qP25_c33 <= qP25_c32;
               qM25_c33 <= qM25_c32;
               qP24_c33 <= qP24_c32;
               qM24_c33 <= qM24_c32;
               qP23_c33 <= qP23_c32;
               qM23_c33 <= qM23_c32;
               qP22_c33 <= qP22_c32;
               qM22_c33 <= qM22_c32;
               qP21_c33 <= qP21_c32;
               qM21_c33 <= qM21_c32;
               qP20_c33 <= qP20_c32;
               qM20_c33 <= qM20_c32;
               qP19_c33 <= qP19_c32;
               qM19_c33 <= qM19_c32;
               qP18_c33 <= qP18_c32;
               qM18_c33 <= qM18_c32;
               qP17_c33 <= qP17_c32;
               qM17_c33 <= qM17_c32;
               qP16_c33 <= qP16_c32;
               qM16_c33 <= qM16_c32;
               qP15_c33 <= qP15_c32;
               qM15_c33 <= qM15_c32;
               qP14_c33 <= qP14_c32;
               qM14_c33 <= qM14_c32;
               qP13_c33 <= qP13_c32;
               qM13_c33 <= qM13_c32;
               qP12_c33 <= qP12_c32;
               qM12_c33 <= qM12_c32;
               qP11_c33 <= qP11_c32;
               qM11_c33 <= qM11_c32;
               qP10_c33 <= qP10_c32;
               qM10_c33 <= qM10_c32;
               qP9_c33 <= qP9_c32;
               qM9_c33 <= qM9_c32;
               qP8_c33 <= qP8_c32;
               qM8_c33 <= qM8_c32;
               qP7_c33 <= qP7_c32;
               qM7_c33 <= qM7_c32;
               qP6_c33 <= qP6_c32;
               qM6_c33 <= qM6_c32;
               qP5_c33 <= qP5_c32;
               qM5_c33 <= qM5_c32;
               qP4_c33 <= qP4_c32;
               qM4_c33 <= qM4_c32;
               qP3_c33 <= qP3_c32;
               qM3_c33 <= qM3_c32;
               qP2_c33 <= qP2_c32;
               qM2_c33 <= qM2_c32;
            end if;
            if ce_34 = '1' then
               expR0_c34 <= expR0_c33;
               sR_c34 <= sR_c33;
               exnR0_c34 <= exnR0_c33;
               betaw1_c34 <= betaw1_c33;
               q1_c34 <= q1_c33;
               absq1D_c34 <= absq1D_c33;
               qM28_c34 <= qM28_c33;
               qM27_c34 <= qM27_c33;
               qM26_c34 <= qM26_c33;
               qM25_c34 <= qM25_c33;
               qM24_c34 <= qM24_c33;
               qM23_c34 <= qM23_c33;
               qM22_c34 <= qM22_c33;
               qM21_c34 <= qM21_c33;
               qM20_c34 <= qM20_c33;
               qM19_c34 <= qM19_c33;
               qM18_c34 <= qM18_c33;
               qM17_c34 <= qM17_c33;
               qM16_c34 <= qM16_c33;
               qM15_c34 <= qM15_c33;
               qM14_c34 <= qM14_c33;
               qM13_c34 <= qM13_c33;
               qM12_c34 <= qM12_c33;
               qM11_c34 <= qM11_c33;
               qM10_c34 <= qM10_c33;
               qM9_c34 <= qM9_c33;
               qM8_c34 <= qM8_c33;
               qM7_c34 <= qM7_c33;
               qM6_c34 <= qM6_c33;
               qM5_c34 <= qM5_c33;
               qM4_c34 <= qM4_c33;
               qM3_c34 <= qM3_c33;
               qM2_c34 <= qM2_c33;
               qM1_c34 <= qM1_c33;
               qP_c34 <= qP_c33;
            end if;
            if ce_35 = '1' then
               expR0_c35 <= expR0_c34;
               sR_c35 <= sR_c34;
               exnR0_c35 <= exnR0_c34;
               qP_c35 <= qP_c34;
               qM_c35 <= qM_c34;
            end if;
            if ce_36 = '1' then
               expR0_c36 <= expR0_c35;
               sR_c36 <= sR_c35;
               exnR0_c36 <= exnR0_c35;
               mR_c36 <= mR_c35;
               fRnorm_c36 <= fRnorm_c35;
               round_c36 <= round_c35;
            end if;
         end if;
      end process;
   fX_c0 <= "1" & X(51 downto 0);
   fY_c0 <= "1" & Y(51 downto 0);
   -- exponent difference, sign and exception combination computed early, to have fewer bits to pipeline
   expR0_c0 <= ("00" & X(62 downto 52)) - ("00" & Y(62 downto 52));
   sR_c0 <= X(63) xor Y(63);
   -- early exception handling 
   exnXY_c0 <= X(65 downto 64) & Y(65 downto 64);
   with exnXY_c0  select 
      exnR0_c0 <= 
         "01"	 when "0101",										-- normal
         "00"	 when "0001" | "0010" | "0110", -- zero
         "10"	 when "0100" | "1000" | "1001", -- overflow
         "11"	 when others;										-- NaN
   D_c0 <= fY_c0 ;
   psX_c0 <= "0" & fX_c0 ;
   betaw28_c0 <=  "00" & psX_c0;
   sel28_c0 <= betaw28_c0(55 downto 50) & D_c0(51 downto 49);
   SelFunctionTable28: selFunction_Freq500_uid4
      port map ( X => sel28_c0,
                 Y => q28_copy5_c0);
   q28_c0 <= q28_copy5_c0; -- output copy to hold a pipeline register if needed

   with q28_c0  select 
      absq28D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q28_c1(2)  select 
   w27_c1<= betaw28_c1 - absq28D_c1 when '0',
         betaw28_c1 + absq28D_c1 when others;

   betaw27_c1 <= w27_c1(53 downto 0) & "00"; -- multiplication by the radix
   sel27_c1 <= betaw27_c1(55 downto 50) & D_c1(51 downto 49);
   SelFunctionTable27: selFunction_Freq500_uid4
      port map ( X => sel27_c1,
                 Y => q27_copy6_c1);
   q27_c1 <= q27_copy6_c1; -- output copy to hold a pipeline register if needed

   with q27_c1  select 
      absq27D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q27_c2(2)  select 
   w26_c2<= betaw27_c2 - absq27D_c2 when '0',
         betaw27_c2 + absq27D_c2 when others;

   betaw26_c2 <= w26_c2(53 downto 0) & "00"; -- multiplication by the radix
   sel26_c2 <= betaw26_c2(55 downto 50) & D_c2(51 downto 49);
   SelFunctionTable26: selFunction_Freq500_uid4
      port map ( X => sel26_c2,
                 Y => q26_copy7_c2);
   q26_c2 <= q26_copy7_c2; -- output copy to hold a pipeline register if needed

   with q26_c2  select 
      absq26D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q26_c3(2)  select 
   w25_c3<= betaw26_c3 - absq26D_c3 when '0',
         betaw26_c3 + absq26D_c3 when others;

   betaw25_c3 <= w25_c3(53 downto 0) & "00"; -- multiplication by the radix
   sel25_c3 <= betaw25_c3(55 downto 50) & D_c3(51 downto 49);
   SelFunctionTable25: selFunction_Freq500_uid4
      port map ( X => sel25_c3,
                 Y => q25_copy8_c3);
   q25_c4 <= q25_copy8_c4; -- output copy to hold a pipeline register if needed

   with q25_c4  select 
      absq25D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q25_c4(2)  select 
   w24_c4<= betaw25_c4 - absq25D_c4 when '0',
         betaw25_c4 + absq25D_c4 when others;

   betaw24_c4 <= w24_c4(53 downto 0) & "00"; -- multiplication by the radix
   sel24_c4 <= betaw24_c4(55 downto 50) & D_c4(51 downto 49);
   SelFunctionTable24: selFunction_Freq500_uid4
      port map ( X => sel24_c4,
                 Y => q24_copy9_c4);
   q24_c5 <= q24_copy9_c5; -- output copy to hold a pipeline register if needed

   with q24_c5  select 
      absq24D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q24_c6(2)  select 
   w23_c6<= betaw24_c6 - absq24D_c6 when '0',
         betaw24_c6 + absq24D_c6 when others;

   betaw23_c6 <= w23_c6(53 downto 0) & "00"; -- multiplication by the radix
   sel23_c6 <= betaw23_c6(55 downto 50) & D_c6(51 downto 49);
   SelFunctionTable23: selFunction_Freq500_uid4
      port map ( X => sel23_c6,
                 Y => q23_copy10_c6);
   q23_c6 <= q23_copy10_c6; -- output copy to hold a pipeline register if needed

   with q23_c6  select 
      absq23D_c6 <= 
         "000" & D_c6						 when "001" | "111", -- mult by 1
         "00" & D_c6 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q23_c7(2)  select 
   w22_c7<= betaw23_c7 - absq23D_c7 when '0',
         betaw23_c7 + absq23D_c7 when others;

   betaw22_c7 <= w22_c7(53 downto 0) & "00"; -- multiplication by the radix
   sel22_c7 <= betaw22_c7(55 downto 50) & D_c7(51 downto 49);
   SelFunctionTable22: selFunction_Freq500_uid4
      port map ( X => sel22_c7,
                 Y => q22_copy11_c7);
   q22_c7 <= q22_copy11_c7; -- output copy to hold a pipeline register if needed

   with q22_c7  select 
      absq22D_c7 <= 
         "000" & D_c7						 when "001" | "111", -- mult by 1
         "00" & D_c7 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q22_c8(2)  select 
   w21_c8<= betaw22_c8 - absq22D_c8 when '0',
         betaw22_c8 + absq22D_c8 when others;

   betaw21_c8 <= w21_c8(53 downto 0) & "00"; -- multiplication by the radix
   sel21_c8 <= betaw21_c8(55 downto 50) & D_c8(51 downto 49);
   SelFunctionTable21: selFunction_Freq500_uid4
      port map ( X => sel21_c8,
                 Y => q21_copy12_c8);
   q21_c9 <= q21_copy12_c9; -- output copy to hold a pipeline register if needed

   with q21_c9  select 
      absq21D_c9 <= 
         "000" & D_c9						 when "001" | "111", -- mult by 1
         "00" & D_c9 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q21_c9(2)  select 
   w20_c9<= betaw21_c9 - absq21D_c9 when '0',
         betaw21_c9 + absq21D_c9 when others;

   betaw20_c9 <= w20_c9(53 downto 0) & "00"; -- multiplication by the radix
   sel20_c9 <= betaw20_c9(55 downto 50) & D_c9(51 downto 49);
   SelFunctionTable20: selFunction_Freq500_uid4
      port map ( X => sel20_c9,
                 Y => q20_copy13_c9);
   q20_c10 <= q20_copy13_c10; -- output copy to hold a pipeline register if needed

   with q20_c10  select 
      absq20D_c10 <= 
         "000" & D_c10						 when "001" | "111", -- mult by 1
         "00" & D_c10 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q20_c11(2)  select 
   w19_c11<= betaw20_c11 - absq20D_c11 when '0',
         betaw20_c11 + absq20D_c11 when others;

   betaw19_c11 <= w19_c11(53 downto 0) & "00"; -- multiplication by the radix
   sel19_c11 <= betaw19_c11(55 downto 50) & D_c11(51 downto 49);
   SelFunctionTable19: selFunction_Freq500_uid4
      port map ( X => sel19_c11,
                 Y => q19_copy14_c11);
   q19_c11 <= q19_copy14_c11; -- output copy to hold a pipeline register if needed

   with q19_c11  select 
      absq19D_c11 <= 
         "000" & D_c11						 when "001" | "111", -- mult by 1
         "00" & D_c11 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q19_c12(2)  select 
   w18_c12<= betaw19_c12 - absq19D_c12 when '0',
         betaw19_c12 + absq19D_c12 when others;

   betaw18_c12 <= w18_c12(53 downto 0) & "00"; -- multiplication by the radix
   sel18_c12 <= betaw18_c12(55 downto 50) & D_c12(51 downto 49);
   SelFunctionTable18: selFunction_Freq500_uid4
      port map ( X => sel18_c12,
                 Y => q18_copy15_c12);
   q18_c12 <= q18_copy15_c12; -- output copy to hold a pipeline register if needed

   with q18_c12  select 
      absq18D_c12 <= 
         "000" & D_c12						 when "001" | "111", -- mult by 1
         "00" & D_c12 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q18_c13(2)  select 
   w17_c13<= betaw18_c13 - absq18D_c13 when '0',
         betaw18_c13 + absq18D_c13 when others;

   betaw17_c13 <= w17_c13(53 downto 0) & "00"; -- multiplication by the radix
   sel17_c13 <= betaw17_c13(55 downto 50) & D_c13(51 downto 49);
   SelFunctionTable17: selFunction_Freq500_uid4
      port map ( X => sel17_c13,
                 Y => q17_copy16_c13);
   q17_c14 <= q17_copy16_c14; -- output copy to hold a pipeline register if needed

   with q17_c14  select 
      absq17D_c14 <= 
         "000" & D_c14						 when "001" | "111", -- mult by 1
         "00" & D_c14 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q17_c14(2)  select 
   w16_c14<= betaw17_c14 - absq17D_c14 when '0',
         betaw17_c14 + absq17D_c14 when others;

   betaw16_c14 <= w16_c14(53 downto 0) & "00"; -- multiplication by the radix
   sel16_c14 <= betaw16_c14(55 downto 50) & D_c14(51 downto 49);
   SelFunctionTable16: selFunction_Freq500_uid4
      port map ( X => sel16_c14,
                 Y => q16_copy17_c14);
   q16_c15 <= q16_copy17_c15; -- output copy to hold a pipeline register if needed

   with q16_c15  select 
      absq16D_c15 <= 
         "000" & D_c15						 when "001" | "111", -- mult by 1
         "00" & D_c15 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q16_c16(2)  select 
   w15_c16<= betaw16_c16 - absq16D_c16 when '0',
         betaw16_c16 + absq16D_c16 when others;

   betaw15_c16 <= w15_c16(53 downto 0) & "00"; -- multiplication by the radix
   sel15_c16 <= betaw15_c16(55 downto 50) & D_c16(51 downto 49);
   SelFunctionTable15: selFunction_Freq500_uid4
      port map ( X => sel15_c16,
                 Y => q15_copy18_c16);
   q15_c16 <= q15_copy18_c16; -- output copy to hold a pipeline register if needed

   with q15_c16  select 
      absq15D_c16 <= 
         "000" & D_c16						 when "001" | "111", -- mult by 1
         "00" & D_c16 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q15_c17(2)  select 
   w14_c17<= betaw15_c17 - absq15D_c17 when '0',
         betaw15_c17 + absq15D_c17 when others;

   betaw14_c17 <= w14_c17(53 downto 0) & "00"; -- multiplication by the radix
   sel14_c17 <= betaw14_c17(55 downto 50) & D_c17(51 downto 49);
   SelFunctionTable14: selFunction_Freq500_uid4
      port map ( X => sel14_c17,
                 Y => q14_copy19_c17);
   q14_c17 <= q14_copy19_c17; -- output copy to hold a pipeline register if needed

   with q14_c17  select 
      absq14D_c17 <= 
         "000" & D_c17						 when "001" | "111", -- mult by 1
         "00" & D_c17 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q14_c18(2)  select 
   w13_c18<= betaw14_c18 - absq14D_c18 when '0',
         betaw14_c18 + absq14D_c18 when others;

   betaw13_c18 <= w13_c18(53 downto 0) & "00"; -- multiplication by the radix
   sel13_c18 <= betaw13_c18(55 downto 50) & D_c18(51 downto 49);
   SelFunctionTable13: selFunction_Freq500_uid4
      port map ( X => sel13_c18,
                 Y => q13_copy20_c18);
   q13_c18 <= q13_copy20_c18; -- output copy to hold a pipeline register if needed

   with q13_c18  select 
      absq13D_c18 <= 
         "000" & D_c18						 when "001" | "111", -- mult by 1
         "00" & D_c18 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q13_c19(2)  select 
   w12_c19<= betaw13_c19 - absq13D_c19 when '0',
         betaw13_c19 + absq13D_c19 when others;

   betaw12_c19 <= w12_c19(53 downto 0) & "00"; -- multiplication by the radix
   sel12_c19 <= betaw12_c19(55 downto 50) & D_c19(51 downto 49);
   SelFunctionTable12: selFunction_Freq500_uid4
      port map ( X => sel12_c19,
                 Y => q12_copy21_c19);
   q12_c20 <= q12_copy21_c20; -- output copy to hold a pipeline register if needed

   with q12_c20  select 
      absq12D_c20 <= 
         "000" & D_c20						 when "001" | "111", -- mult by 1
         "00" & D_c20 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q12_c21(2)  select 
   w11_c21<= betaw12_c21 - absq12D_c21 when '0',
         betaw12_c21 + absq12D_c21 when others;

   betaw11_c21 <= w11_c21(53 downto 0) & "00"; -- multiplication by the radix
   sel11_c21 <= betaw11_c21(55 downto 50) & D_c21(51 downto 49);
   SelFunctionTable11: selFunction_Freq500_uid4
      port map ( X => sel11_c21,
                 Y => q11_copy22_c21);
   q11_c21 <= q11_copy22_c21; -- output copy to hold a pipeline register if needed

   with q11_c21  select 
      absq11D_c21 <= 
         "000" & D_c21						 when "001" | "111", -- mult by 1
         "00" & D_c21 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q11_c22(2)  select 
   w10_c22<= betaw11_c22 - absq11D_c22 when '0',
         betaw11_c22 + absq11D_c22 when others;

   betaw10_c22 <= w10_c22(53 downto 0) & "00"; -- multiplication by the radix
   sel10_c22 <= betaw10_c22(55 downto 50) & D_c22(51 downto 49);
   SelFunctionTable10: selFunction_Freq500_uid4
      port map ( X => sel10_c22,
                 Y => q10_copy23_c22);
   q10_c22 <= q10_copy23_c22; -- output copy to hold a pipeline register if needed

   with q10_c22  select 
      absq10D_c22 <= 
         "000" & D_c22						 when "001" | "111", -- mult by 1
         "00" & D_c22 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q10_c23(2)  select 
   w9_c23<= betaw10_c23 - absq10D_c23 when '0',
         betaw10_c23 + absq10D_c23 when others;

   betaw9_c23 <= w9_c23(53 downto 0) & "00"; -- multiplication by the radix
   sel9_c23 <= betaw9_c23(55 downto 50) & D_c23(51 downto 49);
   SelFunctionTable9: selFunction_Freq500_uid4
      port map ( X => sel9_c23,
                 Y => q9_copy24_c23);
   q9_c23 <= q9_copy24_c23; -- output copy to hold a pipeline register if needed

   with q9_c23  select 
      absq9D_c23 <= 
         "000" & D_c23						 when "001" | "111", -- mult by 1
         "00" & D_c23 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q9_c24(2)  select 
   w8_c24<= betaw9_c24 - absq9D_c24 when '0',
         betaw9_c24 + absq9D_c24 when others;

   betaw8_c24 <= w8_c24(53 downto 0) & "00"; -- multiplication by the radix
   sel8_c24 <= betaw8_c24(55 downto 50) & D_c24(51 downto 49);
   SelFunctionTable8: selFunction_Freq500_uid4
      port map ( X => sel8_c24,
                 Y => q8_copy25_c24);
   q8_c25 <= q8_copy25_c25; -- output copy to hold a pipeline register if needed

   with q8_c25  select 
      absq8D_c25 <= 
         "000" & D_c25						 when "001" | "111", -- mult by 1
         "00" & D_c25 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q8_c26(2)  select 
   w7_c26<= betaw8_c26 - absq8D_c26 when '0',
         betaw8_c26 + absq8D_c26 when others;

   betaw7_c26 <= w7_c26(53 downto 0) & "00"; -- multiplication by the radix
   sel7_c26 <= betaw7_c26(55 downto 50) & D_c26(51 downto 49);
   SelFunctionTable7: selFunction_Freq500_uid4
      port map ( X => sel7_c26,
                 Y => q7_copy26_c26);
   q7_c26 <= q7_copy26_c26; -- output copy to hold a pipeline register if needed

   with q7_c26  select 
      absq7D_c26 <= 
         "000" & D_c26						 when "001" | "111", -- mult by 1
         "00" & D_c26 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q7_c27(2)  select 
   w6_c27<= betaw7_c27 - absq7D_c27 when '0',
         betaw7_c27 + absq7D_c27 when others;

   betaw6_c27 <= w6_c27(53 downto 0) & "00"; -- multiplication by the radix
   sel6_c27 <= betaw6_c27(55 downto 50) & D_c27(51 downto 49);
   SelFunctionTable6: selFunction_Freq500_uid4
      port map ( X => sel6_c27,
                 Y => q6_copy27_c27);
   q6_c27 <= q6_copy27_c27; -- output copy to hold a pipeline register if needed

   with q6_c27  select 
      absq6D_c27 <= 
         "000" & D_c27						 when "001" | "111", -- mult by 1
         "00" & D_c27 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q6_c28(2)  select 
   w5_c28<= betaw6_c28 - absq6D_c28 when '0',
         betaw6_c28 + absq6D_c28 when others;

   betaw5_c28 <= w5_c28(53 downto 0) & "00"; -- multiplication by the radix
   sel5_c28 <= betaw5_c28(55 downto 50) & D_c28(51 downto 49);
   SelFunctionTable5: selFunction_Freq500_uid4
      port map ( X => sel5_c28,
                 Y => q5_copy28_c28);
   q5_c28 <= q5_copy28_c28; -- output copy to hold a pipeline register if needed

   with q5_c28  select 
      absq5D_c28 <= 
         "000" & D_c28						 when "001" | "111", -- mult by 1
         "00" & D_c28 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q5_c29(2)  select 
   w4_c29<= betaw5_c29 - absq5D_c29 when '0',
         betaw5_c29 + absq5D_c29 when others;

   betaw4_c29 <= w4_c29(53 downto 0) & "00"; -- multiplication by the radix
   sel4_c29 <= betaw4_c29(55 downto 50) & D_c29(51 downto 49);
   SelFunctionTable4: selFunction_Freq500_uid4
      port map ( X => sel4_c29,
                 Y => q4_copy29_c29);
   q4_c30 <= q4_copy29_c30; -- output copy to hold a pipeline register if needed

   with q4_c30  select 
      absq4D_c30 <= 
         "000" & D_c30						 when "001" | "111", -- mult by 1
         "00" & D_c30 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q4_c31(2)  select 
   w3_c31<= betaw4_c31 - absq4D_c31 when '0',
         betaw4_c31 + absq4D_c31 when others;

   betaw3_c31 <= w3_c31(53 downto 0) & "00"; -- multiplication by the radix
   sel3_c31 <= betaw3_c31(55 downto 50) & D_c31(51 downto 49);
   SelFunctionTable3: selFunction_Freq500_uid4
      port map ( X => sel3_c31,
                 Y => q3_copy30_c31);
   q3_c31 <= q3_copy30_c31; -- output copy to hold a pipeline register if needed

   with q3_c31  select 
      absq3D_c31 <= 
         "000" & D_c31						 when "001" | "111", -- mult by 1
         "00" & D_c31 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q3_c32(2)  select 
   w2_c32<= betaw3_c32 - absq3D_c32 when '0',
         betaw3_c32 + absq3D_c32 when others;

   betaw2_c32 <= w2_c32(53 downto 0) & "00"; -- multiplication by the radix
   sel2_c32 <= betaw2_c32(55 downto 50) & D_c32(51 downto 49);
   SelFunctionTable2: selFunction_Freq500_uid4
      port map ( X => sel2_c32,
                 Y => q2_copy31_c32);
   q2_c32 <= q2_copy31_c32; -- output copy to hold a pipeline register if needed

   with q2_c32  select 
      absq2D_c32 <= 
         "000" & D_c32						 when "001" | "111", -- mult by 1
         "00" & D_c32 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q2_c33(2)  select 
   w1_c33<= betaw2_c33 - absq2D_c33 when '0',
         betaw2_c33 + absq2D_c33 when others;

   betaw1_c33 <= w1_c33(53 downto 0) & "00"; -- multiplication by the radix
   sel1_c33 <= betaw1_c33(55 downto 50) & D_c33(51 downto 49);
   SelFunctionTable1: selFunction_Freq500_uid4
      port map ( X => sel1_c33,
                 Y => q1_copy32_c33);
   q1_c33 <= q1_copy32_c33; -- output copy to hold a pipeline register if needed

   with q1_c33  select 
      absq1D_c33 <= 
         "000" & D_c33						 when "001" | "111", -- mult by 1
         "00" & D_c33 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q1_c34(2)  select 
   w0_c34<= betaw1_c34 - absq1D_c34 when '0',
         betaw1_c34 + absq1D_c34 when others;

   wfinal_c34 <= w0_c34(53 downto 0);
   qM0_c34 <= wfinal_c34(53); -- rounding bit is the sign of the remainder
   qP28_c0 <=      q28_c0(1 downto 0);
   qM28_c0 <=      q28_c0(2) & "0";
   qP27_c1 <=      q27_c1(1 downto 0);
   qM27_c1 <=      q27_c1(2) & "0";
   qP26_c2 <=      q26_c2(1 downto 0);
   qM26_c2 <=      q26_c2(2) & "0";
   qP25_c4 <=      q25_c4(1 downto 0);
   qM25_c4 <=      q25_c4(2) & "0";
   qP24_c5 <=      q24_c5(1 downto 0);
   qM24_c5 <=      q24_c5(2) & "0";
   qP23_c6 <=      q23_c6(1 downto 0);
   qM23_c6 <=      q23_c6(2) & "0";
   qP22_c7 <=      q22_c7(1 downto 0);
   qM22_c7 <=      q22_c7(2) & "0";
   qP21_c9 <=      q21_c9(1 downto 0);
   qM21_c9 <=      q21_c9(2) & "0";
   qP20_c10 <=      q20_c10(1 downto 0);
   qM20_c10 <=      q20_c10(2) & "0";
   qP19_c11 <=      q19_c11(1 downto 0);
   qM19_c11 <=      q19_c11(2) & "0";
   qP18_c12 <=      q18_c12(1 downto 0);
   qM18_c12 <=      q18_c12(2) & "0";
   qP17_c14 <=      q17_c14(1 downto 0);
   qM17_c14 <=      q17_c14(2) & "0";
   qP16_c15 <=      q16_c15(1 downto 0);
   qM16_c15 <=      q16_c15(2) & "0";
   qP15_c16 <=      q15_c16(1 downto 0);
   qM15_c16 <=      q15_c16(2) & "0";
   qP14_c17 <=      q14_c17(1 downto 0);
   qM14_c17 <=      q14_c17(2) & "0";
   qP13_c18 <=      q13_c18(1 downto 0);
   qM13_c18 <=      q13_c18(2) & "0";
   qP12_c20 <=      q12_c20(1 downto 0);
   qM12_c20 <=      q12_c20(2) & "0";
   qP11_c21 <=      q11_c21(1 downto 0);
   qM11_c21 <=      q11_c21(2) & "0";
   qP10_c22 <=      q10_c22(1 downto 0);
   qM10_c22 <=      q10_c22(2) & "0";
   qP9_c23 <=      q9_c23(1 downto 0);
   qM9_c23 <=      q9_c23(2) & "0";
   qP8_c25 <=      q8_c25(1 downto 0);
   qM8_c25 <=      q8_c25(2) & "0";
   qP7_c26 <=      q7_c26(1 downto 0);
   qM7_c26 <=      q7_c26(2) & "0";
   qP6_c27 <=      q6_c27(1 downto 0);
   qM6_c27 <=      q6_c27(2) & "0";
   qP5_c28 <=      q5_c28(1 downto 0);
   qM5_c28 <=      q5_c28(2) & "0";
   qP4_c30 <=      q4_c30(1 downto 0);
   qM4_c30 <=      q4_c30(2) & "0";
   qP3_c31 <=      q3_c31(1 downto 0);
   qM3_c31 <=      q3_c31(2) & "0";
   qP2_c32 <=      q2_c32(1 downto 0);
   qM2_c32 <=      q2_c32(2) & "0";
   qP1_c33 <=      q1_c33(1 downto 0);
   qM1_c33 <=      q1_c33(2) & "0";
   qP_c33 <= qP28_c33 & qP27_c33 & qP26_c33 & qP25_c33 & qP24_c33 & qP23_c33 & qP22_c33 & qP21_c33 & qP20_c33 & qP19_c33 & qP18_c33 & qP17_c33 & qP16_c33 & qP15_c33 & qP14_c33 & qP13_c33 & qP12_c33 & qP11_c33 & qP10_c33 & qP9_c33 & qP8_c33 & qP7_c33 & qP6_c33 & qP5_c33 & qP4_c33 & qP3_c33 & qP2_c33 & qP1_c33;
   qM_c34 <= qM28_c34(0) & qM27_c34 & qM26_c34 & qM25_c34 & qM24_c34 & qM23_c34 & qM22_c34 & qM21_c34 & qM20_c34 & qM19_c34 & qM18_c34 & qM17_c34 & qM16_c34 & qM15_c34 & qM14_c34 & qM13_c34 & qM12_c34 & qM11_c34 & qM10_c34 & qM9_c34 & qM8_c34 & qM7_c34 & qM6_c34 & qM5_c34 & qM4_c34 & qM3_c34 & qM2_c34 & qM1_c34 & qM0_c34;
   quotient_c35 <= qP_c35 - qM_c35;
   -- We need a mR in (0, -wf-2) format: 1+wF fraction bits, 1 round bit, and 1 guard bit for the normalisation,
   -- quotient is the truncation of the exact quotient to at least 2^(-wF-2) bits
   -- now discarding its possible known MSB zeroes, and dropping the possible extra LSB bit (due to radix 4) 
   mR_c35 <= quotient_c35(54 downto 0); 
   -- normalisation
   fRnorm_c35 <=    mR_c35(53 downto 1)  when mR_c35(54)= '1'
           else mR_c35(52 downto 0);  -- now fRnorm is a (-1, -wF-1) fraction
   round_c35 <= fRnorm_c35(0); 
   expR1_c36 <= expR0_c36 + ("000" & (9 downto 1 => '1') & mR_c36(54)); -- add back bias
   -- final rounding
   expfrac_c36 <= expR1_c36 & fRnorm_c36(52 downto 1) ;
   expfracR_c36 <= expfrac_c36 + ((64 downto 1 => '0') & round_c36);
   exnR_c36 <=      "00"  when expfracR_c36(64) = '1'   -- underflow
           else "10"  when  expfracR_c36(64 downto 63) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_c36  select 
      exnRfinal_c36 <= 
         exnR_c36   when "01", -- normal
         exnR0_c36  when others;
   R <= exnRfinal_c36 & sR_c36 & expfracR_c36(62 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          selFunction_Freq300_uid4
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity selFunction_Freq300_uid4 is
    port (X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of selFunction_Freq300_uid4 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000000000",
      "000" when "000000001",
      "000" when "000000010",
      "000" when "000000011",
      "000" when "000000100",
      "000" when "000000101",
      "000" when "000000110",
      "000" when "000000111",
      "000" when "000001000",
      "000" when "000001001",
      "000" when "000001010",
      "000" when "000001011",
      "000" when "000001100",
      "000" when "000001101",
      "000" when "000001110",
      "000" when "000001111",
      "001" when "000010000",
      "000" when "000010001",
      "000" when "000010010",
      "000" when "000010011",
      "000" when "000010100",
      "000" when "000010101",
      "000" when "000010110",
      "000" when "000010111",
      "001" when "000011000",
      "001" when "000011001",
      "001" when "000011010",
      "001" when "000011011",
      "000" when "000011100",
      "000" when "000011101",
      "000" when "000011110",
      "000" when "000011111",
      "001" when "000100000",
      "001" when "000100001",
      "001" when "000100010",
      "001" when "000100011",
      "001" when "000100100",
      "001" when "000100101",
      "001" when "000100110",
      "000" when "000100111",
      "001" when "000101000",
      "001" when "000101001",
      "001" when "000101010",
      "001" when "000101011",
      "001" when "000101100",
      "001" when "000101101",
      "001" when "000101110",
      "001" when "000101111",
      "010" when "000110000",
      "001" when "000110001",
      "001" when "000110010",
      "001" when "000110011",
      "001" when "000110100",
      "001" when "000110101",
      "001" when "000110110",
      "001" when "000110111",
      "010" when "000111000",
      "010" when "000111001",
      "001" when "000111010",
      "001" when "000111011",
      "001" when "000111100",
      "001" when "000111101",
      "001" when "000111110",
      "001" when "000111111",
      "010" when "001000000",
      "010" when "001000001",
      "010" when "001000010",
      "001" when "001000011",
      "001" when "001000100",
      "001" when "001000101",
      "001" when "001000110",
      "001" when "001000111",
      "010" when "001001000",
      "010" when "001001001",
      "010" when "001001010",
      "010" when "001001011",
      "001" when "001001100",
      "001" when "001001101",
      "001" when "001001110",
      "001" when "001001111",
      "010" when "001010000",
      "010" when "001010001",
      "010" when "001010010",
      "010" when "001010011",
      "010" when "001010100",
      "010" when "001010101",
      "001" when "001010110",
      "001" when "001010111",
      "010" when "001011000",
      "010" when "001011001",
      "010" when "001011010",
      "010" when "001011011",
      "010" when "001011100",
      "010" when "001011101",
      "010" when "001011110",
      "001" when "001011111",
      "010" when "001100000",
      "010" when "001100001",
      "010" when "001100010",
      "010" when "001100011",
      "010" when "001100100",
      "010" when "001100101",
      "010" when "001100110",
      "010" when "001100111",
      "010" when "001101000",
      "010" when "001101001",
      "010" when "001101010",
      "010" when "001101011",
      "010" when "001101100",
      "010" when "001101101",
      "010" when "001101110",
      "010" when "001101111",
      "010" when "001110000",
      "010" when "001110001",
      "010" when "001110010",
      "010" when "001110011",
      "010" when "001110100",
      "010" when "001110101",
      "010" when "001110110",
      "010" when "001110111",
      "010" when "001111000",
      "010" when "001111001",
      "010" when "001111010",
      "010" when "001111011",
      "010" when "001111100",
      "010" when "001111101",
      "010" when "001111110",
      "010" when "001111111",
      "010" when "010000000",
      "010" when "010000001",
      "010" when "010000010",
      "010" when "010000011",
      "010" when "010000100",
      "010" when "010000101",
      "010" when "010000110",
      "010" when "010000111",
      "010" when "010001000",
      "010" when "010001001",
      "010" when "010001010",
      "010" when "010001011",
      "010" when "010001100",
      "010" when "010001101",
      "010" when "010001110",
      "010" when "010001111",
      "010" when "010010000",
      "010" when "010010001",
      "010" when "010010010",
      "010" when "010010011",
      "010" when "010010100",
      "010" when "010010101",
      "010" when "010010110",
      "010" when "010010111",
      "010" when "010011000",
      "010" when "010011001",
      "010" when "010011010",
      "010" when "010011011",
      "010" when "010011100",
      "010" when "010011101",
      "010" when "010011110",
      "010" when "010011111",
      "010" when "010100000",
      "010" when "010100001",
      "010" when "010100010",
      "010" when "010100011",
      "010" when "010100100",
      "010" when "010100101",
      "010" when "010100110",
      "010" when "010100111",
      "010" when "010101000",
      "010" when "010101001",
      "010" when "010101010",
      "010" when "010101011",
      "010" when "010101100",
      "010" when "010101101",
      "010" when "010101110",
      "010" when "010101111",
      "010" when "010110000",
      "010" when "010110001",
      "010" when "010110010",
      "010" when "010110011",
      "010" when "010110100",
      "010" when "010110101",
      "010" when "010110110",
      "010" when "010110111",
      "010" when "010111000",
      "010" when "010111001",
      "010" when "010111010",
      "010" when "010111011",
      "010" when "010111100",
      "010" when "010111101",
      "010" when "010111110",
      "010" when "010111111",
      "010" when "011000000",
      "010" when "011000001",
      "010" when "011000010",
      "010" when "011000011",
      "010" when "011000100",
      "010" when "011000101",
      "010" when "011000110",
      "010" when "011000111",
      "010" when "011001000",
      "010" when "011001001",
      "010" when "011001010",
      "010" when "011001011",
      "010" when "011001100",
      "010" when "011001101",
      "010" when "011001110",
      "010" when "011001111",
      "010" when "011010000",
      "010" when "011010001",
      "010" when "011010010",
      "010" when "011010011",
      "010" when "011010100",
      "010" when "011010101",
      "010" when "011010110",
      "010" when "011010111",
      "010" when "011011000",
      "010" when "011011001",
      "010" when "011011010",
      "010" when "011011011",
      "010" when "011011100",
      "010" when "011011101",
      "010" when "011011110",
      "010" when "011011111",
      "010" when "011100000",
      "010" when "011100001",
      "010" when "011100010",
      "010" when "011100011",
      "010" when "011100100",
      "010" when "011100101",
      "010" when "011100110",
      "010" when "011100111",
      "010" when "011101000",
      "010" when "011101001",
      "010" when "011101010",
      "010" when "011101011",
      "010" when "011101100",
      "010" when "011101101",
      "010" when "011101110",
      "010" when "011101111",
      "010" when "011110000",
      "010" when "011110001",
      "010" when "011110010",
      "010" when "011110011",
      "010" when "011110100",
      "010" when "011110101",
      "010" when "011110110",
      "010" when "011110111",
      "010" when "011111000",
      "010" when "011111001",
      "010" when "011111010",
      "010" when "011111011",
      "010" when "011111100",
      "010" when "011111101",
      "010" when "011111110",
      "010" when "011111111",
      "110" when "100000000",
      "110" when "100000001",
      "110" when "100000010",
      "110" when "100000011",
      "110" when "100000100",
      "110" when "100000101",
      "110" when "100000110",
      "110" when "100000111",
      "110" when "100001000",
      "110" when "100001001",
      "110" when "100001010",
      "110" when "100001011",
      "110" when "100001100",
      "110" when "100001101",
      "110" when "100001110",
      "110" when "100001111",
      "110" when "100010000",
      "110" when "100010001",
      "110" when "100010010",
      "110" when "100010011",
      "110" when "100010100",
      "110" when "100010101",
      "110" when "100010110",
      "110" when "100010111",
      "110" when "100011000",
      "110" when "100011001",
      "110" when "100011010",
      "110" when "100011011",
      "110" when "100011100",
      "110" when "100011101",
      "110" when "100011110",
      "110" when "100011111",
      "110" when "100100000",
      "110" when "100100001",
      "110" when "100100010",
      "110" when "100100011",
      "110" when "100100100",
      "110" when "100100101",
      "110" when "100100110",
      "110" when "100100111",
      "110" when "100101000",
      "110" when "100101001",
      "110" when "100101010",
      "110" when "100101011",
      "110" when "100101100",
      "110" when "100101101",
      "110" when "100101110",
      "110" when "100101111",
      "110" when "100110000",
      "110" when "100110001",
      "110" when "100110010",
      "110" when "100110011",
      "110" when "100110100",
      "110" when "100110101",
      "110" when "100110110",
      "110" when "100110111",
      "110" when "100111000",
      "110" when "100111001",
      "110" when "100111010",
      "110" when "100111011",
      "110" when "100111100",
      "110" when "100111101",
      "110" when "100111110",
      "110" when "100111111",
      "110" when "101000000",
      "110" when "101000001",
      "110" when "101000010",
      "110" when "101000011",
      "110" when "101000100",
      "110" when "101000101",
      "110" when "101000110",
      "110" when "101000111",
      "110" when "101001000",
      "110" when "101001001",
      "110" when "101001010",
      "110" when "101001011",
      "110" when "101001100",
      "110" when "101001101",
      "110" when "101001110",
      "110" when "101001111",
      "110" when "101010000",
      "110" when "101010001",
      "110" when "101010010",
      "110" when "101010011",
      "110" when "101010100",
      "110" when "101010101",
      "110" when "101010110",
      "110" when "101010111",
      "110" when "101011000",
      "110" when "101011001",
      "110" when "101011010",
      "110" when "101011011",
      "110" when "101011100",
      "110" when "101011101",
      "110" when "101011110",
      "110" when "101011111",
      "110" when "101100000",
      "110" when "101100001",
      "110" when "101100010",
      "110" when "101100011",
      "110" when "101100100",
      "110" when "101100101",
      "110" when "101100110",
      "110" when "101100111",
      "110" when "101101000",
      "110" when "101101001",
      "110" when "101101010",
      "110" when "101101011",
      "110" when "101101100",
      "110" when "101101101",
      "110" when "101101110",
      "110" when "101101111",
      "110" when "101110000",
      "110" when "101110001",
      "110" when "101110010",
      "110" when "101110011",
      "110" when "101110100",
      "110" when "101110101",
      "110" when "101110110",
      "110" when "101110111",
      "110" when "101111000",
      "110" when "101111001",
      "110" when "101111010",
      "110" when "101111011",
      "110" when "101111100",
      "110" when "101111101",
      "110" when "101111110",
      "110" when "101111111",
      "110" when "110000000",
      "110" when "110000001",
      "110" when "110000010",
      "110" when "110000011",
      "110" when "110000100",
      "110" when "110000101",
      "110" when "110000110",
      "110" when "110000111",
      "110" when "110001000",
      "110" when "110001001",
      "110" when "110001010",
      "110" when "110001011",
      "110" when "110001100",
      "110" when "110001101",
      "110" when "110001110",
      "110" when "110001111",
      "110" when "110010000",
      "110" when "110010001",
      "110" when "110010010",
      "110" when "110010011",
      "110" when "110010100",
      "110" when "110010101",
      "110" when "110010110",
      "110" when "110010111",
      "110" when "110011000",
      "110" when "110011001",
      "110" when "110011010",
      "110" when "110011011",
      "110" when "110011100",
      "110" when "110011101",
      "110" when "110011110",
      "110" when "110011111",
      "110" when "110100000",
      "110" when "110100001",
      "110" when "110100010",
      "110" when "110100011",
      "110" when "110100100",
      "110" when "110100101",
      "110" when "110100110",
      "110" when "110100111",
      "110" when "110101000",
      "110" when "110101001",
      "110" when "110101010",
      "110" when "110101011",
      "110" when "110101100",
      "110" when "110101101",
      "110" when "110101110",
      "111" when "110101111",
      "110" when "110110000",
      "110" when "110110001",
      "110" when "110110010",
      "110" when "110110011",
      "110" when "110110100",
      "111" when "110110101",
      "111" when "110110110",
      "111" when "110110111",
      "110" when "110111000",
      "110" when "110111001",
      "110" when "110111010",
      "110" when "110111011",
      "111" when "110111100",
      "111" when "110111101",
      "111" when "110111110",
      "111" when "110111111",
      "110" when "111000000",
      "110" when "111000001",
      "111" when "111000010",
      "111" when "111000011",
      "111" when "111000100",
      "111" when "111000101",
      "111" when "111000110",
      "111" when "111000111",
      "110" when "111001000",
      "111" when "111001001",
      "111" when "111001010",
      "111" when "111001011",
      "111" when "111001100",
      "111" when "111001101",
      "111" when "111001110",
      "111" when "111001111",
      "111" when "111010000",
      "111" when "111010001",
      "111" when "111010010",
      "111" when "111010011",
      "111" when "111010100",
      "111" when "111010101",
      "111" when "111010110",
      "111" when "111010111",
      "111" when "111011000",
      "111" when "111011001",
      "111" when "111011010",
      "111" when "111011011",
      "111" when "111011100",
      "111" when "111011101",
      "111" when "111011110",
      "111" when "111011111",
      "111" when "111100000",
      "111" when "111100001",
      "111" when "111100010",
      "111" when "111100011",
      "111" when "111100100",
      "111" when "111100101",
      "111" when "111100110",
      "111" when "111100111",
      "111" when "111101000",
      "111" when "111101001",
      "111" when "111101010",
      "111" when "111101011",
      "000" when "111101100",
      "000" when "111101101",
      "000" when "111101110",
      "000" when "111101111",
      "000" when "111110000",
      "000" when "111110001",
      "000" when "111110010",
      "000" when "111110011",
      "000" when "111110100",
      "000" when "111110101",
      "000" when "111110110",
      "000" when "111110111",
      "000" when "111111000",
      "000" when "111111001",
      "000" when "111111010",
      "000" when "111111011",
      "000" when "111111100",
      "000" when "111111101",
      "000" when "111111110",
      "000" when "111111111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            FloatingPointDivider
--                         (FPDiv_11_52_Freq300_uid2)
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 20 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointDivider_64_6_859333 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15, ce_16, ce_17, ce_18, ce_19, ce_20 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointDivider_64_6_859333 is
   component selFunction_Freq300_uid4 is
      port ( X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal fX_c0 :  std_logic_vector(52 downto 0);
signal fY_c0 :  std_logic_vector(52 downto 0);
signal expR0_c0, expR0_c1, expR0_c2, expR0_c3, expR0_c4, expR0_c5, expR0_c6, expR0_c7, expR0_c8, expR0_c9, expR0_c10, expR0_c11, expR0_c12, expR0_c13, expR0_c14, expR0_c15, expR0_c16, expR0_c17, expR0_c18, expR0_c19, expR0_c20 :  std_logic_vector(12 downto 0);
signal sR_c0, sR_c1, sR_c2, sR_c3, sR_c4, sR_c5, sR_c6, sR_c7, sR_c8, sR_c9, sR_c10, sR_c11, sR_c12, sR_c13, sR_c14, sR_c15, sR_c16, sR_c17, sR_c18, sR_c19, sR_c20 :  std_logic;
signal exnXY_c0 :  std_logic_vector(3 downto 0);
signal exnR0_c0, exnR0_c1, exnR0_c2, exnR0_c3, exnR0_c4, exnR0_c5, exnR0_c6, exnR0_c7, exnR0_c8, exnR0_c9, exnR0_c10, exnR0_c11, exnR0_c12, exnR0_c13, exnR0_c14, exnR0_c15, exnR0_c16, exnR0_c17, exnR0_c18, exnR0_c19, exnR0_c20 :  std_logic_vector(1 downto 0);
signal D_c0, D_c1, D_c2, D_c3, D_c4, D_c5, D_c6, D_c7, D_c8, D_c9, D_c10, D_c11, D_c12, D_c13, D_c14, D_c15, D_c16, D_c17, D_c18, D_c19 :  std_logic_vector(52 downto 0);
signal psX_c0 :  std_logic_vector(53 downto 0);
signal betaw28_c0 :  std_logic_vector(55 downto 0);
signal sel28_c0 :  std_logic_vector(8 downto 0);
signal q28_c0 :  std_logic_vector(2 downto 0);
signal q28_copy5_c0 :  std_logic_vector(2 downto 0);
signal absq28D_c0 :  std_logic_vector(55 downto 0);
signal w27_c0 :  std_logic_vector(55 downto 0);
signal betaw27_c0, betaw27_c1 :  std_logic_vector(55 downto 0);
signal sel27_c0 :  std_logic_vector(8 downto 0);
signal q27_c0, q27_c1 :  std_logic_vector(2 downto 0);
signal q27_copy6_c0 :  std_logic_vector(2 downto 0);
signal absq27D_c0, absq27D_c1 :  std_logic_vector(55 downto 0);
signal w26_c1 :  std_logic_vector(55 downto 0);
signal betaw26_c1, betaw26_c2 :  std_logic_vector(55 downto 0);
signal sel26_c1 :  std_logic_vector(8 downto 0);
signal q26_c1, q26_c2 :  std_logic_vector(2 downto 0);
signal q26_copy7_c1 :  std_logic_vector(2 downto 0);
signal absq26D_c1, absq26D_c2 :  std_logic_vector(55 downto 0);
signal w25_c2 :  std_logic_vector(55 downto 0);
signal betaw25_c2 :  std_logic_vector(55 downto 0);
signal sel25_c2 :  std_logic_vector(8 downto 0);
signal q25_c2 :  std_logic_vector(2 downto 0);
signal q25_copy8_c2 :  std_logic_vector(2 downto 0);
signal absq25D_c2 :  std_logic_vector(55 downto 0);
signal w24_c2 :  std_logic_vector(55 downto 0);
signal betaw24_c2, betaw24_c3 :  std_logic_vector(55 downto 0);
signal sel24_c2 :  std_logic_vector(8 downto 0);
signal q24_c3 :  std_logic_vector(2 downto 0);
signal q24_copy9_c2, q24_copy9_c3 :  std_logic_vector(2 downto 0);
signal absq24D_c3 :  std_logic_vector(55 downto 0);
signal w23_c3 :  std_logic_vector(55 downto 0);
signal betaw23_c3, betaw23_c4 :  std_logic_vector(55 downto 0);
signal sel23_c3 :  std_logic_vector(8 downto 0);
signal q23_c3, q23_c4 :  std_logic_vector(2 downto 0);
signal q23_copy10_c3 :  std_logic_vector(2 downto 0);
signal absq23D_c3, absq23D_c4 :  std_logic_vector(55 downto 0);
signal w22_c4 :  std_logic_vector(55 downto 0);
signal betaw22_c4 :  std_logic_vector(55 downto 0);
signal sel22_c4 :  std_logic_vector(8 downto 0);
signal q22_c4 :  std_logic_vector(2 downto 0);
signal q22_copy11_c4 :  std_logic_vector(2 downto 0);
signal absq22D_c4 :  std_logic_vector(55 downto 0);
signal w21_c4 :  std_logic_vector(55 downto 0);
signal betaw21_c4, betaw21_c5 :  std_logic_vector(55 downto 0);
signal sel21_c4 :  std_logic_vector(8 downto 0);
signal q21_c5 :  std_logic_vector(2 downto 0);
signal q21_copy12_c4, q21_copy12_c5 :  std_logic_vector(2 downto 0);
signal absq21D_c5 :  std_logic_vector(55 downto 0);
signal w20_c5 :  std_logic_vector(55 downto 0);
signal betaw20_c5, betaw20_c6 :  std_logic_vector(55 downto 0);
signal sel20_c5 :  std_logic_vector(8 downto 0);
signal q20_c5, q20_c6 :  std_logic_vector(2 downto 0);
signal q20_copy13_c5 :  std_logic_vector(2 downto 0);
signal absq20D_c5, absq20D_c6 :  std_logic_vector(55 downto 0);
signal w19_c6 :  std_logic_vector(55 downto 0);
signal betaw19_c6, betaw19_c7 :  std_logic_vector(55 downto 0);
signal sel19_c6 :  std_logic_vector(8 downto 0);
signal q19_c6, q19_c7 :  std_logic_vector(2 downto 0);
signal q19_copy14_c6 :  std_logic_vector(2 downto 0);
signal absq19D_c6, absq19D_c7 :  std_logic_vector(55 downto 0);
signal w18_c7 :  std_logic_vector(55 downto 0);
signal betaw18_c7 :  std_logic_vector(55 downto 0);
signal sel18_c7 :  std_logic_vector(8 downto 0);
signal q18_c7 :  std_logic_vector(2 downto 0);
signal q18_copy15_c7 :  std_logic_vector(2 downto 0);
signal absq18D_c7 :  std_logic_vector(55 downto 0);
signal w17_c7 :  std_logic_vector(55 downto 0);
signal betaw17_c7, betaw17_c8 :  std_logic_vector(55 downto 0);
signal sel17_c7 :  std_logic_vector(8 downto 0);
signal q17_c8 :  std_logic_vector(2 downto 0);
signal q17_copy16_c7, q17_copy16_c8 :  std_logic_vector(2 downto 0);
signal absq17D_c8 :  std_logic_vector(55 downto 0);
signal w16_c8 :  std_logic_vector(55 downto 0);
signal betaw16_c8, betaw16_c9 :  std_logic_vector(55 downto 0);
signal sel16_c8 :  std_logic_vector(8 downto 0);
signal q16_c8, q16_c9 :  std_logic_vector(2 downto 0);
signal q16_copy17_c8 :  std_logic_vector(2 downto 0);
signal absq16D_c8, absq16D_c9 :  std_logic_vector(55 downto 0);
signal w15_c9 :  std_logic_vector(55 downto 0);
signal betaw15_c9 :  std_logic_vector(55 downto 0);
signal sel15_c9 :  std_logic_vector(8 downto 0);
signal q15_c9 :  std_logic_vector(2 downto 0);
signal q15_copy18_c9 :  std_logic_vector(2 downto 0);
signal absq15D_c9 :  std_logic_vector(55 downto 0);
signal w14_c9 :  std_logic_vector(55 downto 0);
signal betaw14_c9, betaw14_c10 :  std_logic_vector(55 downto 0);
signal sel14_c9 :  std_logic_vector(8 downto 0);
signal q14_c10 :  std_logic_vector(2 downto 0);
signal q14_copy19_c9, q14_copy19_c10 :  std_logic_vector(2 downto 0);
signal absq14D_c10 :  std_logic_vector(55 downto 0);
signal w13_c10 :  std_logic_vector(55 downto 0);
signal betaw13_c10, betaw13_c11 :  std_logic_vector(55 downto 0);
signal sel13_c10 :  std_logic_vector(8 downto 0);
signal q13_c10, q13_c11 :  std_logic_vector(2 downto 0);
signal q13_copy20_c10 :  std_logic_vector(2 downto 0);
signal absq13D_c10, absq13D_c11 :  std_logic_vector(55 downto 0);
signal w12_c11 :  std_logic_vector(55 downto 0);
signal betaw12_c11, betaw12_c12 :  std_logic_vector(55 downto 0);
signal sel12_c11 :  std_logic_vector(8 downto 0);
signal q12_c11, q12_c12 :  std_logic_vector(2 downto 0);
signal q12_copy21_c11 :  std_logic_vector(2 downto 0);
signal absq12D_c11, absq12D_c12 :  std_logic_vector(55 downto 0);
signal w11_c12 :  std_logic_vector(55 downto 0);
signal betaw11_c12 :  std_logic_vector(55 downto 0);
signal sel11_c12 :  std_logic_vector(8 downto 0);
signal q11_c12 :  std_logic_vector(2 downto 0);
signal q11_copy22_c12 :  std_logic_vector(2 downto 0);
signal absq11D_c12 :  std_logic_vector(55 downto 0);
signal w10_c12 :  std_logic_vector(55 downto 0);
signal betaw10_c12, betaw10_c13 :  std_logic_vector(55 downto 0);
signal sel10_c12 :  std_logic_vector(8 downto 0);
signal q10_c13 :  std_logic_vector(2 downto 0);
signal q10_copy23_c12, q10_copy23_c13 :  std_logic_vector(2 downto 0);
signal absq10D_c13 :  std_logic_vector(55 downto 0);
signal w9_c13 :  std_logic_vector(55 downto 0);
signal betaw9_c13, betaw9_c14 :  std_logic_vector(55 downto 0);
signal sel9_c13 :  std_logic_vector(8 downto 0);
signal q9_c13, q9_c14 :  std_logic_vector(2 downto 0);
signal q9_copy24_c13 :  std_logic_vector(2 downto 0);
signal absq9D_c13, absq9D_c14 :  std_logic_vector(55 downto 0);
signal w8_c14 :  std_logic_vector(55 downto 0);
signal betaw8_c14 :  std_logic_vector(55 downto 0);
signal sel8_c14 :  std_logic_vector(8 downto 0);
signal q8_c14 :  std_logic_vector(2 downto 0);
signal q8_copy25_c14 :  std_logic_vector(2 downto 0);
signal absq8D_c14 :  std_logic_vector(55 downto 0);
signal w7_c14 :  std_logic_vector(55 downto 0);
signal betaw7_c14, betaw7_c15 :  std_logic_vector(55 downto 0);
signal sel7_c14 :  std_logic_vector(8 downto 0);
signal q7_c15 :  std_logic_vector(2 downto 0);
signal q7_copy26_c14, q7_copy26_c15 :  std_logic_vector(2 downto 0);
signal absq7D_c15 :  std_logic_vector(55 downto 0);
signal w6_c15 :  std_logic_vector(55 downto 0);
signal betaw6_c15, betaw6_c16 :  std_logic_vector(55 downto 0);
signal sel6_c15 :  std_logic_vector(8 downto 0);
signal q6_c15, q6_c16 :  std_logic_vector(2 downto 0);
signal q6_copy27_c15 :  std_logic_vector(2 downto 0);
signal absq6D_c15, absq6D_c16 :  std_logic_vector(55 downto 0);
signal w5_c16 :  std_logic_vector(55 downto 0);
signal betaw5_c16, betaw5_c17 :  std_logic_vector(55 downto 0);
signal sel5_c16 :  std_logic_vector(8 downto 0);
signal q5_c16, q5_c17 :  std_logic_vector(2 downto 0);
signal q5_copy28_c16 :  std_logic_vector(2 downto 0);
signal absq5D_c16, absq5D_c17 :  std_logic_vector(55 downto 0);
signal w4_c17 :  std_logic_vector(55 downto 0);
signal betaw4_c17 :  std_logic_vector(55 downto 0);
signal sel4_c17 :  std_logic_vector(8 downto 0);
signal q4_c17 :  std_logic_vector(2 downto 0);
signal q4_copy29_c17 :  std_logic_vector(2 downto 0);
signal absq4D_c17 :  std_logic_vector(55 downto 0);
signal w3_c17 :  std_logic_vector(55 downto 0);
signal betaw3_c17, betaw3_c18 :  std_logic_vector(55 downto 0);
signal sel3_c17 :  std_logic_vector(8 downto 0);
signal q3_c18 :  std_logic_vector(2 downto 0);
signal q3_copy30_c17, q3_copy30_c18 :  std_logic_vector(2 downto 0);
signal absq3D_c18 :  std_logic_vector(55 downto 0);
signal w2_c18 :  std_logic_vector(55 downto 0);
signal betaw2_c18, betaw2_c19 :  std_logic_vector(55 downto 0);
signal sel2_c18 :  std_logic_vector(8 downto 0);
signal q2_c18, q2_c19 :  std_logic_vector(2 downto 0);
signal q2_copy31_c18 :  std_logic_vector(2 downto 0);
signal absq2D_c18, absq2D_c19 :  std_logic_vector(55 downto 0);
signal w1_c19 :  std_logic_vector(55 downto 0);
signal betaw1_c19 :  std_logic_vector(55 downto 0);
signal sel1_c19 :  std_logic_vector(8 downto 0);
signal q1_c19 :  std_logic_vector(2 downto 0);
signal q1_copy32_c19 :  std_logic_vector(2 downto 0);
signal absq1D_c19 :  std_logic_vector(55 downto 0);
signal w0_c19 :  std_logic_vector(55 downto 0);
signal wfinal_c19 :  std_logic_vector(53 downto 0);
signal qM0_c19 :  std_logic;
signal qP28_c0, qP28_c1, qP28_c2, qP28_c3, qP28_c4, qP28_c5, qP28_c6, qP28_c7, qP28_c8, qP28_c9, qP28_c10, qP28_c11, qP28_c12, qP28_c13, qP28_c14, qP28_c15, qP28_c16, qP28_c17, qP28_c18, qP28_c19 :  std_logic_vector(1 downto 0);
signal qM28_c0, qM28_c1, qM28_c2, qM28_c3, qM28_c4, qM28_c5, qM28_c6, qM28_c7, qM28_c8, qM28_c9, qM28_c10, qM28_c11, qM28_c12, qM28_c13, qM28_c14, qM28_c15, qM28_c16, qM28_c17, qM28_c18, qM28_c19 :  std_logic_vector(1 downto 0);
signal qP27_c0, qP27_c1, qP27_c2, qP27_c3, qP27_c4, qP27_c5, qP27_c6, qP27_c7, qP27_c8, qP27_c9, qP27_c10, qP27_c11, qP27_c12, qP27_c13, qP27_c14, qP27_c15, qP27_c16, qP27_c17, qP27_c18, qP27_c19 :  std_logic_vector(1 downto 0);
signal qM27_c0, qM27_c1, qM27_c2, qM27_c3, qM27_c4, qM27_c5, qM27_c6, qM27_c7, qM27_c8, qM27_c9, qM27_c10, qM27_c11, qM27_c12, qM27_c13, qM27_c14, qM27_c15, qM27_c16, qM27_c17, qM27_c18, qM27_c19 :  std_logic_vector(1 downto 0);
signal qP26_c1, qP26_c2, qP26_c3, qP26_c4, qP26_c5, qP26_c6, qP26_c7, qP26_c8, qP26_c9, qP26_c10, qP26_c11, qP26_c12, qP26_c13, qP26_c14, qP26_c15, qP26_c16, qP26_c17, qP26_c18, qP26_c19 :  std_logic_vector(1 downto 0);
signal qM26_c1, qM26_c2, qM26_c3, qM26_c4, qM26_c5, qM26_c6, qM26_c7, qM26_c8, qM26_c9, qM26_c10, qM26_c11, qM26_c12, qM26_c13, qM26_c14, qM26_c15, qM26_c16, qM26_c17, qM26_c18, qM26_c19 :  std_logic_vector(1 downto 0);
signal qP25_c2, qP25_c3, qP25_c4, qP25_c5, qP25_c6, qP25_c7, qP25_c8, qP25_c9, qP25_c10, qP25_c11, qP25_c12, qP25_c13, qP25_c14, qP25_c15, qP25_c16, qP25_c17, qP25_c18, qP25_c19 :  std_logic_vector(1 downto 0);
signal qM25_c2, qM25_c3, qM25_c4, qM25_c5, qM25_c6, qM25_c7, qM25_c8, qM25_c9, qM25_c10, qM25_c11, qM25_c12, qM25_c13, qM25_c14, qM25_c15, qM25_c16, qM25_c17, qM25_c18, qM25_c19 :  std_logic_vector(1 downto 0);
signal qP24_c3, qP24_c4, qP24_c5, qP24_c6, qP24_c7, qP24_c8, qP24_c9, qP24_c10, qP24_c11, qP24_c12, qP24_c13, qP24_c14, qP24_c15, qP24_c16, qP24_c17, qP24_c18, qP24_c19 :  std_logic_vector(1 downto 0);
signal qM24_c3, qM24_c4, qM24_c5, qM24_c6, qM24_c7, qM24_c8, qM24_c9, qM24_c10, qM24_c11, qM24_c12, qM24_c13, qM24_c14, qM24_c15, qM24_c16, qM24_c17, qM24_c18, qM24_c19 :  std_logic_vector(1 downto 0);
signal qP23_c3, qP23_c4, qP23_c5, qP23_c6, qP23_c7, qP23_c8, qP23_c9, qP23_c10, qP23_c11, qP23_c12, qP23_c13, qP23_c14, qP23_c15, qP23_c16, qP23_c17, qP23_c18, qP23_c19 :  std_logic_vector(1 downto 0);
signal qM23_c3, qM23_c4, qM23_c5, qM23_c6, qM23_c7, qM23_c8, qM23_c9, qM23_c10, qM23_c11, qM23_c12, qM23_c13, qM23_c14, qM23_c15, qM23_c16, qM23_c17, qM23_c18, qM23_c19 :  std_logic_vector(1 downto 0);
signal qP22_c4, qP22_c5, qP22_c6, qP22_c7, qP22_c8, qP22_c9, qP22_c10, qP22_c11, qP22_c12, qP22_c13, qP22_c14, qP22_c15, qP22_c16, qP22_c17, qP22_c18, qP22_c19 :  std_logic_vector(1 downto 0);
signal qM22_c4, qM22_c5, qM22_c6, qM22_c7, qM22_c8, qM22_c9, qM22_c10, qM22_c11, qM22_c12, qM22_c13, qM22_c14, qM22_c15, qM22_c16, qM22_c17, qM22_c18, qM22_c19 :  std_logic_vector(1 downto 0);
signal qP21_c5, qP21_c6, qP21_c7, qP21_c8, qP21_c9, qP21_c10, qP21_c11, qP21_c12, qP21_c13, qP21_c14, qP21_c15, qP21_c16, qP21_c17, qP21_c18, qP21_c19 :  std_logic_vector(1 downto 0);
signal qM21_c5, qM21_c6, qM21_c7, qM21_c8, qM21_c9, qM21_c10, qM21_c11, qM21_c12, qM21_c13, qM21_c14, qM21_c15, qM21_c16, qM21_c17, qM21_c18, qM21_c19 :  std_logic_vector(1 downto 0);
signal qP20_c5, qP20_c6, qP20_c7, qP20_c8, qP20_c9, qP20_c10, qP20_c11, qP20_c12, qP20_c13, qP20_c14, qP20_c15, qP20_c16, qP20_c17, qP20_c18, qP20_c19 :  std_logic_vector(1 downto 0);
signal qM20_c5, qM20_c6, qM20_c7, qM20_c8, qM20_c9, qM20_c10, qM20_c11, qM20_c12, qM20_c13, qM20_c14, qM20_c15, qM20_c16, qM20_c17, qM20_c18, qM20_c19 :  std_logic_vector(1 downto 0);
signal qP19_c6, qP19_c7, qP19_c8, qP19_c9, qP19_c10, qP19_c11, qP19_c12, qP19_c13, qP19_c14, qP19_c15, qP19_c16, qP19_c17, qP19_c18, qP19_c19 :  std_logic_vector(1 downto 0);
signal qM19_c6, qM19_c7, qM19_c8, qM19_c9, qM19_c10, qM19_c11, qM19_c12, qM19_c13, qM19_c14, qM19_c15, qM19_c16, qM19_c17, qM19_c18, qM19_c19 :  std_logic_vector(1 downto 0);
signal qP18_c7, qP18_c8, qP18_c9, qP18_c10, qP18_c11, qP18_c12, qP18_c13, qP18_c14, qP18_c15, qP18_c16, qP18_c17, qP18_c18, qP18_c19 :  std_logic_vector(1 downto 0);
signal qM18_c7, qM18_c8, qM18_c9, qM18_c10, qM18_c11, qM18_c12, qM18_c13, qM18_c14, qM18_c15, qM18_c16, qM18_c17, qM18_c18, qM18_c19 :  std_logic_vector(1 downto 0);
signal qP17_c8, qP17_c9, qP17_c10, qP17_c11, qP17_c12, qP17_c13, qP17_c14, qP17_c15, qP17_c16, qP17_c17, qP17_c18, qP17_c19 :  std_logic_vector(1 downto 0);
signal qM17_c8, qM17_c9, qM17_c10, qM17_c11, qM17_c12, qM17_c13, qM17_c14, qM17_c15, qM17_c16, qM17_c17, qM17_c18, qM17_c19 :  std_logic_vector(1 downto 0);
signal qP16_c8, qP16_c9, qP16_c10, qP16_c11, qP16_c12, qP16_c13, qP16_c14, qP16_c15, qP16_c16, qP16_c17, qP16_c18, qP16_c19 :  std_logic_vector(1 downto 0);
signal qM16_c8, qM16_c9, qM16_c10, qM16_c11, qM16_c12, qM16_c13, qM16_c14, qM16_c15, qM16_c16, qM16_c17, qM16_c18, qM16_c19 :  std_logic_vector(1 downto 0);
signal qP15_c9, qP15_c10, qP15_c11, qP15_c12, qP15_c13, qP15_c14, qP15_c15, qP15_c16, qP15_c17, qP15_c18, qP15_c19 :  std_logic_vector(1 downto 0);
signal qM15_c9, qM15_c10, qM15_c11, qM15_c12, qM15_c13, qM15_c14, qM15_c15, qM15_c16, qM15_c17, qM15_c18, qM15_c19 :  std_logic_vector(1 downto 0);
signal qP14_c10, qP14_c11, qP14_c12, qP14_c13, qP14_c14, qP14_c15, qP14_c16, qP14_c17, qP14_c18, qP14_c19 :  std_logic_vector(1 downto 0);
signal qM14_c10, qM14_c11, qM14_c12, qM14_c13, qM14_c14, qM14_c15, qM14_c16, qM14_c17, qM14_c18, qM14_c19 :  std_logic_vector(1 downto 0);
signal qP13_c10, qP13_c11, qP13_c12, qP13_c13, qP13_c14, qP13_c15, qP13_c16, qP13_c17, qP13_c18, qP13_c19 :  std_logic_vector(1 downto 0);
signal qM13_c10, qM13_c11, qM13_c12, qM13_c13, qM13_c14, qM13_c15, qM13_c16, qM13_c17, qM13_c18, qM13_c19 :  std_logic_vector(1 downto 0);
signal qP12_c11, qP12_c12, qP12_c13, qP12_c14, qP12_c15, qP12_c16, qP12_c17, qP12_c18, qP12_c19 :  std_logic_vector(1 downto 0);
signal qM12_c11, qM12_c12, qM12_c13, qM12_c14, qM12_c15, qM12_c16, qM12_c17, qM12_c18, qM12_c19 :  std_logic_vector(1 downto 0);
signal qP11_c12, qP11_c13, qP11_c14, qP11_c15, qP11_c16, qP11_c17, qP11_c18, qP11_c19 :  std_logic_vector(1 downto 0);
signal qM11_c12, qM11_c13, qM11_c14, qM11_c15, qM11_c16, qM11_c17, qM11_c18, qM11_c19 :  std_logic_vector(1 downto 0);
signal qP10_c13, qP10_c14, qP10_c15, qP10_c16, qP10_c17, qP10_c18, qP10_c19 :  std_logic_vector(1 downto 0);
signal qM10_c13, qM10_c14, qM10_c15, qM10_c16, qM10_c17, qM10_c18, qM10_c19 :  std_logic_vector(1 downto 0);
signal qP9_c13, qP9_c14, qP9_c15, qP9_c16, qP9_c17, qP9_c18, qP9_c19 :  std_logic_vector(1 downto 0);
signal qM9_c13, qM9_c14, qM9_c15, qM9_c16, qM9_c17, qM9_c18, qM9_c19 :  std_logic_vector(1 downto 0);
signal qP8_c14, qP8_c15, qP8_c16, qP8_c17, qP8_c18, qP8_c19 :  std_logic_vector(1 downto 0);
signal qM8_c14, qM8_c15, qM8_c16, qM8_c17, qM8_c18, qM8_c19 :  std_logic_vector(1 downto 0);
signal qP7_c15, qP7_c16, qP7_c17, qP7_c18, qP7_c19 :  std_logic_vector(1 downto 0);
signal qM7_c15, qM7_c16, qM7_c17, qM7_c18, qM7_c19 :  std_logic_vector(1 downto 0);
signal qP6_c15, qP6_c16, qP6_c17, qP6_c18, qP6_c19 :  std_logic_vector(1 downto 0);
signal qM6_c15, qM6_c16, qM6_c17, qM6_c18, qM6_c19 :  std_logic_vector(1 downto 0);
signal qP5_c16, qP5_c17, qP5_c18, qP5_c19 :  std_logic_vector(1 downto 0);
signal qM5_c16, qM5_c17, qM5_c18, qM5_c19 :  std_logic_vector(1 downto 0);
signal qP4_c17, qP4_c18, qP4_c19 :  std_logic_vector(1 downto 0);
signal qM4_c17, qM4_c18, qM4_c19 :  std_logic_vector(1 downto 0);
signal qP3_c18, qP3_c19 :  std_logic_vector(1 downto 0);
signal qM3_c18, qM3_c19 :  std_logic_vector(1 downto 0);
signal qP2_c18, qP2_c19 :  std_logic_vector(1 downto 0);
signal qM2_c18, qM2_c19 :  std_logic_vector(1 downto 0);
signal qP1_c19 :  std_logic_vector(1 downto 0);
signal qM1_c19 :  std_logic_vector(1 downto 0);
signal qP_c19, qP_c20 :  std_logic_vector(55 downto 0);
signal qM_c19, qM_c20 :  std_logic_vector(55 downto 0);
signal quotient_c20 :  std_logic_vector(55 downto 0);
signal mR_c20 :  std_logic_vector(54 downto 0);
signal fRnorm_c20 :  std_logic_vector(52 downto 0);
signal round_c20 :  std_logic;
signal expR1_c20 :  std_logic_vector(12 downto 0);
signal expfrac_c20 :  std_logic_vector(64 downto 0);
signal expfracR_c20 :  std_logic_vector(64 downto 0);
signal exnR_c20 :  std_logic_vector(1 downto 0);
signal exnRfinal_c20 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               expR0_c1 <= expR0_c0;
               sR_c1 <= sR_c0;
               exnR0_c1 <= exnR0_c0;
               D_c1 <= D_c0;
               betaw27_c1 <= betaw27_c0;
               q27_c1 <= q27_c0;
               absq27D_c1 <= absq27D_c0;
               qP28_c1 <= qP28_c0;
               qM28_c1 <= qM28_c0;
               qP27_c1 <= qP27_c0;
               qM27_c1 <= qM27_c0;
            end if;
            if ce_2 = '1' then
               expR0_c2 <= expR0_c1;
               sR_c2 <= sR_c1;
               exnR0_c2 <= exnR0_c1;
               D_c2 <= D_c1;
               betaw26_c2 <= betaw26_c1;
               q26_c2 <= q26_c1;
               absq26D_c2 <= absq26D_c1;
               qP28_c2 <= qP28_c1;
               qM28_c2 <= qM28_c1;
               qP27_c2 <= qP27_c1;
               qM27_c2 <= qM27_c1;
               qP26_c2 <= qP26_c1;
               qM26_c2 <= qM26_c1;
            end if;
            if ce_3 = '1' then
               expR0_c3 <= expR0_c2;
               sR_c3 <= sR_c2;
               exnR0_c3 <= exnR0_c2;
               D_c3 <= D_c2;
               betaw24_c3 <= betaw24_c2;
               q24_copy9_c3 <= q24_copy9_c2;
               qP28_c3 <= qP28_c2;
               qM28_c3 <= qM28_c2;
               qP27_c3 <= qP27_c2;
               qM27_c3 <= qM27_c2;
               qP26_c3 <= qP26_c2;
               qM26_c3 <= qM26_c2;
               qP25_c3 <= qP25_c2;
               qM25_c3 <= qM25_c2;
            end if;
            if ce_4 = '1' then
               expR0_c4 <= expR0_c3;
               sR_c4 <= sR_c3;
               exnR0_c4 <= exnR0_c3;
               D_c4 <= D_c3;
               betaw23_c4 <= betaw23_c3;
               q23_c4 <= q23_c3;
               absq23D_c4 <= absq23D_c3;
               qP28_c4 <= qP28_c3;
               qM28_c4 <= qM28_c3;
               qP27_c4 <= qP27_c3;
               qM27_c4 <= qM27_c3;
               qP26_c4 <= qP26_c3;
               qM26_c4 <= qM26_c3;
               qP25_c4 <= qP25_c3;
               qM25_c4 <= qM25_c3;
               qP24_c4 <= qP24_c3;
               qM24_c4 <= qM24_c3;
               qP23_c4 <= qP23_c3;
               qM23_c4 <= qM23_c3;
            end if;
            if ce_5 = '1' then
               expR0_c5 <= expR0_c4;
               sR_c5 <= sR_c4;
               exnR0_c5 <= exnR0_c4;
               D_c5 <= D_c4;
               betaw21_c5 <= betaw21_c4;
               q21_copy12_c5 <= q21_copy12_c4;
               qP28_c5 <= qP28_c4;
               qM28_c5 <= qM28_c4;
               qP27_c5 <= qP27_c4;
               qM27_c5 <= qM27_c4;
               qP26_c5 <= qP26_c4;
               qM26_c5 <= qM26_c4;
               qP25_c5 <= qP25_c4;
               qM25_c5 <= qM25_c4;
               qP24_c5 <= qP24_c4;
               qM24_c5 <= qM24_c4;
               qP23_c5 <= qP23_c4;
               qM23_c5 <= qM23_c4;
               qP22_c5 <= qP22_c4;
               qM22_c5 <= qM22_c4;
            end if;
            if ce_6 = '1' then
               expR0_c6 <= expR0_c5;
               sR_c6 <= sR_c5;
               exnR0_c6 <= exnR0_c5;
               D_c6 <= D_c5;
               betaw20_c6 <= betaw20_c5;
               q20_c6 <= q20_c5;
               absq20D_c6 <= absq20D_c5;
               qP28_c6 <= qP28_c5;
               qM28_c6 <= qM28_c5;
               qP27_c6 <= qP27_c5;
               qM27_c6 <= qM27_c5;
               qP26_c6 <= qP26_c5;
               qM26_c6 <= qM26_c5;
               qP25_c6 <= qP25_c5;
               qM25_c6 <= qM25_c5;
               qP24_c6 <= qP24_c5;
               qM24_c6 <= qM24_c5;
               qP23_c6 <= qP23_c5;
               qM23_c6 <= qM23_c5;
               qP22_c6 <= qP22_c5;
               qM22_c6 <= qM22_c5;
               qP21_c6 <= qP21_c5;
               qM21_c6 <= qM21_c5;
               qP20_c6 <= qP20_c5;
               qM20_c6 <= qM20_c5;
            end if;
            if ce_7 = '1' then
               expR0_c7 <= expR0_c6;
               sR_c7 <= sR_c6;
               exnR0_c7 <= exnR0_c6;
               D_c7 <= D_c6;
               betaw19_c7 <= betaw19_c6;
               q19_c7 <= q19_c6;
               absq19D_c7 <= absq19D_c6;
               qP28_c7 <= qP28_c6;
               qM28_c7 <= qM28_c6;
               qP27_c7 <= qP27_c6;
               qM27_c7 <= qM27_c6;
               qP26_c7 <= qP26_c6;
               qM26_c7 <= qM26_c6;
               qP25_c7 <= qP25_c6;
               qM25_c7 <= qM25_c6;
               qP24_c7 <= qP24_c6;
               qM24_c7 <= qM24_c6;
               qP23_c7 <= qP23_c6;
               qM23_c7 <= qM23_c6;
               qP22_c7 <= qP22_c6;
               qM22_c7 <= qM22_c6;
               qP21_c7 <= qP21_c6;
               qM21_c7 <= qM21_c6;
               qP20_c7 <= qP20_c6;
               qM20_c7 <= qM20_c6;
               qP19_c7 <= qP19_c6;
               qM19_c7 <= qM19_c6;
            end if;
            if ce_8 = '1' then
               expR0_c8 <= expR0_c7;
               sR_c8 <= sR_c7;
               exnR0_c8 <= exnR0_c7;
               D_c8 <= D_c7;
               betaw17_c8 <= betaw17_c7;
               q17_copy16_c8 <= q17_copy16_c7;
               qP28_c8 <= qP28_c7;
               qM28_c8 <= qM28_c7;
               qP27_c8 <= qP27_c7;
               qM27_c8 <= qM27_c7;
               qP26_c8 <= qP26_c7;
               qM26_c8 <= qM26_c7;
               qP25_c8 <= qP25_c7;
               qM25_c8 <= qM25_c7;
               qP24_c8 <= qP24_c7;
               qM24_c8 <= qM24_c7;
               qP23_c8 <= qP23_c7;
               qM23_c8 <= qM23_c7;
               qP22_c8 <= qP22_c7;
               qM22_c8 <= qM22_c7;
               qP21_c8 <= qP21_c7;
               qM21_c8 <= qM21_c7;
               qP20_c8 <= qP20_c7;
               qM20_c8 <= qM20_c7;
               qP19_c8 <= qP19_c7;
               qM19_c8 <= qM19_c7;
               qP18_c8 <= qP18_c7;
               qM18_c8 <= qM18_c7;
            end if;
            if ce_9 = '1' then
               expR0_c9 <= expR0_c8;
               sR_c9 <= sR_c8;
               exnR0_c9 <= exnR0_c8;
               D_c9 <= D_c8;
               betaw16_c9 <= betaw16_c8;
               q16_c9 <= q16_c8;
               absq16D_c9 <= absq16D_c8;
               qP28_c9 <= qP28_c8;
               qM28_c9 <= qM28_c8;
               qP27_c9 <= qP27_c8;
               qM27_c9 <= qM27_c8;
               qP26_c9 <= qP26_c8;
               qM26_c9 <= qM26_c8;
               qP25_c9 <= qP25_c8;
               qM25_c9 <= qM25_c8;
               qP24_c9 <= qP24_c8;
               qM24_c9 <= qM24_c8;
               qP23_c9 <= qP23_c8;
               qM23_c9 <= qM23_c8;
               qP22_c9 <= qP22_c8;
               qM22_c9 <= qM22_c8;
               qP21_c9 <= qP21_c8;
               qM21_c9 <= qM21_c8;
               qP20_c9 <= qP20_c8;
               qM20_c9 <= qM20_c8;
               qP19_c9 <= qP19_c8;
               qM19_c9 <= qM19_c8;
               qP18_c9 <= qP18_c8;
               qM18_c9 <= qM18_c8;
               qP17_c9 <= qP17_c8;
               qM17_c9 <= qM17_c8;
               qP16_c9 <= qP16_c8;
               qM16_c9 <= qM16_c8;
            end if;
            if ce_10 = '1' then
               expR0_c10 <= expR0_c9;
               sR_c10 <= sR_c9;
               exnR0_c10 <= exnR0_c9;
               D_c10 <= D_c9;
               betaw14_c10 <= betaw14_c9;
               q14_copy19_c10 <= q14_copy19_c9;
               qP28_c10 <= qP28_c9;
               qM28_c10 <= qM28_c9;
               qP27_c10 <= qP27_c9;
               qM27_c10 <= qM27_c9;
               qP26_c10 <= qP26_c9;
               qM26_c10 <= qM26_c9;
               qP25_c10 <= qP25_c9;
               qM25_c10 <= qM25_c9;
               qP24_c10 <= qP24_c9;
               qM24_c10 <= qM24_c9;
               qP23_c10 <= qP23_c9;
               qM23_c10 <= qM23_c9;
               qP22_c10 <= qP22_c9;
               qM22_c10 <= qM22_c9;
               qP21_c10 <= qP21_c9;
               qM21_c10 <= qM21_c9;
               qP20_c10 <= qP20_c9;
               qM20_c10 <= qM20_c9;
               qP19_c10 <= qP19_c9;
               qM19_c10 <= qM19_c9;
               qP18_c10 <= qP18_c9;
               qM18_c10 <= qM18_c9;
               qP17_c10 <= qP17_c9;
               qM17_c10 <= qM17_c9;
               qP16_c10 <= qP16_c9;
               qM16_c10 <= qM16_c9;
               qP15_c10 <= qP15_c9;
               qM15_c10 <= qM15_c9;
            end if;
            if ce_11 = '1' then
               expR0_c11 <= expR0_c10;
               sR_c11 <= sR_c10;
               exnR0_c11 <= exnR0_c10;
               D_c11 <= D_c10;
               betaw13_c11 <= betaw13_c10;
               q13_c11 <= q13_c10;
               absq13D_c11 <= absq13D_c10;
               qP28_c11 <= qP28_c10;
               qM28_c11 <= qM28_c10;
               qP27_c11 <= qP27_c10;
               qM27_c11 <= qM27_c10;
               qP26_c11 <= qP26_c10;
               qM26_c11 <= qM26_c10;
               qP25_c11 <= qP25_c10;
               qM25_c11 <= qM25_c10;
               qP24_c11 <= qP24_c10;
               qM24_c11 <= qM24_c10;
               qP23_c11 <= qP23_c10;
               qM23_c11 <= qM23_c10;
               qP22_c11 <= qP22_c10;
               qM22_c11 <= qM22_c10;
               qP21_c11 <= qP21_c10;
               qM21_c11 <= qM21_c10;
               qP20_c11 <= qP20_c10;
               qM20_c11 <= qM20_c10;
               qP19_c11 <= qP19_c10;
               qM19_c11 <= qM19_c10;
               qP18_c11 <= qP18_c10;
               qM18_c11 <= qM18_c10;
               qP17_c11 <= qP17_c10;
               qM17_c11 <= qM17_c10;
               qP16_c11 <= qP16_c10;
               qM16_c11 <= qM16_c10;
               qP15_c11 <= qP15_c10;
               qM15_c11 <= qM15_c10;
               qP14_c11 <= qP14_c10;
               qM14_c11 <= qM14_c10;
               qP13_c11 <= qP13_c10;
               qM13_c11 <= qM13_c10;
            end if;
            if ce_12 = '1' then
               expR0_c12 <= expR0_c11;
               sR_c12 <= sR_c11;
               exnR0_c12 <= exnR0_c11;
               D_c12 <= D_c11;
               betaw12_c12 <= betaw12_c11;
               q12_c12 <= q12_c11;
               absq12D_c12 <= absq12D_c11;
               qP28_c12 <= qP28_c11;
               qM28_c12 <= qM28_c11;
               qP27_c12 <= qP27_c11;
               qM27_c12 <= qM27_c11;
               qP26_c12 <= qP26_c11;
               qM26_c12 <= qM26_c11;
               qP25_c12 <= qP25_c11;
               qM25_c12 <= qM25_c11;
               qP24_c12 <= qP24_c11;
               qM24_c12 <= qM24_c11;
               qP23_c12 <= qP23_c11;
               qM23_c12 <= qM23_c11;
               qP22_c12 <= qP22_c11;
               qM22_c12 <= qM22_c11;
               qP21_c12 <= qP21_c11;
               qM21_c12 <= qM21_c11;
               qP20_c12 <= qP20_c11;
               qM20_c12 <= qM20_c11;
               qP19_c12 <= qP19_c11;
               qM19_c12 <= qM19_c11;
               qP18_c12 <= qP18_c11;
               qM18_c12 <= qM18_c11;
               qP17_c12 <= qP17_c11;
               qM17_c12 <= qM17_c11;
               qP16_c12 <= qP16_c11;
               qM16_c12 <= qM16_c11;
               qP15_c12 <= qP15_c11;
               qM15_c12 <= qM15_c11;
               qP14_c12 <= qP14_c11;
               qM14_c12 <= qM14_c11;
               qP13_c12 <= qP13_c11;
               qM13_c12 <= qM13_c11;
               qP12_c12 <= qP12_c11;
               qM12_c12 <= qM12_c11;
            end if;
            if ce_13 = '1' then
               expR0_c13 <= expR0_c12;
               sR_c13 <= sR_c12;
               exnR0_c13 <= exnR0_c12;
               D_c13 <= D_c12;
               betaw10_c13 <= betaw10_c12;
               q10_copy23_c13 <= q10_copy23_c12;
               qP28_c13 <= qP28_c12;
               qM28_c13 <= qM28_c12;
               qP27_c13 <= qP27_c12;
               qM27_c13 <= qM27_c12;
               qP26_c13 <= qP26_c12;
               qM26_c13 <= qM26_c12;
               qP25_c13 <= qP25_c12;
               qM25_c13 <= qM25_c12;
               qP24_c13 <= qP24_c12;
               qM24_c13 <= qM24_c12;
               qP23_c13 <= qP23_c12;
               qM23_c13 <= qM23_c12;
               qP22_c13 <= qP22_c12;
               qM22_c13 <= qM22_c12;
               qP21_c13 <= qP21_c12;
               qM21_c13 <= qM21_c12;
               qP20_c13 <= qP20_c12;
               qM20_c13 <= qM20_c12;
               qP19_c13 <= qP19_c12;
               qM19_c13 <= qM19_c12;
               qP18_c13 <= qP18_c12;
               qM18_c13 <= qM18_c12;
               qP17_c13 <= qP17_c12;
               qM17_c13 <= qM17_c12;
               qP16_c13 <= qP16_c12;
               qM16_c13 <= qM16_c12;
               qP15_c13 <= qP15_c12;
               qM15_c13 <= qM15_c12;
               qP14_c13 <= qP14_c12;
               qM14_c13 <= qM14_c12;
               qP13_c13 <= qP13_c12;
               qM13_c13 <= qM13_c12;
               qP12_c13 <= qP12_c12;
               qM12_c13 <= qM12_c12;
               qP11_c13 <= qP11_c12;
               qM11_c13 <= qM11_c12;
            end if;
            if ce_14 = '1' then
               expR0_c14 <= expR0_c13;
               sR_c14 <= sR_c13;
               exnR0_c14 <= exnR0_c13;
               D_c14 <= D_c13;
               betaw9_c14 <= betaw9_c13;
               q9_c14 <= q9_c13;
               absq9D_c14 <= absq9D_c13;
               qP28_c14 <= qP28_c13;
               qM28_c14 <= qM28_c13;
               qP27_c14 <= qP27_c13;
               qM27_c14 <= qM27_c13;
               qP26_c14 <= qP26_c13;
               qM26_c14 <= qM26_c13;
               qP25_c14 <= qP25_c13;
               qM25_c14 <= qM25_c13;
               qP24_c14 <= qP24_c13;
               qM24_c14 <= qM24_c13;
               qP23_c14 <= qP23_c13;
               qM23_c14 <= qM23_c13;
               qP22_c14 <= qP22_c13;
               qM22_c14 <= qM22_c13;
               qP21_c14 <= qP21_c13;
               qM21_c14 <= qM21_c13;
               qP20_c14 <= qP20_c13;
               qM20_c14 <= qM20_c13;
               qP19_c14 <= qP19_c13;
               qM19_c14 <= qM19_c13;
               qP18_c14 <= qP18_c13;
               qM18_c14 <= qM18_c13;
               qP17_c14 <= qP17_c13;
               qM17_c14 <= qM17_c13;
               qP16_c14 <= qP16_c13;
               qM16_c14 <= qM16_c13;
               qP15_c14 <= qP15_c13;
               qM15_c14 <= qM15_c13;
               qP14_c14 <= qP14_c13;
               qM14_c14 <= qM14_c13;
               qP13_c14 <= qP13_c13;
               qM13_c14 <= qM13_c13;
               qP12_c14 <= qP12_c13;
               qM12_c14 <= qM12_c13;
               qP11_c14 <= qP11_c13;
               qM11_c14 <= qM11_c13;
               qP10_c14 <= qP10_c13;
               qM10_c14 <= qM10_c13;
               qP9_c14 <= qP9_c13;
               qM9_c14 <= qM9_c13;
            end if;
            if ce_15 = '1' then
               expR0_c15 <= expR0_c14;
               sR_c15 <= sR_c14;
               exnR0_c15 <= exnR0_c14;
               D_c15 <= D_c14;
               betaw7_c15 <= betaw7_c14;
               q7_copy26_c15 <= q7_copy26_c14;
               qP28_c15 <= qP28_c14;
               qM28_c15 <= qM28_c14;
               qP27_c15 <= qP27_c14;
               qM27_c15 <= qM27_c14;
               qP26_c15 <= qP26_c14;
               qM26_c15 <= qM26_c14;
               qP25_c15 <= qP25_c14;
               qM25_c15 <= qM25_c14;
               qP24_c15 <= qP24_c14;
               qM24_c15 <= qM24_c14;
               qP23_c15 <= qP23_c14;
               qM23_c15 <= qM23_c14;
               qP22_c15 <= qP22_c14;
               qM22_c15 <= qM22_c14;
               qP21_c15 <= qP21_c14;
               qM21_c15 <= qM21_c14;
               qP20_c15 <= qP20_c14;
               qM20_c15 <= qM20_c14;
               qP19_c15 <= qP19_c14;
               qM19_c15 <= qM19_c14;
               qP18_c15 <= qP18_c14;
               qM18_c15 <= qM18_c14;
               qP17_c15 <= qP17_c14;
               qM17_c15 <= qM17_c14;
               qP16_c15 <= qP16_c14;
               qM16_c15 <= qM16_c14;
               qP15_c15 <= qP15_c14;
               qM15_c15 <= qM15_c14;
               qP14_c15 <= qP14_c14;
               qM14_c15 <= qM14_c14;
               qP13_c15 <= qP13_c14;
               qM13_c15 <= qM13_c14;
               qP12_c15 <= qP12_c14;
               qM12_c15 <= qM12_c14;
               qP11_c15 <= qP11_c14;
               qM11_c15 <= qM11_c14;
               qP10_c15 <= qP10_c14;
               qM10_c15 <= qM10_c14;
               qP9_c15 <= qP9_c14;
               qM9_c15 <= qM9_c14;
               qP8_c15 <= qP8_c14;
               qM8_c15 <= qM8_c14;
            end if;
            if ce_16 = '1' then
               expR0_c16 <= expR0_c15;
               sR_c16 <= sR_c15;
               exnR0_c16 <= exnR0_c15;
               D_c16 <= D_c15;
               betaw6_c16 <= betaw6_c15;
               q6_c16 <= q6_c15;
               absq6D_c16 <= absq6D_c15;
               qP28_c16 <= qP28_c15;
               qM28_c16 <= qM28_c15;
               qP27_c16 <= qP27_c15;
               qM27_c16 <= qM27_c15;
               qP26_c16 <= qP26_c15;
               qM26_c16 <= qM26_c15;
               qP25_c16 <= qP25_c15;
               qM25_c16 <= qM25_c15;
               qP24_c16 <= qP24_c15;
               qM24_c16 <= qM24_c15;
               qP23_c16 <= qP23_c15;
               qM23_c16 <= qM23_c15;
               qP22_c16 <= qP22_c15;
               qM22_c16 <= qM22_c15;
               qP21_c16 <= qP21_c15;
               qM21_c16 <= qM21_c15;
               qP20_c16 <= qP20_c15;
               qM20_c16 <= qM20_c15;
               qP19_c16 <= qP19_c15;
               qM19_c16 <= qM19_c15;
               qP18_c16 <= qP18_c15;
               qM18_c16 <= qM18_c15;
               qP17_c16 <= qP17_c15;
               qM17_c16 <= qM17_c15;
               qP16_c16 <= qP16_c15;
               qM16_c16 <= qM16_c15;
               qP15_c16 <= qP15_c15;
               qM15_c16 <= qM15_c15;
               qP14_c16 <= qP14_c15;
               qM14_c16 <= qM14_c15;
               qP13_c16 <= qP13_c15;
               qM13_c16 <= qM13_c15;
               qP12_c16 <= qP12_c15;
               qM12_c16 <= qM12_c15;
               qP11_c16 <= qP11_c15;
               qM11_c16 <= qM11_c15;
               qP10_c16 <= qP10_c15;
               qM10_c16 <= qM10_c15;
               qP9_c16 <= qP9_c15;
               qM9_c16 <= qM9_c15;
               qP8_c16 <= qP8_c15;
               qM8_c16 <= qM8_c15;
               qP7_c16 <= qP7_c15;
               qM7_c16 <= qM7_c15;
               qP6_c16 <= qP6_c15;
               qM6_c16 <= qM6_c15;
            end if;
            if ce_17 = '1' then
               expR0_c17 <= expR0_c16;
               sR_c17 <= sR_c16;
               exnR0_c17 <= exnR0_c16;
               D_c17 <= D_c16;
               betaw5_c17 <= betaw5_c16;
               q5_c17 <= q5_c16;
               absq5D_c17 <= absq5D_c16;
               qP28_c17 <= qP28_c16;
               qM28_c17 <= qM28_c16;
               qP27_c17 <= qP27_c16;
               qM27_c17 <= qM27_c16;
               qP26_c17 <= qP26_c16;
               qM26_c17 <= qM26_c16;
               qP25_c17 <= qP25_c16;
               qM25_c17 <= qM25_c16;
               qP24_c17 <= qP24_c16;
               qM24_c17 <= qM24_c16;
               qP23_c17 <= qP23_c16;
               qM23_c17 <= qM23_c16;
               qP22_c17 <= qP22_c16;
               qM22_c17 <= qM22_c16;
               qP21_c17 <= qP21_c16;
               qM21_c17 <= qM21_c16;
               qP20_c17 <= qP20_c16;
               qM20_c17 <= qM20_c16;
               qP19_c17 <= qP19_c16;
               qM19_c17 <= qM19_c16;
               qP18_c17 <= qP18_c16;
               qM18_c17 <= qM18_c16;
               qP17_c17 <= qP17_c16;
               qM17_c17 <= qM17_c16;
               qP16_c17 <= qP16_c16;
               qM16_c17 <= qM16_c16;
               qP15_c17 <= qP15_c16;
               qM15_c17 <= qM15_c16;
               qP14_c17 <= qP14_c16;
               qM14_c17 <= qM14_c16;
               qP13_c17 <= qP13_c16;
               qM13_c17 <= qM13_c16;
               qP12_c17 <= qP12_c16;
               qM12_c17 <= qM12_c16;
               qP11_c17 <= qP11_c16;
               qM11_c17 <= qM11_c16;
               qP10_c17 <= qP10_c16;
               qM10_c17 <= qM10_c16;
               qP9_c17 <= qP9_c16;
               qM9_c17 <= qM9_c16;
               qP8_c17 <= qP8_c16;
               qM8_c17 <= qM8_c16;
               qP7_c17 <= qP7_c16;
               qM7_c17 <= qM7_c16;
               qP6_c17 <= qP6_c16;
               qM6_c17 <= qM6_c16;
               qP5_c17 <= qP5_c16;
               qM5_c17 <= qM5_c16;
            end if;
            if ce_18 = '1' then
               expR0_c18 <= expR0_c17;
               sR_c18 <= sR_c17;
               exnR0_c18 <= exnR0_c17;
               D_c18 <= D_c17;
               betaw3_c18 <= betaw3_c17;
               q3_copy30_c18 <= q3_copy30_c17;
               qP28_c18 <= qP28_c17;
               qM28_c18 <= qM28_c17;
               qP27_c18 <= qP27_c17;
               qM27_c18 <= qM27_c17;
               qP26_c18 <= qP26_c17;
               qM26_c18 <= qM26_c17;
               qP25_c18 <= qP25_c17;
               qM25_c18 <= qM25_c17;
               qP24_c18 <= qP24_c17;
               qM24_c18 <= qM24_c17;
               qP23_c18 <= qP23_c17;
               qM23_c18 <= qM23_c17;
               qP22_c18 <= qP22_c17;
               qM22_c18 <= qM22_c17;
               qP21_c18 <= qP21_c17;
               qM21_c18 <= qM21_c17;
               qP20_c18 <= qP20_c17;
               qM20_c18 <= qM20_c17;
               qP19_c18 <= qP19_c17;
               qM19_c18 <= qM19_c17;
               qP18_c18 <= qP18_c17;
               qM18_c18 <= qM18_c17;
               qP17_c18 <= qP17_c17;
               qM17_c18 <= qM17_c17;
               qP16_c18 <= qP16_c17;
               qM16_c18 <= qM16_c17;
               qP15_c18 <= qP15_c17;
               qM15_c18 <= qM15_c17;
               qP14_c18 <= qP14_c17;
               qM14_c18 <= qM14_c17;
               qP13_c18 <= qP13_c17;
               qM13_c18 <= qM13_c17;
               qP12_c18 <= qP12_c17;
               qM12_c18 <= qM12_c17;
               qP11_c18 <= qP11_c17;
               qM11_c18 <= qM11_c17;
               qP10_c18 <= qP10_c17;
               qM10_c18 <= qM10_c17;
               qP9_c18 <= qP9_c17;
               qM9_c18 <= qM9_c17;
               qP8_c18 <= qP8_c17;
               qM8_c18 <= qM8_c17;
               qP7_c18 <= qP7_c17;
               qM7_c18 <= qM7_c17;
               qP6_c18 <= qP6_c17;
               qM6_c18 <= qM6_c17;
               qP5_c18 <= qP5_c17;
               qM5_c18 <= qM5_c17;
               qP4_c18 <= qP4_c17;
               qM4_c18 <= qM4_c17;
            end if;
            if ce_19 = '1' then
               expR0_c19 <= expR0_c18;
               sR_c19 <= sR_c18;
               exnR0_c19 <= exnR0_c18;
               D_c19 <= D_c18;
               betaw2_c19 <= betaw2_c18;
               q2_c19 <= q2_c18;
               absq2D_c19 <= absq2D_c18;
               qP28_c19 <= qP28_c18;
               qM28_c19 <= qM28_c18;
               qP27_c19 <= qP27_c18;
               qM27_c19 <= qM27_c18;
               qP26_c19 <= qP26_c18;
               qM26_c19 <= qM26_c18;
               qP25_c19 <= qP25_c18;
               qM25_c19 <= qM25_c18;
               qP24_c19 <= qP24_c18;
               qM24_c19 <= qM24_c18;
               qP23_c19 <= qP23_c18;
               qM23_c19 <= qM23_c18;
               qP22_c19 <= qP22_c18;
               qM22_c19 <= qM22_c18;
               qP21_c19 <= qP21_c18;
               qM21_c19 <= qM21_c18;
               qP20_c19 <= qP20_c18;
               qM20_c19 <= qM20_c18;
               qP19_c19 <= qP19_c18;
               qM19_c19 <= qM19_c18;
               qP18_c19 <= qP18_c18;
               qM18_c19 <= qM18_c18;
               qP17_c19 <= qP17_c18;
               qM17_c19 <= qM17_c18;
               qP16_c19 <= qP16_c18;
               qM16_c19 <= qM16_c18;
               qP15_c19 <= qP15_c18;
               qM15_c19 <= qM15_c18;
               qP14_c19 <= qP14_c18;
               qM14_c19 <= qM14_c18;
               qP13_c19 <= qP13_c18;
               qM13_c19 <= qM13_c18;
               qP12_c19 <= qP12_c18;
               qM12_c19 <= qM12_c18;
               qP11_c19 <= qP11_c18;
               qM11_c19 <= qM11_c18;
               qP10_c19 <= qP10_c18;
               qM10_c19 <= qM10_c18;
               qP9_c19 <= qP9_c18;
               qM9_c19 <= qM9_c18;
               qP8_c19 <= qP8_c18;
               qM8_c19 <= qM8_c18;
               qP7_c19 <= qP7_c18;
               qM7_c19 <= qM7_c18;
               qP6_c19 <= qP6_c18;
               qM6_c19 <= qM6_c18;
               qP5_c19 <= qP5_c18;
               qM5_c19 <= qM5_c18;
               qP4_c19 <= qP4_c18;
               qM4_c19 <= qM4_c18;
               qP3_c19 <= qP3_c18;
               qM3_c19 <= qM3_c18;
               qP2_c19 <= qP2_c18;
               qM2_c19 <= qM2_c18;
            end if;
            if ce_20 = '1' then
               expR0_c20 <= expR0_c19;
               sR_c20 <= sR_c19;
               exnR0_c20 <= exnR0_c19;
               qP_c20 <= qP_c19;
               qM_c20 <= qM_c19;
            end if;
         end if;
      end process;
   fX_c0 <= "1" & X(51 downto 0);
   fY_c0 <= "1" & Y(51 downto 0);
   -- exponent difference, sign and exception combination computed early, to have fewer bits to pipeline
   expR0_c0 <= ("00" & X(62 downto 52)) - ("00" & Y(62 downto 52));
   sR_c0 <= X(63) xor Y(63);
   -- early exception handling 
   exnXY_c0 <= X(65 downto 64) & Y(65 downto 64);
   with exnXY_c0  select 
      exnR0_c0 <= 
         "01"	 when "0101",										-- normal
         "00"	 when "0001" | "0010" | "0110", -- zero
         "10"	 when "0100" | "1000" | "1001", -- overflow
         "11"	 when others;										-- NaN
   D_c0 <= fY_c0 ;
   psX_c0 <= "0" & fX_c0 ;
   betaw28_c0 <=  "00" & psX_c0;
   sel28_c0 <= betaw28_c0(55 downto 50) & D_c0(51 downto 49);
   SelFunctionTable28: selFunction_Freq300_uid4
      port map ( X => sel28_c0,
                 Y => q28_copy5_c0);
   q28_c0 <= q28_copy5_c0; -- output copy to hold a pipeline register if needed

   with q28_c0  select 
      absq28D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q28_c0(2)  select 
   w27_c0<= betaw28_c0 - absq28D_c0 when '0',
         betaw28_c0 + absq28D_c0 when others;

   betaw27_c0 <= w27_c0(53 downto 0) & "00"; -- multiplication by the radix
   sel27_c0 <= betaw27_c0(55 downto 50) & D_c0(51 downto 49);
   SelFunctionTable27: selFunction_Freq300_uid4
      port map ( X => sel27_c0,
                 Y => q27_copy6_c0);
   q27_c0 <= q27_copy6_c0; -- output copy to hold a pipeline register if needed

   with q27_c0  select 
      absq27D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q27_c1(2)  select 
   w26_c1<= betaw27_c1 - absq27D_c1 when '0',
         betaw27_c1 + absq27D_c1 when others;

   betaw26_c1 <= w26_c1(53 downto 0) & "00"; -- multiplication by the radix
   sel26_c1 <= betaw26_c1(55 downto 50) & D_c1(51 downto 49);
   SelFunctionTable26: selFunction_Freq300_uid4
      port map ( X => sel26_c1,
                 Y => q26_copy7_c1);
   q26_c1 <= q26_copy7_c1; -- output copy to hold a pipeline register if needed

   with q26_c1  select 
      absq26D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q26_c2(2)  select 
   w25_c2<= betaw26_c2 - absq26D_c2 when '0',
         betaw26_c2 + absq26D_c2 when others;

   betaw25_c2 <= w25_c2(53 downto 0) & "00"; -- multiplication by the radix
   sel25_c2 <= betaw25_c2(55 downto 50) & D_c2(51 downto 49);
   SelFunctionTable25: selFunction_Freq300_uid4
      port map ( X => sel25_c2,
                 Y => q25_copy8_c2);
   q25_c2 <= q25_copy8_c2; -- output copy to hold a pipeline register if needed

   with q25_c2  select 
      absq25D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q25_c2(2)  select 
   w24_c2<= betaw25_c2 - absq25D_c2 when '0',
         betaw25_c2 + absq25D_c2 when others;

   betaw24_c2 <= w24_c2(53 downto 0) & "00"; -- multiplication by the radix
   sel24_c2 <= betaw24_c2(55 downto 50) & D_c2(51 downto 49);
   SelFunctionTable24: selFunction_Freq300_uid4
      port map ( X => sel24_c2,
                 Y => q24_copy9_c2);
   q24_c3 <= q24_copy9_c3; -- output copy to hold a pipeline register if needed

   with q24_c3  select 
      absq24D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q24_c3(2)  select 
   w23_c3<= betaw24_c3 - absq24D_c3 when '0',
         betaw24_c3 + absq24D_c3 when others;

   betaw23_c3 <= w23_c3(53 downto 0) & "00"; -- multiplication by the radix
   sel23_c3 <= betaw23_c3(55 downto 50) & D_c3(51 downto 49);
   SelFunctionTable23: selFunction_Freq300_uid4
      port map ( X => sel23_c3,
                 Y => q23_copy10_c3);
   q23_c3 <= q23_copy10_c3; -- output copy to hold a pipeline register if needed

   with q23_c3  select 
      absq23D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q23_c4(2)  select 
   w22_c4<= betaw23_c4 - absq23D_c4 when '0',
         betaw23_c4 + absq23D_c4 when others;

   betaw22_c4 <= w22_c4(53 downto 0) & "00"; -- multiplication by the radix
   sel22_c4 <= betaw22_c4(55 downto 50) & D_c4(51 downto 49);
   SelFunctionTable22: selFunction_Freq300_uid4
      port map ( X => sel22_c4,
                 Y => q22_copy11_c4);
   q22_c4 <= q22_copy11_c4; -- output copy to hold a pipeline register if needed

   with q22_c4  select 
      absq22D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q22_c4(2)  select 
   w21_c4<= betaw22_c4 - absq22D_c4 when '0',
         betaw22_c4 + absq22D_c4 when others;

   betaw21_c4 <= w21_c4(53 downto 0) & "00"; -- multiplication by the radix
   sel21_c4 <= betaw21_c4(55 downto 50) & D_c4(51 downto 49);
   SelFunctionTable21: selFunction_Freq300_uid4
      port map ( X => sel21_c4,
                 Y => q21_copy12_c4);
   q21_c5 <= q21_copy12_c5; -- output copy to hold a pipeline register if needed

   with q21_c5  select 
      absq21D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q21_c5(2)  select 
   w20_c5<= betaw21_c5 - absq21D_c5 when '0',
         betaw21_c5 + absq21D_c5 when others;

   betaw20_c5 <= w20_c5(53 downto 0) & "00"; -- multiplication by the radix
   sel20_c5 <= betaw20_c5(55 downto 50) & D_c5(51 downto 49);
   SelFunctionTable20: selFunction_Freq300_uid4
      port map ( X => sel20_c5,
                 Y => q20_copy13_c5);
   q20_c5 <= q20_copy13_c5; -- output copy to hold a pipeline register if needed

   with q20_c5  select 
      absq20D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q20_c6(2)  select 
   w19_c6<= betaw20_c6 - absq20D_c6 when '0',
         betaw20_c6 + absq20D_c6 when others;

   betaw19_c6 <= w19_c6(53 downto 0) & "00"; -- multiplication by the radix
   sel19_c6 <= betaw19_c6(55 downto 50) & D_c6(51 downto 49);
   SelFunctionTable19: selFunction_Freq300_uid4
      port map ( X => sel19_c6,
                 Y => q19_copy14_c6);
   q19_c6 <= q19_copy14_c6; -- output copy to hold a pipeline register if needed

   with q19_c6  select 
      absq19D_c6 <= 
         "000" & D_c6						 when "001" | "111", -- mult by 1
         "00" & D_c6 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q19_c7(2)  select 
   w18_c7<= betaw19_c7 - absq19D_c7 when '0',
         betaw19_c7 + absq19D_c7 when others;

   betaw18_c7 <= w18_c7(53 downto 0) & "00"; -- multiplication by the radix
   sel18_c7 <= betaw18_c7(55 downto 50) & D_c7(51 downto 49);
   SelFunctionTable18: selFunction_Freq300_uid4
      port map ( X => sel18_c7,
                 Y => q18_copy15_c7);
   q18_c7 <= q18_copy15_c7; -- output copy to hold a pipeline register if needed

   with q18_c7  select 
      absq18D_c7 <= 
         "000" & D_c7						 when "001" | "111", -- mult by 1
         "00" & D_c7 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q18_c7(2)  select 
   w17_c7<= betaw18_c7 - absq18D_c7 when '0',
         betaw18_c7 + absq18D_c7 when others;

   betaw17_c7 <= w17_c7(53 downto 0) & "00"; -- multiplication by the radix
   sel17_c7 <= betaw17_c7(55 downto 50) & D_c7(51 downto 49);
   SelFunctionTable17: selFunction_Freq300_uid4
      port map ( X => sel17_c7,
                 Y => q17_copy16_c7);
   q17_c8 <= q17_copy16_c8; -- output copy to hold a pipeline register if needed

   with q17_c8  select 
      absq17D_c8 <= 
         "000" & D_c8						 when "001" | "111", -- mult by 1
         "00" & D_c8 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q17_c8(2)  select 
   w16_c8<= betaw17_c8 - absq17D_c8 when '0',
         betaw17_c8 + absq17D_c8 when others;

   betaw16_c8 <= w16_c8(53 downto 0) & "00"; -- multiplication by the radix
   sel16_c8 <= betaw16_c8(55 downto 50) & D_c8(51 downto 49);
   SelFunctionTable16: selFunction_Freq300_uid4
      port map ( X => sel16_c8,
                 Y => q16_copy17_c8);
   q16_c8 <= q16_copy17_c8; -- output copy to hold a pipeline register if needed

   with q16_c8  select 
      absq16D_c8 <= 
         "000" & D_c8						 when "001" | "111", -- mult by 1
         "00" & D_c8 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q16_c9(2)  select 
   w15_c9<= betaw16_c9 - absq16D_c9 when '0',
         betaw16_c9 + absq16D_c9 when others;

   betaw15_c9 <= w15_c9(53 downto 0) & "00"; -- multiplication by the radix
   sel15_c9 <= betaw15_c9(55 downto 50) & D_c9(51 downto 49);
   SelFunctionTable15: selFunction_Freq300_uid4
      port map ( X => sel15_c9,
                 Y => q15_copy18_c9);
   q15_c9 <= q15_copy18_c9; -- output copy to hold a pipeline register if needed

   with q15_c9  select 
      absq15D_c9 <= 
         "000" & D_c9						 when "001" | "111", -- mult by 1
         "00" & D_c9 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q15_c9(2)  select 
   w14_c9<= betaw15_c9 - absq15D_c9 when '0',
         betaw15_c9 + absq15D_c9 when others;

   betaw14_c9 <= w14_c9(53 downto 0) & "00"; -- multiplication by the radix
   sel14_c9 <= betaw14_c9(55 downto 50) & D_c9(51 downto 49);
   SelFunctionTable14: selFunction_Freq300_uid4
      port map ( X => sel14_c9,
                 Y => q14_copy19_c9);
   q14_c10 <= q14_copy19_c10; -- output copy to hold a pipeline register if needed

   with q14_c10  select 
      absq14D_c10 <= 
         "000" & D_c10						 when "001" | "111", -- mult by 1
         "00" & D_c10 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q14_c10(2)  select 
   w13_c10<= betaw14_c10 - absq14D_c10 when '0',
         betaw14_c10 + absq14D_c10 when others;

   betaw13_c10 <= w13_c10(53 downto 0) & "00"; -- multiplication by the radix
   sel13_c10 <= betaw13_c10(55 downto 50) & D_c10(51 downto 49);
   SelFunctionTable13: selFunction_Freq300_uid4
      port map ( X => sel13_c10,
                 Y => q13_copy20_c10);
   q13_c10 <= q13_copy20_c10; -- output copy to hold a pipeline register if needed

   with q13_c10  select 
      absq13D_c10 <= 
         "000" & D_c10						 when "001" | "111", -- mult by 1
         "00" & D_c10 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q13_c11(2)  select 
   w12_c11<= betaw13_c11 - absq13D_c11 when '0',
         betaw13_c11 + absq13D_c11 when others;

   betaw12_c11 <= w12_c11(53 downto 0) & "00"; -- multiplication by the radix
   sel12_c11 <= betaw12_c11(55 downto 50) & D_c11(51 downto 49);
   SelFunctionTable12: selFunction_Freq300_uid4
      port map ( X => sel12_c11,
                 Y => q12_copy21_c11);
   q12_c11 <= q12_copy21_c11; -- output copy to hold a pipeline register if needed

   with q12_c11  select 
      absq12D_c11 <= 
         "000" & D_c11						 when "001" | "111", -- mult by 1
         "00" & D_c11 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q12_c12(2)  select 
   w11_c12<= betaw12_c12 - absq12D_c12 when '0',
         betaw12_c12 + absq12D_c12 when others;

   betaw11_c12 <= w11_c12(53 downto 0) & "00"; -- multiplication by the radix
   sel11_c12 <= betaw11_c12(55 downto 50) & D_c12(51 downto 49);
   SelFunctionTable11: selFunction_Freq300_uid4
      port map ( X => sel11_c12,
                 Y => q11_copy22_c12);
   q11_c12 <= q11_copy22_c12; -- output copy to hold a pipeline register if needed

   with q11_c12  select 
      absq11D_c12 <= 
         "000" & D_c12						 when "001" | "111", -- mult by 1
         "00" & D_c12 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q11_c12(2)  select 
   w10_c12<= betaw11_c12 - absq11D_c12 when '0',
         betaw11_c12 + absq11D_c12 when others;

   betaw10_c12 <= w10_c12(53 downto 0) & "00"; -- multiplication by the radix
   sel10_c12 <= betaw10_c12(55 downto 50) & D_c12(51 downto 49);
   SelFunctionTable10: selFunction_Freq300_uid4
      port map ( X => sel10_c12,
                 Y => q10_copy23_c12);
   q10_c13 <= q10_copy23_c13; -- output copy to hold a pipeline register if needed

   with q10_c13  select 
      absq10D_c13 <= 
         "000" & D_c13						 when "001" | "111", -- mult by 1
         "00" & D_c13 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q10_c13(2)  select 
   w9_c13<= betaw10_c13 - absq10D_c13 when '0',
         betaw10_c13 + absq10D_c13 when others;

   betaw9_c13 <= w9_c13(53 downto 0) & "00"; -- multiplication by the radix
   sel9_c13 <= betaw9_c13(55 downto 50) & D_c13(51 downto 49);
   SelFunctionTable9: selFunction_Freq300_uid4
      port map ( X => sel9_c13,
                 Y => q9_copy24_c13);
   q9_c13 <= q9_copy24_c13; -- output copy to hold a pipeline register if needed

   with q9_c13  select 
      absq9D_c13 <= 
         "000" & D_c13						 when "001" | "111", -- mult by 1
         "00" & D_c13 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q9_c14(2)  select 
   w8_c14<= betaw9_c14 - absq9D_c14 when '0',
         betaw9_c14 + absq9D_c14 when others;

   betaw8_c14 <= w8_c14(53 downto 0) & "00"; -- multiplication by the radix
   sel8_c14 <= betaw8_c14(55 downto 50) & D_c14(51 downto 49);
   SelFunctionTable8: selFunction_Freq300_uid4
      port map ( X => sel8_c14,
                 Y => q8_copy25_c14);
   q8_c14 <= q8_copy25_c14; -- output copy to hold a pipeline register if needed

   with q8_c14  select 
      absq8D_c14 <= 
         "000" & D_c14						 when "001" | "111", -- mult by 1
         "00" & D_c14 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q8_c14(2)  select 
   w7_c14<= betaw8_c14 - absq8D_c14 when '0',
         betaw8_c14 + absq8D_c14 when others;

   betaw7_c14 <= w7_c14(53 downto 0) & "00"; -- multiplication by the radix
   sel7_c14 <= betaw7_c14(55 downto 50) & D_c14(51 downto 49);
   SelFunctionTable7: selFunction_Freq300_uid4
      port map ( X => sel7_c14,
                 Y => q7_copy26_c14);
   q7_c15 <= q7_copy26_c15; -- output copy to hold a pipeline register if needed

   with q7_c15  select 
      absq7D_c15 <= 
         "000" & D_c15						 when "001" | "111", -- mult by 1
         "00" & D_c15 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q7_c15(2)  select 
   w6_c15<= betaw7_c15 - absq7D_c15 when '0',
         betaw7_c15 + absq7D_c15 when others;

   betaw6_c15 <= w6_c15(53 downto 0) & "00"; -- multiplication by the radix
   sel6_c15 <= betaw6_c15(55 downto 50) & D_c15(51 downto 49);
   SelFunctionTable6: selFunction_Freq300_uid4
      port map ( X => sel6_c15,
                 Y => q6_copy27_c15);
   q6_c15 <= q6_copy27_c15; -- output copy to hold a pipeline register if needed

   with q6_c15  select 
      absq6D_c15 <= 
         "000" & D_c15						 when "001" | "111", -- mult by 1
         "00" & D_c15 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q6_c16(2)  select 
   w5_c16<= betaw6_c16 - absq6D_c16 when '0',
         betaw6_c16 + absq6D_c16 when others;

   betaw5_c16 <= w5_c16(53 downto 0) & "00"; -- multiplication by the radix
   sel5_c16 <= betaw5_c16(55 downto 50) & D_c16(51 downto 49);
   SelFunctionTable5: selFunction_Freq300_uid4
      port map ( X => sel5_c16,
                 Y => q5_copy28_c16);
   q5_c16 <= q5_copy28_c16; -- output copy to hold a pipeline register if needed

   with q5_c16  select 
      absq5D_c16 <= 
         "000" & D_c16						 when "001" | "111", -- mult by 1
         "00" & D_c16 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q5_c17(2)  select 
   w4_c17<= betaw5_c17 - absq5D_c17 when '0',
         betaw5_c17 + absq5D_c17 when others;

   betaw4_c17 <= w4_c17(53 downto 0) & "00"; -- multiplication by the radix
   sel4_c17 <= betaw4_c17(55 downto 50) & D_c17(51 downto 49);
   SelFunctionTable4: selFunction_Freq300_uid4
      port map ( X => sel4_c17,
                 Y => q4_copy29_c17);
   q4_c17 <= q4_copy29_c17; -- output copy to hold a pipeline register if needed

   with q4_c17  select 
      absq4D_c17 <= 
         "000" & D_c17						 when "001" | "111", -- mult by 1
         "00" & D_c17 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q4_c17(2)  select 
   w3_c17<= betaw4_c17 - absq4D_c17 when '0',
         betaw4_c17 + absq4D_c17 when others;

   betaw3_c17 <= w3_c17(53 downto 0) & "00"; -- multiplication by the radix
   sel3_c17 <= betaw3_c17(55 downto 50) & D_c17(51 downto 49);
   SelFunctionTable3: selFunction_Freq300_uid4
      port map ( X => sel3_c17,
                 Y => q3_copy30_c17);
   q3_c18 <= q3_copy30_c18; -- output copy to hold a pipeline register if needed

   with q3_c18  select 
      absq3D_c18 <= 
         "000" & D_c18						 when "001" | "111", -- mult by 1
         "00" & D_c18 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q3_c18(2)  select 
   w2_c18<= betaw3_c18 - absq3D_c18 when '0',
         betaw3_c18 + absq3D_c18 when others;

   betaw2_c18 <= w2_c18(53 downto 0) & "00"; -- multiplication by the radix
   sel2_c18 <= betaw2_c18(55 downto 50) & D_c18(51 downto 49);
   SelFunctionTable2: selFunction_Freq300_uid4
      port map ( X => sel2_c18,
                 Y => q2_copy31_c18);
   q2_c18 <= q2_copy31_c18; -- output copy to hold a pipeline register if needed

   with q2_c18  select 
      absq2D_c18 <= 
         "000" & D_c18						 when "001" | "111", -- mult by 1
         "00" & D_c18 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q2_c19(2)  select 
   w1_c19<= betaw2_c19 - absq2D_c19 when '0',
         betaw2_c19 + absq2D_c19 when others;

   betaw1_c19 <= w1_c19(53 downto 0) & "00"; -- multiplication by the radix
   sel1_c19 <= betaw1_c19(55 downto 50) & D_c19(51 downto 49);
   SelFunctionTable1: selFunction_Freq300_uid4
      port map ( X => sel1_c19,
                 Y => q1_copy32_c19);
   q1_c19 <= q1_copy32_c19; -- output copy to hold a pipeline register if needed

   with q1_c19  select 
      absq1D_c19 <= 
         "000" & D_c19						 when "001" | "111", -- mult by 1
         "00" & D_c19 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q1_c19(2)  select 
   w0_c19<= betaw1_c19 - absq1D_c19 when '0',
         betaw1_c19 + absq1D_c19 when others;

   wfinal_c19 <= w0_c19(53 downto 0);
   qM0_c19 <= wfinal_c19(53); -- rounding bit is the sign of the remainder
   qP28_c0 <=      q28_c0(1 downto 0);
   qM28_c0 <=      q28_c0(2) & "0";
   qP27_c0 <=      q27_c0(1 downto 0);
   qM27_c0 <=      q27_c0(2) & "0";
   qP26_c1 <=      q26_c1(1 downto 0);
   qM26_c1 <=      q26_c1(2) & "0";
   qP25_c2 <=      q25_c2(1 downto 0);
   qM25_c2 <=      q25_c2(2) & "0";
   qP24_c3 <=      q24_c3(1 downto 0);
   qM24_c3 <=      q24_c3(2) & "0";
   qP23_c3 <=      q23_c3(1 downto 0);
   qM23_c3 <=      q23_c3(2) & "0";
   qP22_c4 <=      q22_c4(1 downto 0);
   qM22_c4 <=      q22_c4(2) & "0";
   qP21_c5 <=      q21_c5(1 downto 0);
   qM21_c5 <=      q21_c5(2) & "0";
   qP20_c5 <=      q20_c5(1 downto 0);
   qM20_c5 <=      q20_c5(2) & "0";
   qP19_c6 <=      q19_c6(1 downto 0);
   qM19_c6 <=      q19_c6(2) & "0";
   qP18_c7 <=      q18_c7(1 downto 0);
   qM18_c7 <=      q18_c7(2) & "0";
   qP17_c8 <=      q17_c8(1 downto 0);
   qM17_c8 <=      q17_c8(2) & "0";
   qP16_c8 <=      q16_c8(1 downto 0);
   qM16_c8 <=      q16_c8(2) & "0";
   qP15_c9 <=      q15_c9(1 downto 0);
   qM15_c9 <=      q15_c9(2) & "0";
   qP14_c10 <=      q14_c10(1 downto 0);
   qM14_c10 <=      q14_c10(2) & "0";
   qP13_c10 <=      q13_c10(1 downto 0);
   qM13_c10 <=      q13_c10(2) & "0";
   qP12_c11 <=      q12_c11(1 downto 0);
   qM12_c11 <=      q12_c11(2) & "0";
   qP11_c12 <=      q11_c12(1 downto 0);
   qM11_c12 <=      q11_c12(2) & "0";
   qP10_c13 <=      q10_c13(1 downto 0);
   qM10_c13 <=      q10_c13(2) & "0";
   qP9_c13 <=      q9_c13(1 downto 0);
   qM9_c13 <=      q9_c13(2) & "0";
   qP8_c14 <=      q8_c14(1 downto 0);
   qM8_c14 <=      q8_c14(2) & "0";
   qP7_c15 <=      q7_c15(1 downto 0);
   qM7_c15 <=      q7_c15(2) & "0";
   qP6_c15 <=      q6_c15(1 downto 0);
   qM6_c15 <=      q6_c15(2) & "0";
   qP5_c16 <=      q5_c16(1 downto 0);
   qM5_c16 <=      q5_c16(2) & "0";
   qP4_c17 <=      q4_c17(1 downto 0);
   qM4_c17 <=      q4_c17(2) & "0";
   qP3_c18 <=      q3_c18(1 downto 0);
   qM3_c18 <=      q3_c18(2) & "0";
   qP2_c18 <=      q2_c18(1 downto 0);
   qM2_c18 <=      q2_c18(2) & "0";
   qP1_c19 <=      q1_c19(1 downto 0);
   qM1_c19 <=      q1_c19(2) & "0";
   qP_c19 <= qP28_c19 & qP27_c19 & qP26_c19 & qP25_c19 & qP24_c19 & qP23_c19 & qP22_c19 & qP21_c19 & qP20_c19 & qP19_c19 & qP18_c19 & qP17_c19 & qP16_c19 & qP15_c19 & qP14_c19 & qP13_c19 & qP12_c19 & qP11_c19 & qP10_c19 & qP9_c19 & qP8_c19 & qP7_c19 & qP6_c19 & qP5_c19 & qP4_c19 & qP3_c19 & qP2_c19 & qP1_c19;
   qM_c19 <= qM28_c19(0) & qM27_c19 & qM26_c19 & qM25_c19 & qM24_c19 & qM23_c19 & qM22_c19 & qM21_c19 & qM20_c19 & qM19_c19 & qM18_c19 & qM17_c19 & qM16_c19 & qM15_c19 & qM14_c19 & qM13_c19 & qM12_c19 & qM11_c19 & qM10_c19 & qM9_c19 & qM8_c19 & qM7_c19 & qM6_c19 & qM5_c19 & qM4_c19 & qM3_c19 & qM2_c19 & qM1_c19 & qM0_c19;
   quotient_c20 <= qP_c20 - qM_c20;
   -- We need a mR in (0, -wf-2) format: 1+wF fraction bits, 1 round bit, and 1 guard bit for the normalisation,
   -- quotient is the truncation of the exact quotient to at least 2^(-wF-2) bits
   -- now discarding its possible known MSB zeroes, and dropping the possible extra LSB bit (due to radix 4) 
   mR_c20 <= quotient_c20(54 downto 0); 
   -- normalisation
   fRnorm_c20 <=    mR_c20(53 downto 1)  when mR_c20(54)= '1'
           else mR_c20(52 downto 0);  -- now fRnorm is a (-1, -wF-1) fraction
   round_c20 <= fRnorm_c20(0); 
   expR1_c20 <= expR0_c20 + ("000" & (9 downto 1 => '1') & mR_c20(54)); -- add back bias
   -- final rounding
   expfrac_c20 <= expR1_c20 & fRnorm_c20(52 downto 1) ;
   expfracR_c20 <= expfrac_c20 + ((64 downto 1 => '0') & round_c20);
   exnR_c20 <=      "00"  when expfracR_c20(64) = '1'   -- underflow
           else "10"  when  expfracR_c20(64 downto 63) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_c20  select 
      exnRfinal_c20 <= 
         exnR_c20   when "01", -- normal
         exnR0_c20  when others;
   R <= exnRfinal_c20 & sR_c20 & expfracR_c20(62 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          selFunction_Freq100_uid4
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity selFunction_Freq100_uid4 is
    port (X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of selFunction_Freq100_uid4 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000000000",
      "000" when "000000001",
      "000" when "000000010",
      "000" when "000000011",
      "000" when "000000100",
      "000" when "000000101",
      "000" when "000000110",
      "000" when "000000111",
      "000" when "000001000",
      "000" when "000001001",
      "000" when "000001010",
      "000" when "000001011",
      "000" when "000001100",
      "000" when "000001101",
      "000" when "000001110",
      "000" when "000001111",
      "001" when "000010000",
      "000" when "000010001",
      "000" when "000010010",
      "000" when "000010011",
      "000" when "000010100",
      "000" when "000010101",
      "000" when "000010110",
      "000" when "000010111",
      "001" when "000011000",
      "001" when "000011001",
      "001" when "000011010",
      "001" when "000011011",
      "000" when "000011100",
      "000" when "000011101",
      "000" when "000011110",
      "000" when "000011111",
      "001" when "000100000",
      "001" when "000100001",
      "001" when "000100010",
      "001" when "000100011",
      "001" when "000100100",
      "001" when "000100101",
      "001" when "000100110",
      "000" when "000100111",
      "001" when "000101000",
      "001" when "000101001",
      "001" when "000101010",
      "001" when "000101011",
      "001" when "000101100",
      "001" when "000101101",
      "001" when "000101110",
      "001" when "000101111",
      "010" when "000110000",
      "001" when "000110001",
      "001" when "000110010",
      "001" when "000110011",
      "001" when "000110100",
      "001" when "000110101",
      "001" when "000110110",
      "001" when "000110111",
      "010" when "000111000",
      "010" when "000111001",
      "001" when "000111010",
      "001" when "000111011",
      "001" when "000111100",
      "001" when "000111101",
      "001" when "000111110",
      "001" when "000111111",
      "010" when "001000000",
      "010" when "001000001",
      "010" when "001000010",
      "001" when "001000011",
      "001" when "001000100",
      "001" when "001000101",
      "001" when "001000110",
      "001" when "001000111",
      "010" when "001001000",
      "010" when "001001001",
      "010" when "001001010",
      "010" when "001001011",
      "001" when "001001100",
      "001" when "001001101",
      "001" when "001001110",
      "001" when "001001111",
      "010" when "001010000",
      "010" when "001010001",
      "010" when "001010010",
      "010" when "001010011",
      "010" when "001010100",
      "010" when "001010101",
      "001" when "001010110",
      "001" when "001010111",
      "010" when "001011000",
      "010" when "001011001",
      "010" when "001011010",
      "010" when "001011011",
      "010" when "001011100",
      "010" when "001011101",
      "010" when "001011110",
      "001" when "001011111",
      "010" when "001100000",
      "010" when "001100001",
      "010" when "001100010",
      "010" when "001100011",
      "010" when "001100100",
      "010" when "001100101",
      "010" when "001100110",
      "010" when "001100111",
      "010" when "001101000",
      "010" when "001101001",
      "010" when "001101010",
      "010" when "001101011",
      "010" when "001101100",
      "010" when "001101101",
      "010" when "001101110",
      "010" when "001101111",
      "010" when "001110000",
      "010" when "001110001",
      "010" when "001110010",
      "010" when "001110011",
      "010" when "001110100",
      "010" when "001110101",
      "010" when "001110110",
      "010" when "001110111",
      "010" when "001111000",
      "010" when "001111001",
      "010" when "001111010",
      "010" when "001111011",
      "010" when "001111100",
      "010" when "001111101",
      "010" when "001111110",
      "010" when "001111111",
      "010" when "010000000",
      "010" when "010000001",
      "010" when "010000010",
      "010" when "010000011",
      "010" when "010000100",
      "010" when "010000101",
      "010" when "010000110",
      "010" when "010000111",
      "010" when "010001000",
      "010" when "010001001",
      "010" when "010001010",
      "010" when "010001011",
      "010" when "010001100",
      "010" when "010001101",
      "010" when "010001110",
      "010" when "010001111",
      "010" when "010010000",
      "010" when "010010001",
      "010" when "010010010",
      "010" when "010010011",
      "010" when "010010100",
      "010" when "010010101",
      "010" when "010010110",
      "010" when "010010111",
      "010" when "010011000",
      "010" when "010011001",
      "010" when "010011010",
      "010" when "010011011",
      "010" when "010011100",
      "010" when "010011101",
      "010" when "010011110",
      "010" when "010011111",
      "010" when "010100000",
      "010" when "010100001",
      "010" when "010100010",
      "010" when "010100011",
      "010" when "010100100",
      "010" when "010100101",
      "010" when "010100110",
      "010" when "010100111",
      "010" when "010101000",
      "010" when "010101001",
      "010" when "010101010",
      "010" when "010101011",
      "010" when "010101100",
      "010" when "010101101",
      "010" when "010101110",
      "010" when "010101111",
      "010" when "010110000",
      "010" when "010110001",
      "010" when "010110010",
      "010" when "010110011",
      "010" when "010110100",
      "010" when "010110101",
      "010" when "010110110",
      "010" when "010110111",
      "010" when "010111000",
      "010" when "010111001",
      "010" when "010111010",
      "010" when "010111011",
      "010" when "010111100",
      "010" when "010111101",
      "010" when "010111110",
      "010" when "010111111",
      "010" when "011000000",
      "010" when "011000001",
      "010" when "011000010",
      "010" when "011000011",
      "010" when "011000100",
      "010" when "011000101",
      "010" when "011000110",
      "010" when "011000111",
      "010" when "011001000",
      "010" when "011001001",
      "010" when "011001010",
      "010" when "011001011",
      "010" when "011001100",
      "010" when "011001101",
      "010" when "011001110",
      "010" when "011001111",
      "010" when "011010000",
      "010" when "011010001",
      "010" when "011010010",
      "010" when "011010011",
      "010" when "011010100",
      "010" when "011010101",
      "010" when "011010110",
      "010" when "011010111",
      "010" when "011011000",
      "010" when "011011001",
      "010" when "011011010",
      "010" when "011011011",
      "010" when "011011100",
      "010" when "011011101",
      "010" when "011011110",
      "010" when "011011111",
      "010" when "011100000",
      "010" when "011100001",
      "010" when "011100010",
      "010" when "011100011",
      "010" when "011100100",
      "010" when "011100101",
      "010" when "011100110",
      "010" when "011100111",
      "010" when "011101000",
      "010" when "011101001",
      "010" when "011101010",
      "010" when "011101011",
      "010" when "011101100",
      "010" when "011101101",
      "010" when "011101110",
      "010" when "011101111",
      "010" when "011110000",
      "010" when "011110001",
      "010" when "011110010",
      "010" when "011110011",
      "010" when "011110100",
      "010" when "011110101",
      "010" when "011110110",
      "010" when "011110111",
      "010" when "011111000",
      "010" when "011111001",
      "010" when "011111010",
      "010" when "011111011",
      "010" when "011111100",
      "010" when "011111101",
      "010" when "011111110",
      "010" when "011111111",
      "110" when "100000000",
      "110" when "100000001",
      "110" when "100000010",
      "110" when "100000011",
      "110" when "100000100",
      "110" when "100000101",
      "110" when "100000110",
      "110" when "100000111",
      "110" when "100001000",
      "110" when "100001001",
      "110" when "100001010",
      "110" when "100001011",
      "110" when "100001100",
      "110" when "100001101",
      "110" when "100001110",
      "110" when "100001111",
      "110" when "100010000",
      "110" when "100010001",
      "110" when "100010010",
      "110" when "100010011",
      "110" when "100010100",
      "110" when "100010101",
      "110" when "100010110",
      "110" when "100010111",
      "110" when "100011000",
      "110" when "100011001",
      "110" when "100011010",
      "110" when "100011011",
      "110" when "100011100",
      "110" when "100011101",
      "110" when "100011110",
      "110" when "100011111",
      "110" when "100100000",
      "110" when "100100001",
      "110" when "100100010",
      "110" when "100100011",
      "110" when "100100100",
      "110" when "100100101",
      "110" when "100100110",
      "110" when "100100111",
      "110" when "100101000",
      "110" when "100101001",
      "110" when "100101010",
      "110" when "100101011",
      "110" when "100101100",
      "110" when "100101101",
      "110" when "100101110",
      "110" when "100101111",
      "110" when "100110000",
      "110" when "100110001",
      "110" when "100110010",
      "110" when "100110011",
      "110" when "100110100",
      "110" when "100110101",
      "110" when "100110110",
      "110" when "100110111",
      "110" when "100111000",
      "110" when "100111001",
      "110" when "100111010",
      "110" when "100111011",
      "110" when "100111100",
      "110" when "100111101",
      "110" when "100111110",
      "110" when "100111111",
      "110" when "101000000",
      "110" when "101000001",
      "110" when "101000010",
      "110" when "101000011",
      "110" when "101000100",
      "110" when "101000101",
      "110" when "101000110",
      "110" when "101000111",
      "110" when "101001000",
      "110" when "101001001",
      "110" when "101001010",
      "110" when "101001011",
      "110" when "101001100",
      "110" when "101001101",
      "110" when "101001110",
      "110" when "101001111",
      "110" when "101010000",
      "110" when "101010001",
      "110" when "101010010",
      "110" when "101010011",
      "110" when "101010100",
      "110" when "101010101",
      "110" when "101010110",
      "110" when "101010111",
      "110" when "101011000",
      "110" when "101011001",
      "110" when "101011010",
      "110" when "101011011",
      "110" when "101011100",
      "110" when "101011101",
      "110" when "101011110",
      "110" when "101011111",
      "110" when "101100000",
      "110" when "101100001",
      "110" when "101100010",
      "110" when "101100011",
      "110" when "101100100",
      "110" when "101100101",
      "110" when "101100110",
      "110" when "101100111",
      "110" when "101101000",
      "110" when "101101001",
      "110" when "101101010",
      "110" when "101101011",
      "110" when "101101100",
      "110" when "101101101",
      "110" when "101101110",
      "110" when "101101111",
      "110" when "101110000",
      "110" when "101110001",
      "110" when "101110010",
      "110" when "101110011",
      "110" when "101110100",
      "110" when "101110101",
      "110" when "101110110",
      "110" when "101110111",
      "110" when "101111000",
      "110" when "101111001",
      "110" when "101111010",
      "110" when "101111011",
      "110" when "101111100",
      "110" when "101111101",
      "110" when "101111110",
      "110" when "101111111",
      "110" when "110000000",
      "110" when "110000001",
      "110" when "110000010",
      "110" when "110000011",
      "110" when "110000100",
      "110" when "110000101",
      "110" when "110000110",
      "110" when "110000111",
      "110" when "110001000",
      "110" when "110001001",
      "110" when "110001010",
      "110" when "110001011",
      "110" when "110001100",
      "110" when "110001101",
      "110" when "110001110",
      "110" when "110001111",
      "110" when "110010000",
      "110" when "110010001",
      "110" when "110010010",
      "110" when "110010011",
      "110" when "110010100",
      "110" when "110010101",
      "110" when "110010110",
      "110" when "110010111",
      "110" when "110011000",
      "110" when "110011001",
      "110" when "110011010",
      "110" when "110011011",
      "110" when "110011100",
      "110" when "110011101",
      "110" when "110011110",
      "110" when "110011111",
      "110" when "110100000",
      "110" when "110100001",
      "110" when "110100010",
      "110" when "110100011",
      "110" when "110100100",
      "110" when "110100101",
      "110" when "110100110",
      "110" when "110100111",
      "110" when "110101000",
      "110" when "110101001",
      "110" when "110101010",
      "110" when "110101011",
      "110" when "110101100",
      "110" when "110101101",
      "110" when "110101110",
      "111" when "110101111",
      "110" when "110110000",
      "110" when "110110001",
      "110" when "110110010",
      "110" when "110110011",
      "110" when "110110100",
      "111" when "110110101",
      "111" when "110110110",
      "111" when "110110111",
      "110" when "110111000",
      "110" when "110111001",
      "110" when "110111010",
      "110" when "110111011",
      "111" when "110111100",
      "111" when "110111101",
      "111" when "110111110",
      "111" when "110111111",
      "110" when "111000000",
      "110" when "111000001",
      "111" when "111000010",
      "111" when "111000011",
      "111" when "111000100",
      "111" when "111000101",
      "111" when "111000110",
      "111" when "111000111",
      "110" when "111001000",
      "111" when "111001001",
      "111" when "111001010",
      "111" when "111001011",
      "111" when "111001100",
      "111" when "111001101",
      "111" when "111001110",
      "111" when "111001111",
      "111" when "111010000",
      "111" when "111010001",
      "111" when "111010010",
      "111" when "111010011",
      "111" when "111010100",
      "111" when "111010101",
      "111" when "111010110",
      "111" when "111010111",
      "111" when "111011000",
      "111" when "111011001",
      "111" when "111011010",
      "111" when "111011011",
      "111" when "111011100",
      "111" when "111011101",
      "111" when "111011110",
      "111" when "111011111",
      "111" when "111100000",
      "111" when "111100001",
      "111" when "111100010",
      "111" when "111100011",
      "111" when "111100100",
      "111" when "111100101",
      "111" when "111100110",
      "111" when "111100111",
      "111" when "111101000",
      "111" when "111101001",
      "111" when "111101010",
      "111" when "111101011",
      "000" when "111101100",
      "000" when "111101101",
      "000" when "111101110",
      "000" when "111101111",
      "000" when "111110000",
      "000" when "111110001",
      "000" when "111110010",
      "000" when "111110011",
      "000" when "111110100",
      "000" when "111110101",
      "000" when "111110110",
      "000" when "111110111",
      "000" when "111111000",
      "000" when "111111001",
      "000" when "111111010",
      "000" when "111111011",
      "000" when "111111100",
      "000" when "111111101",
      "000" when "111111110",
      "000" when "111111111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            FloatingPointDivider
--                         (FPDiv_11_52_Freq100_uid2)
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 6 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointDivider_64_16_008000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6 : in std_logic;
          X : in  std_logic_vector(11+52+2 downto 0);
          Y : in  std_logic_vector(11+52+2 downto 0);
          R : out  std_logic_vector(11+52+2 downto 0)   );
end entity;

architecture arch of FloatingPointDivider_64_16_008000 is
   component selFunction_Freq100_uid4 is
      port ( X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal fX_c0 :  std_logic_vector(52 downto 0);
signal fY_c0 :  std_logic_vector(52 downto 0);
signal expR0_c0, expR0_c1, expR0_c2, expR0_c3, expR0_c4, expR0_c5, expR0_c6 :  std_logic_vector(12 downto 0);
signal sR_c0, sR_c1, sR_c2, sR_c3, sR_c4, sR_c5, sR_c6 :  std_logic;
signal exnXY_c0 :  std_logic_vector(3 downto 0);
signal exnR0_c0, exnR0_c1, exnR0_c2, exnR0_c3, exnR0_c4, exnR0_c5, exnR0_c6 :  std_logic_vector(1 downto 0);
signal D_c0, D_c1, D_c2, D_c3, D_c4, D_c5, D_c6 :  std_logic_vector(52 downto 0);
signal psX_c0 :  std_logic_vector(53 downto 0);
signal betaw28_c0 :  std_logic_vector(55 downto 0);
signal sel28_c0 :  std_logic_vector(8 downto 0);
signal q28_c0 :  std_logic_vector(2 downto 0);
signal q28_copy5_c0 :  std_logic_vector(2 downto 0);
signal absq28D_c0 :  std_logic_vector(55 downto 0);
signal w27_c0 :  std_logic_vector(55 downto 0);
signal betaw27_c0 :  std_logic_vector(55 downto 0);
signal sel27_c0 :  std_logic_vector(8 downto 0);
signal q27_c0 :  std_logic_vector(2 downto 0);
signal q27_copy6_c0 :  std_logic_vector(2 downto 0);
signal absq27D_c0 :  std_logic_vector(55 downto 0);
signal w26_c0 :  std_logic_vector(55 downto 0);
signal betaw26_c0 :  std_logic_vector(55 downto 0);
signal sel26_c0 :  std_logic_vector(8 downto 0);
signal q26_c0 :  std_logic_vector(2 downto 0);
signal q26_copy7_c0 :  std_logic_vector(2 downto 0);
signal absq26D_c0 :  std_logic_vector(55 downto 0);
signal w25_c0 :  std_logic_vector(55 downto 0);
signal betaw25_c0 :  std_logic_vector(55 downto 0);
signal sel25_c0 :  std_logic_vector(8 downto 0);
signal q25_c0 :  std_logic_vector(2 downto 0);
signal q25_copy8_c0 :  std_logic_vector(2 downto 0);
signal absq25D_c0 :  std_logic_vector(55 downto 0);
signal w24_c0 :  std_logic_vector(55 downto 0);
signal betaw24_c0, betaw24_c1 :  std_logic_vector(55 downto 0);
signal sel24_c0 :  std_logic_vector(8 downto 0);
signal q24_c0, q24_c1 :  std_logic_vector(2 downto 0);
signal q24_copy9_c0 :  std_logic_vector(2 downto 0);
signal absq24D_c0, absq24D_c1 :  std_logic_vector(55 downto 0);
signal w23_c1 :  std_logic_vector(55 downto 0);
signal betaw23_c1 :  std_logic_vector(55 downto 0);
signal sel23_c1 :  std_logic_vector(8 downto 0);
signal q23_c1 :  std_logic_vector(2 downto 0);
signal q23_copy10_c1 :  std_logic_vector(2 downto 0);
signal absq23D_c1 :  std_logic_vector(55 downto 0);
signal w22_c1 :  std_logic_vector(55 downto 0);
signal betaw22_c1 :  std_logic_vector(55 downto 0);
signal sel22_c1 :  std_logic_vector(8 downto 0);
signal q22_c1 :  std_logic_vector(2 downto 0);
signal q22_copy11_c1 :  std_logic_vector(2 downto 0);
signal absq22D_c1 :  std_logic_vector(55 downto 0);
signal w21_c1 :  std_logic_vector(55 downto 0);
signal betaw21_c1 :  std_logic_vector(55 downto 0);
signal sel21_c1 :  std_logic_vector(8 downto 0);
signal q21_c1 :  std_logic_vector(2 downto 0);
signal q21_copy12_c1 :  std_logic_vector(2 downto 0);
signal absq21D_c1 :  std_logic_vector(55 downto 0);
signal w20_c1 :  std_logic_vector(55 downto 0);
signal betaw20_c1, betaw20_c2 :  std_logic_vector(55 downto 0);
signal sel20_c1 :  std_logic_vector(8 downto 0);
signal q20_c1, q20_c2 :  std_logic_vector(2 downto 0);
signal q20_copy13_c1 :  std_logic_vector(2 downto 0);
signal absq20D_c1, absq20D_c2 :  std_logic_vector(55 downto 0);
signal w19_c2 :  std_logic_vector(55 downto 0);
signal betaw19_c2 :  std_logic_vector(55 downto 0);
signal sel19_c2 :  std_logic_vector(8 downto 0);
signal q19_c2 :  std_logic_vector(2 downto 0);
signal q19_copy14_c2 :  std_logic_vector(2 downto 0);
signal absq19D_c2 :  std_logic_vector(55 downto 0);
signal w18_c2 :  std_logic_vector(55 downto 0);
signal betaw18_c2 :  std_logic_vector(55 downto 0);
signal sel18_c2 :  std_logic_vector(8 downto 0);
signal q18_c2 :  std_logic_vector(2 downto 0);
signal q18_copy15_c2 :  std_logic_vector(2 downto 0);
signal absq18D_c2 :  std_logic_vector(55 downto 0);
signal w17_c2 :  std_logic_vector(55 downto 0);
signal betaw17_c2 :  std_logic_vector(55 downto 0);
signal sel17_c2 :  std_logic_vector(8 downto 0);
signal q17_c2 :  std_logic_vector(2 downto 0);
signal q17_copy16_c2 :  std_logic_vector(2 downto 0);
signal absq17D_c2 :  std_logic_vector(55 downto 0);
signal w16_c2 :  std_logic_vector(55 downto 0);
signal betaw16_c2 :  std_logic_vector(55 downto 0);
signal sel16_c2 :  std_logic_vector(8 downto 0);
signal q16_c2 :  std_logic_vector(2 downto 0);
signal q16_copy17_c2 :  std_logic_vector(2 downto 0);
signal absq16D_c2 :  std_logic_vector(55 downto 0);
signal w15_c2 :  std_logic_vector(55 downto 0);
signal betaw15_c2, betaw15_c3 :  std_logic_vector(55 downto 0);
signal sel15_c2 :  std_logic_vector(8 downto 0);
signal q15_c3 :  std_logic_vector(2 downto 0);
signal q15_copy18_c2, q15_copy18_c3 :  std_logic_vector(2 downto 0);
signal absq15D_c3 :  std_logic_vector(55 downto 0);
signal w14_c3 :  std_logic_vector(55 downto 0);
signal betaw14_c3 :  std_logic_vector(55 downto 0);
signal sel14_c3 :  std_logic_vector(8 downto 0);
signal q14_c3 :  std_logic_vector(2 downto 0);
signal q14_copy19_c3 :  std_logic_vector(2 downto 0);
signal absq14D_c3 :  std_logic_vector(55 downto 0);
signal w13_c3 :  std_logic_vector(55 downto 0);
signal betaw13_c3 :  std_logic_vector(55 downto 0);
signal sel13_c3 :  std_logic_vector(8 downto 0);
signal q13_c3 :  std_logic_vector(2 downto 0);
signal q13_copy20_c3 :  std_logic_vector(2 downto 0);
signal absq13D_c3 :  std_logic_vector(55 downto 0);
signal w12_c3 :  std_logic_vector(55 downto 0);
signal betaw12_c3 :  std_logic_vector(55 downto 0);
signal sel12_c3 :  std_logic_vector(8 downto 0);
signal q12_c3 :  std_logic_vector(2 downto 0);
signal q12_copy21_c3 :  std_logic_vector(2 downto 0);
signal absq12D_c3 :  std_logic_vector(55 downto 0);
signal w11_c3 :  std_logic_vector(55 downto 0);
signal betaw11_c3, betaw11_c4 :  std_logic_vector(55 downto 0);
signal sel11_c3 :  std_logic_vector(8 downto 0);
signal q11_c3, q11_c4 :  std_logic_vector(2 downto 0);
signal q11_copy22_c3 :  std_logic_vector(2 downto 0);
signal absq11D_c3, absq11D_c4 :  std_logic_vector(55 downto 0);
signal w10_c4 :  std_logic_vector(55 downto 0);
signal betaw10_c4 :  std_logic_vector(55 downto 0);
signal sel10_c4 :  std_logic_vector(8 downto 0);
signal q10_c4 :  std_logic_vector(2 downto 0);
signal q10_copy23_c4 :  std_logic_vector(2 downto 0);
signal absq10D_c4 :  std_logic_vector(55 downto 0);
signal w9_c4 :  std_logic_vector(55 downto 0);
signal betaw9_c4 :  std_logic_vector(55 downto 0);
signal sel9_c4 :  std_logic_vector(8 downto 0);
signal q9_c4 :  std_logic_vector(2 downto 0);
signal q9_copy24_c4 :  std_logic_vector(2 downto 0);
signal absq9D_c4 :  std_logic_vector(55 downto 0);
signal w8_c4 :  std_logic_vector(55 downto 0);
signal betaw8_c4 :  std_logic_vector(55 downto 0);
signal sel8_c4 :  std_logic_vector(8 downto 0);
signal q8_c4 :  std_logic_vector(2 downto 0);
signal q8_copy25_c4 :  std_logic_vector(2 downto 0);
signal absq8D_c4 :  std_logic_vector(55 downto 0);
signal w7_c4 :  std_logic_vector(55 downto 0);
signal betaw7_c4 :  std_logic_vector(55 downto 0);
signal sel7_c4 :  std_logic_vector(8 downto 0);
signal q7_c4 :  std_logic_vector(2 downto 0);
signal q7_copy26_c4 :  std_logic_vector(2 downto 0);
signal absq7D_c4 :  std_logic_vector(55 downto 0);
signal w6_c4 :  std_logic_vector(55 downto 0);
signal betaw6_c4, betaw6_c5 :  std_logic_vector(55 downto 0);
signal sel6_c4 :  std_logic_vector(8 downto 0);
signal q6_c5 :  std_logic_vector(2 downto 0);
signal q6_copy27_c4, q6_copy27_c5 :  std_logic_vector(2 downto 0);
signal absq6D_c5 :  std_logic_vector(55 downto 0);
signal w5_c5 :  std_logic_vector(55 downto 0);
signal betaw5_c5 :  std_logic_vector(55 downto 0);
signal sel5_c5 :  std_logic_vector(8 downto 0);
signal q5_c5 :  std_logic_vector(2 downto 0);
signal q5_copy28_c5 :  std_logic_vector(2 downto 0);
signal absq5D_c5 :  std_logic_vector(55 downto 0);
signal w4_c5 :  std_logic_vector(55 downto 0);
signal betaw4_c5 :  std_logic_vector(55 downto 0);
signal sel4_c5 :  std_logic_vector(8 downto 0);
signal q4_c5 :  std_logic_vector(2 downto 0);
signal q4_copy29_c5 :  std_logic_vector(2 downto 0);
signal absq4D_c5 :  std_logic_vector(55 downto 0);
signal w3_c5 :  std_logic_vector(55 downto 0);
signal betaw3_c5 :  std_logic_vector(55 downto 0);
signal sel3_c5 :  std_logic_vector(8 downto 0);
signal q3_c5 :  std_logic_vector(2 downto 0);
signal q3_copy30_c5 :  std_logic_vector(2 downto 0);
signal absq3D_c5 :  std_logic_vector(55 downto 0);
signal w2_c5 :  std_logic_vector(55 downto 0);
signal betaw2_c5, betaw2_c6 :  std_logic_vector(55 downto 0);
signal sel2_c5 :  std_logic_vector(8 downto 0);
signal q2_c5, q2_c6 :  std_logic_vector(2 downto 0);
signal q2_copy31_c5 :  std_logic_vector(2 downto 0);
signal absq2D_c5, absq2D_c6 :  std_logic_vector(55 downto 0);
signal w1_c6 :  std_logic_vector(55 downto 0);
signal betaw1_c6 :  std_logic_vector(55 downto 0);
signal sel1_c6 :  std_logic_vector(8 downto 0);
signal q1_c6 :  std_logic_vector(2 downto 0);
signal q1_copy32_c6 :  std_logic_vector(2 downto 0);
signal absq1D_c6 :  std_logic_vector(55 downto 0);
signal w0_c6 :  std_logic_vector(55 downto 0);
signal wfinal_c6 :  std_logic_vector(53 downto 0);
signal qM0_c6 :  std_logic;
signal qP28_c0, qP28_c1, qP28_c2, qP28_c3, qP28_c4, qP28_c5, qP28_c6 :  std_logic_vector(1 downto 0);
signal qM28_c0, qM28_c1, qM28_c2, qM28_c3, qM28_c4, qM28_c5, qM28_c6 :  std_logic_vector(1 downto 0);
signal qP27_c0, qP27_c1, qP27_c2, qP27_c3, qP27_c4, qP27_c5, qP27_c6 :  std_logic_vector(1 downto 0);
signal qM27_c0, qM27_c1, qM27_c2, qM27_c3, qM27_c4, qM27_c5, qM27_c6 :  std_logic_vector(1 downto 0);
signal qP26_c0, qP26_c1, qP26_c2, qP26_c3, qP26_c4, qP26_c5, qP26_c6 :  std_logic_vector(1 downto 0);
signal qM26_c0, qM26_c1, qM26_c2, qM26_c3, qM26_c4, qM26_c5, qM26_c6 :  std_logic_vector(1 downto 0);
signal qP25_c0, qP25_c1, qP25_c2, qP25_c3, qP25_c4, qP25_c5, qP25_c6 :  std_logic_vector(1 downto 0);
signal qM25_c0, qM25_c1, qM25_c2, qM25_c3, qM25_c4, qM25_c5, qM25_c6 :  std_logic_vector(1 downto 0);
signal qP24_c0, qP24_c1, qP24_c2, qP24_c3, qP24_c4, qP24_c5, qP24_c6 :  std_logic_vector(1 downto 0);
signal qM24_c0, qM24_c1, qM24_c2, qM24_c3, qM24_c4, qM24_c5, qM24_c6 :  std_logic_vector(1 downto 0);
signal qP23_c1, qP23_c2, qP23_c3, qP23_c4, qP23_c5, qP23_c6 :  std_logic_vector(1 downto 0);
signal qM23_c1, qM23_c2, qM23_c3, qM23_c4, qM23_c5, qM23_c6 :  std_logic_vector(1 downto 0);
signal qP22_c1, qP22_c2, qP22_c3, qP22_c4, qP22_c5, qP22_c6 :  std_logic_vector(1 downto 0);
signal qM22_c1, qM22_c2, qM22_c3, qM22_c4, qM22_c5, qM22_c6 :  std_logic_vector(1 downto 0);
signal qP21_c1, qP21_c2, qP21_c3, qP21_c4, qP21_c5, qP21_c6 :  std_logic_vector(1 downto 0);
signal qM21_c1, qM21_c2, qM21_c3, qM21_c4, qM21_c5, qM21_c6 :  std_logic_vector(1 downto 0);
signal qP20_c1, qP20_c2, qP20_c3, qP20_c4, qP20_c5, qP20_c6 :  std_logic_vector(1 downto 0);
signal qM20_c1, qM20_c2, qM20_c3, qM20_c4, qM20_c5, qM20_c6 :  std_logic_vector(1 downto 0);
signal qP19_c2, qP19_c3, qP19_c4, qP19_c5, qP19_c6 :  std_logic_vector(1 downto 0);
signal qM19_c2, qM19_c3, qM19_c4, qM19_c5, qM19_c6 :  std_logic_vector(1 downto 0);
signal qP18_c2, qP18_c3, qP18_c4, qP18_c5, qP18_c6 :  std_logic_vector(1 downto 0);
signal qM18_c2, qM18_c3, qM18_c4, qM18_c5, qM18_c6 :  std_logic_vector(1 downto 0);
signal qP17_c2, qP17_c3, qP17_c4, qP17_c5, qP17_c6 :  std_logic_vector(1 downto 0);
signal qM17_c2, qM17_c3, qM17_c4, qM17_c5, qM17_c6 :  std_logic_vector(1 downto 0);
signal qP16_c2, qP16_c3, qP16_c4, qP16_c5, qP16_c6 :  std_logic_vector(1 downto 0);
signal qM16_c2, qM16_c3, qM16_c4, qM16_c5, qM16_c6 :  std_logic_vector(1 downto 0);
signal qP15_c3, qP15_c4, qP15_c5, qP15_c6 :  std_logic_vector(1 downto 0);
signal qM15_c3, qM15_c4, qM15_c5, qM15_c6 :  std_logic_vector(1 downto 0);
signal qP14_c3, qP14_c4, qP14_c5, qP14_c6 :  std_logic_vector(1 downto 0);
signal qM14_c3, qM14_c4, qM14_c5, qM14_c6 :  std_logic_vector(1 downto 0);
signal qP13_c3, qP13_c4, qP13_c5, qP13_c6 :  std_logic_vector(1 downto 0);
signal qM13_c3, qM13_c4, qM13_c5, qM13_c6 :  std_logic_vector(1 downto 0);
signal qP12_c3, qP12_c4, qP12_c5, qP12_c6 :  std_logic_vector(1 downto 0);
signal qM12_c3, qM12_c4, qM12_c5, qM12_c6 :  std_logic_vector(1 downto 0);
signal qP11_c3, qP11_c4, qP11_c5, qP11_c6 :  std_logic_vector(1 downto 0);
signal qM11_c3, qM11_c4, qM11_c5, qM11_c6 :  std_logic_vector(1 downto 0);
signal qP10_c4, qP10_c5, qP10_c6 :  std_logic_vector(1 downto 0);
signal qM10_c4, qM10_c5, qM10_c6 :  std_logic_vector(1 downto 0);
signal qP9_c4, qP9_c5, qP9_c6 :  std_logic_vector(1 downto 0);
signal qM9_c4, qM9_c5, qM9_c6 :  std_logic_vector(1 downto 0);
signal qP8_c4, qP8_c5, qP8_c6 :  std_logic_vector(1 downto 0);
signal qM8_c4, qM8_c5, qM8_c6 :  std_logic_vector(1 downto 0);
signal qP7_c4, qP7_c5, qP7_c6 :  std_logic_vector(1 downto 0);
signal qM7_c4, qM7_c5, qM7_c6 :  std_logic_vector(1 downto 0);
signal qP6_c5, qP6_c6 :  std_logic_vector(1 downto 0);
signal qM6_c5, qM6_c6 :  std_logic_vector(1 downto 0);
signal qP5_c5, qP5_c6 :  std_logic_vector(1 downto 0);
signal qM5_c5, qM5_c6 :  std_logic_vector(1 downto 0);
signal qP4_c5, qP4_c6 :  std_logic_vector(1 downto 0);
signal qM4_c5, qM4_c6 :  std_logic_vector(1 downto 0);
signal qP3_c5, qP3_c6 :  std_logic_vector(1 downto 0);
signal qM3_c5, qM3_c6 :  std_logic_vector(1 downto 0);
signal qP2_c5, qP2_c6 :  std_logic_vector(1 downto 0);
signal qM2_c5, qM2_c6 :  std_logic_vector(1 downto 0);
signal qP1_c6 :  std_logic_vector(1 downto 0);
signal qM1_c6 :  std_logic_vector(1 downto 0);
signal qP_c6 :  std_logic_vector(55 downto 0);
signal qM_c6 :  std_logic_vector(55 downto 0);
signal quotient_c6 :  std_logic_vector(55 downto 0);
signal mR_c6 :  std_logic_vector(54 downto 0);
signal fRnorm_c6 :  std_logic_vector(52 downto 0);
signal round_c6 :  std_logic;
signal expR1_c6 :  std_logic_vector(12 downto 0);
signal expfrac_c6 :  std_logic_vector(64 downto 0);
signal expfracR_c6 :  std_logic_vector(64 downto 0);
signal exnR_c6 :  std_logic_vector(1 downto 0);
signal exnRfinal_c6 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               expR0_c1 <= expR0_c0;
               sR_c1 <= sR_c0;
               exnR0_c1 <= exnR0_c0;
               D_c1 <= D_c0;
               betaw24_c1 <= betaw24_c0;
               q24_c1 <= q24_c0;
               absq24D_c1 <= absq24D_c0;
               qP28_c1 <= qP28_c0;
               qM28_c1 <= qM28_c0;
               qP27_c1 <= qP27_c0;
               qM27_c1 <= qM27_c0;
               qP26_c1 <= qP26_c0;
               qM26_c1 <= qM26_c0;
               qP25_c1 <= qP25_c0;
               qM25_c1 <= qM25_c0;
               qP24_c1 <= qP24_c0;
               qM24_c1 <= qM24_c0;
            end if;
            if ce_2 = '1' then
               expR0_c2 <= expR0_c1;
               sR_c2 <= sR_c1;
               exnR0_c2 <= exnR0_c1;
               D_c2 <= D_c1;
               betaw20_c2 <= betaw20_c1;
               q20_c2 <= q20_c1;
               absq20D_c2 <= absq20D_c1;
               qP28_c2 <= qP28_c1;
               qM28_c2 <= qM28_c1;
               qP27_c2 <= qP27_c1;
               qM27_c2 <= qM27_c1;
               qP26_c2 <= qP26_c1;
               qM26_c2 <= qM26_c1;
               qP25_c2 <= qP25_c1;
               qM25_c2 <= qM25_c1;
               qP24_c2 <= qP24_c1;
               qM24_c2 <= qM24_c1;
               qP23_c2 <= qP23_c1;
               qM23_c2 <= qM23_c1;
               qP22_c2 <= qP22_c1;
               qM22_c2 <= qM22_c1;
               qP21_c2 <= qP21_c1;
               qM21_c2 <= qM21_c1;
               qP20_c2 <= qP20_c1;
               qM20_c2 <= qM20_c1;
            end if;
            if ce_3 = '1' then
               expR0_c3 <= expR0_c2;
               sR_c3 <= sR_c2;
               exnR0_c3 <= exnR0_c2;
               D_c3 <= D_c2;
               betaw15_c3 <= betaw15_c2;
               q15_copy18_c3 <= q15_copy18_c2;
               qP28_c3 <= qP28_c2;
               qM28_c3 <= qM28_c2;
               qP27_c3 <= qP27_c2;
               qM27_c3 <= qM27_c2;
               qP26_c3 <= qP26_c2;
               qM26_c3 <= qM26_c2;
               qP25_c3 <= qP25_c2;
               qM25_c3 <= qM25_c2;
               qP24_c3 <= qP24_c2;
               qM24_c3 <= qM24_c2;
               qP23_c3 <= qP23_c2;
               qM23_c3 <= qM23_c2;
               qP22_c3 <= qP22_c2;
               qM22_c3 <= qM22_c2;
               qP21_c3 <= qP21_c2;
               qM21_c3 <= qM21_c2;
               qP20_c3 <= qP20_c2;
               qM20_c3 <= qM20_c2;
               qP19_c3 <= qP19_c2;
               qM19_c3 <= qM19_c2;
               qP18_c3 <= qP18_c2;
               qM18_c3 <= qM18_c2;
               qP17_c3 <= qP17_c2;
               qM17_c3 <= qM17_c2;
               qP16_c3 <= qP16_c2;
               qM16_c3 <= qM16_c2;
            end if;
            if ce_4 = '1' then
               expR0_c4 <= expR0_c3;
               sR_c4 <= sR_c3;
               exnR0_c4 <= exnR0_c3;
               D_c4 <= D_c3;
               betaw11_c4 <= betaw11_c3;
               q11_c4 <= q11_c3;
               absq11D_c4 <= absq11D_c3;
               qP28_c4 <= qP28_c3;
               qM28_c4 <= qM28_c3;
               qP27_c4 <= qP27_c3;
               qM27_c4 <= qM27_c3;
               qP26_c4 <= qP26_c3;
               qM26_c4 <= qM26_c3;
               qP25_c4 <= qP25_c3;
               qM25_c4 <= qM25_c3;
               qP24_c4 <= qP24_c3;
               qM24_c4 <= qM24_c3;
               qP23_c4 <= qP23_c3;
               qM23_c4 <= qM23_c3;
               qP22_c4 <= qP22_c3;
               qM22_c4 <= qM22_c3;
               qP21_c4 <= qP21_c3;
               qM21_c4 <= qM21_c3;
               qP20_c4 <= qP20_c3;
               qM20_c4 <= qM20_c3;
               qP19_c4 <= qP19_c3;
               qM19_c4 <= qM19_c3;
               qP18_c4 <= qP18_c3;
               qM18_c4 <= qM18_c3;
               qP17_c4 <= qP17_c3;
               qM17_c4 <= qM17_c3;
               qP16_c4 <= qP16_c3;
               qM16_c4 <= qM16_c3;
               qP15_c4 <= qP15_c3;
               qM15_c4 <= qM15_c3;
               qP14_c4 <= qP14_c3;
               qM14_c4 <= qM14_c3;
               qP13_c4 <= qP13_c3;
               qM13_c4 <= qM13_c3;
               qP12_c4 <= qP12_c3;
               qM12_c4 <= qM12_c3;
               qP11_c4 <= qP11_c3;
               qM11_c4 <= qM11_c3;
            end if;
            if ce_5 = '1' then
               expR0_c5 <= expR0_c4;
               sR_c5 <= sR_c4;
               exnR0_c5 <= exnR0_c4;
               D_c5 <= D_c4;
               betaw6_c5 <= betaw6_c4;
               q6_copy27_c5 <= q6_copy27_c4;
               qP28_c5 <= qP28_c4;
               qM28_c5 <= qM28_c4;
               qP27_c5 <= qP27_c4;
               qM27_c5 <= qM27_c4;
               qP26_c5 <= qP26_c4;
               qM26_c5 <= qM26_c4;
               qP25_c5 <= qP25_c4;
               qM25_c5 <= qM25_c4;
               qP24_c5 <= qP24_c4;
               qM24_c5 <= qM24_c4;
               qP23_c5 <= qP23_c4;
               qM23_c5 <= qM23_c4;
               qP22_c5 <= qP22_c4;
               qM22_c5 <= qM22_c4;
               qP21_c5 <= qP21_c4;
               qM21_c5 <= qM21_c4;
               qP20_c5 <= qP20_c4;
               qM20_c5 <= qM20_c4;
               qP19_c5 <= qP19_c4;
               qM19_c5 <= qM19_c4;
               qP18_c5 <= qP18_c4;
               qM18_c5 <= qM18_c4;
               qP17_c5 <= qP17_c4;
               qM17_c5 <= qM17_c4;
               qP16_c5 <= qP16_c4;
               qM16_c5 <= qM16_c4;
               qP15_c5 <= qP15_c4;
               qM15_c5 <= qM15_c4;
               qP14_c5 <= qP14_c4;
               qM14_c5 <= qM14_c4;
               qP13_c5 <= qP13_c4;
               qM13_c5 <= qM13_c4;
               qP12_c5 <= qP12_c4;
               qM12_c5 <= qM12_c4;
               qP11_c5 <= qP11_c4;
               qM11_c5 <= qM11_c4;
               qP10_c5 <= qP10_c4;
               qM10_c5 <= qM10_c4;
               qP9_c5 <= qP9_c4;
               qM9_c5 <= qM9_c4;
               qP8_c5 <= qP8_c4;
               qM8_c5 <= qM8_c4;
               qP7_c5 <= qP7_c4;
               qM7_c5 <= qM7_c4;
            end if;
            if ce_6 = '1' then
               expR0_c6 <= expR0_c5;
               sR_c6 <= sR_c5;
               exnR0_c6 <= exnR0_c5;
               D_c6 <= D_c5;
               betaw2_c6 <= betaw2_c5;
               q2_c6 <= q2_c5;
               absq2D_c6 <= absq2D_c5;
               qP28_c6 <= qP28_c5;
               qM28_c6 <= qM28_c5;
               qP27_c6 <= qP27_c5;
               qM27_c6 <= qM27_c5;
               qP26_c6 <= qP26_c5;
               qM26_c6 <= qM26_c5;
               qP25_c6 <= qP25_c5;
               qM25_c6 <= qM25_c5;
               qP24_c6 <= qP24_c5;
               qM24_c6 <= qM24_c5;
               qP23_c6 <= qP23_c5;
               qM23_c6 <= qM23_c5;
               qP22_c6 <= qP22_c5;
               qM22_c6 <= qM22_c5;
               qP21_c6 <= qP21_c5;
               qM21_c6 <= qM21_c5;
               qP20_c6 <= qP20_c5;
               qM20_c6 <= qM20_c5;
               qP19_c6 <= qP19_c5;
               qM19_c6 <= qM19_c5;
               qP18_c6 <= qP18_c5;
               qM18_c6 <= qM18_c5;
               qP17_c6 <= qP17_c5;
               qM17_c6 <= qM17_c5;
               qP16_c6 <= qP16_c5;
               qM16_c6 <= qM16_c5;
               qP15_c6 <= qP15_c5;
               qM15_c6 <= qM15_c5;
               qP14_c6 <= qP14_c5;
               qM14_c6 <= qM14_c5;
               qP13_c6 <= qP13_c5;
               qM13_c6 <= qM13_c5;
               qP12_c6 <= qP12_c5;
               qM12_c6 <= qM12_c5;
               qP11_c6 <= qP11_c5;
               qM11_c6 <= qM11_c5;
               qP10_c6 <= qP10_c5;
               qM10_c6 <= qM10_c5;
               qP9_c6 <= qP9_c5;
               qM9_c6 <= qM9_c5;
               qP8_c6 <= qP8_c5;
               qM8_c6 <= qM8_c5;
               qP7_c6 <= qP7_c5;
               qM7_c6 <= qM7_c5;
               qP6_c6 <= qP6_c5;
               qM6_c6 <= qM6_c5;
               qP5_c6 <= qP5_c5;
               qM5_c6 <= qM5_c5;
               qP4_c6 <= qP4_c5;
               qM4_c6 <= qM4_c5;
               qP3_c6 <= qP3_c5;
               qM3_c6 <= qM3_c5;
               qP2_c6 <= qP2_c5;
               qM2_c6 <= qM2_c5;
            end if;
         end if;
      end process;
   fX_c0 <= "1" & X(51 downto 0);
   fY_c0 <= "1" & Y(51 downto 0);
   -- exponent difference, sign and exception combination computed early, to have fewer bits to pipeline
   expR0_c0 <= ("00" & X(62 downto 52)) - ("00" & Y(62 downto 52));
   sR_c0 <= X(63) xor Y(63);
   -- early exception handling 
   exnXY_c0 <= X(65 downto 64) & Y(65 downto 64);
   with exnXY_c0  select 
      exnR0_c0 <= 
         "01"	 when "0101",										-- normal
         "00"	 when "0001" | "0010" | "0110", -- zero
         "10"	 when "0100" | "1000" | "1001", -- overflow
         "11"	 when others;										-- NaN
   D_c0 <= fY_c0 ;
   psX_c0 <= "0" & fX_c0 ;
   betaw28_c0 <=  "00" & psX_c0;
   sel28_c0 <= betaw28_c0(55 downto 50) & D_c0(51 downto 49);
   SelFunctionTable28: selFunction_Freq100_uid4
      port map ( X => sel28_c0,
                 Y => q28_copy5_c0);
   q28_c0 <= q28_copy5_c0; -- output copy to hold a pipeline register if needed

   with q28_c0  select 
      absq28D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q28_c0(2)  select 
   w27_c0<= betaw28_c0 - absq28D_c0 when '0',
         betaw28_c0 + absq28D_c0 when others;

   betaw27_c0 <= w27_c0(53 downto 0) & "00"; -- multiplication by the radix
   sel27_c0 <= betaw27_c0(55 downto 50) & D_c0(51 downto 49);
   SelFunctionTable27: selFunction_Freq100_uid4
      port map ( X => sel27_c0,
                 Y => q27_copy6_c0);
   q27_c0 <= q27_copy6_c0; -- output copy to hold a pipeline register if needed

   with q27_c0  select 
      absq27D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q27_c0(2)  select 
   w26_c0<= betaw27_c0 - absq27D_c0 when '0',
         betaw27_c0 + absq27D_c0 when others;

   betaw26_c0 <= w26_c0(53 downto 0) & "00"; -- multiplication by the radix
   sel26_c0 <= betaw26_c0(55 downto 50) & D_c0(51 downto 49);
   SelFunctionTable26: selFunction_Freq100_uid4
      port map ( X => sel26_c0,
                 Y => q26_copy7_c0);
   q26_c0 <= q26_copy7_c0; -- output copy to hold a pipeline register if needed

   with q26_c0  select 
      absq26D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q26_c0(2)  select 
   w25_c0<= betaw26_c0 - absq26D_c0 when '0',
         betaw26_c0 + absq26D_c0 when others;

   betaw25_c0 <= w25_c0(53 downto 0) & "00"; -- multiplication by the radix
   sel25_c0 <= betaw25_c0(55 downto 50) & D_c0(51 downto 49);
   SelFunctionTable25: selFunction_Freq100_uid4
      port map ( X => sel25_c0,
                 Y => q25_copy8_c0);
   q25_c0 <= q25_copy8_c0; -- output copy to hold a pipeline register if needed

   with q25_c0  select 
      absq25D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q25_c0(2)  select 
   w24_c0<= betaw25_c0 - absq25D_c0 when '0',
         betaw25_c0 + absq25D_c0 when others;

   betaw24_c0 <= w24_c0(53 downto 0) & "00"; -- multiplication by the radix
   sel24_c0 <= betaw24_c0(55 downto 50) & D_c0(51 downto 49);
   SelFunctionTable24: selFunction_Freq100_uid4
      port map ( X => sel24_c0,
                 Y => q24_copy9_c0);
   q24_c0 <= q24_copy9_c0; -- output copy to hold a pipeline register if needed

   with q24_c0  select 
      absq24D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q24_c1(2)  select 
   w23_c1<= betaw24_c1 - absq24D_c1 when '0',
         betaw24_c1 + absq24D_c1 when others;

   betaw23_c1 <= w23_c1(53 downto 0) & "00"; -- multiplication by the radix
   sel23_c1 <= betaw23_c1(55 downto 50) & D_c1(51 downto 49);
   SelFunctionTable23: selFunction_Freq100_uid4
      port map ( X => sel23_c1,
                 Y => q23_copy10_c1);
   q23_c1 <= q23_copy10_c1; -- output copy to hold a pipeline register if needed

   with q23_c1  select 
      absq23D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q23_c1(2)  select 
   w22_c1<= betaw23_c1 - absq23D_c1 when '0',
         betaw23_c1 + absq23D_c1 when others;

   betaw22_c1 <= w22_c1(53 downto 0) & "00"; -- multiplication by the radix
   sel22_c1 <= betaw22_c1(55 downto 50) & D_c1(51 downto 49);
   SelFunctionTable22: selFunction_Freq100_uid4
      port map ( X => sel22_c1,
                 Y => q22_copy11_c1);
   q22_c1 <= q22_copy11_c1; -- output copy to hold a pipeline register if needed

   with q22_c1  select 
      absq22D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q22_c1(2)  select 
   w21_c1<= betaw22_c1 - absq22D_c1 when '0',
         betaw22_c1 + absq22D_c1 when others;

   betaw21_c1 <= w21_c1(53 downto 0) & "00"; -- multiplication by the radix
   sel21_c1 <= betaw21_c1(55 downto 50) & D_c1(51 downto 49);
   SelFunctionTable21: selFunction_Freq100_uid4
      port map ( X => sel21_c1,
                 Y => q21_copy12_c1);
   q21_c1 <= q21_copy12_c1; -- output copy to hold a pipeline register if needed

   with q21_c1  select 
      absq21D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q21_c1(2)  select 
   w20_c1<= betaw21_c1 - absq21D_c1 when '0',
         betaw21_c1 + absq21D_c1 when others;

   betaw20_c1 <= w20_c1(53 downto 0) & "00"; -- multiplication by the radix
   sel20_c1 <= betaw20_c1(55 downto 50) & D_c1(51 downto 49);
   SelFunctionTable20: selFunction_Freq100_uid4
      port map ( X => sel20_c1,
                 Y => q20_copy13_c1);
   q20_c1 <= q20_copy13_c1; -- output copy to hold a pipeline register if needed

   with q20_c1  select 
      absq20D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q20_c2(2)  select 
   w19_c2<= betaw20_c2 - absq20D_c2 when '0',
         betaw20_c2 + absq20D_c2 when others;

   betaw19_c2 <= w19_c2(53 downto 0) & "00"; -- multiplication by the radix
   sel19_c2 <= betaw19_c2(55 downto 50) & D_c2(51 downto 49);
   SelFunctionTable19: selFunction_Freq100_uid4
      port map ( X => sel19_c2,
                 Y => q19_copy14_c2);
   q19_c2 <= q19_copy14_c2; -- output copy to hold a pipeline register if needed

   with q19_c2  select 
      absq19D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q19_c2(2)  select 
   w18_c2<= betaw19_c2 - absq19D_c2 when '0',
         betaw19_c2 + absq19D_c2 when others;

   betaw18_c2 <= w18_c2(53 downto 0) & "00"; -- multiplication by the radix
   sel18_c2 <= betaw18_c2(55 downto 50) & D_c2(51 downto 49);
   SelFunctionTable18: selFunction_Freq100_uid4
      port map ( X => sel18_c2,
                 Y => q18_copy15_c2);
   q18_c2 <= q18_copy15_c2; -- output copy to hold a pipeline register if needed

   with q18_c2  select 
      absq18D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q18_c2(2)  select 
   w17_c2<= betaw18_c2 - absq18D_c2 when '0',
         betaw18_c2 + absq18D_c2 when others;

   betaw17_c2 <= w17_c2(53 downto 0) & "00"; -- multiplication by the radix
   sel17_c2 <= betaw17_c2(55 downto 50) & D_c2(51 downto 49);
   SelFunctionTable17: selFunction_Freq100_uid4
      port map ( X => sel17_c2,
                 Y => q17_copy16_c2);
   q17_c2 <= q17_copy16_c2; -- output copy to hold a pipeline register if needed

   with q17_c2  select 
      absq17D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q17_c2(2)  select 
   w16_c2<= betaw17_c2 - absq17D_c2 when '0',
         betaw17_c2 + absq17D_c2 when others;

   betaw16_c2 <= w16_c2(53 downto 0) & "00"; -- multiplication by the radix
   sel16_c2 <= betaw16_c2(55 downto 50) & D_c2(51 downto 49);
   SelFunctionTable16: selFunction_Freq100_uid4
      port map ( X => sel16_c2,
                 Y => q16_copy17_c2);
   q16_c2 <= q16_copy17_c2; -- output copy to hold a pipeline register if needed

   with q16_c2  select 
      absq16D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q16_c2(2)  select 
   w15_c2<= betaw16_c2 - absq16D_c2 when '0',
         betaw16_c2 + absq16D_c2 when others;

   betaw15_c2 <= w15_c2(53 downto 0) & "00"; -- multiplication by the radix
   sel15_c2 <= betaw15_c2(55 downto 50) & D_c2(51 downto 49);
   SelFunctionTable15: selFunction_Freq100_uid4
      port map ( X => sel15_c2,
                 Y => q15_copy18_c2);
   q15_c3 <= q15_copy18_c3; -- output copy to hold a pipeline register if needed

   with q15_c3  select 
      absq15D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q15_c3(2)  select 
   w14_c3<= betaw15_c3 - absq15D_c3 when '0',
         betaw15_c3 + absq15D_c3 when others;

   betaw14_c3 <= w14_c3(53 downto 0) & "00"; -- multiplication by the radix
   sel14_c3 <= betaw14_c3(55 downto 50) & D_c3(51 downto 49);
   SelFunctionTable14: selFunction_Freq100_uid4
      port map ( X => sel14_c3,
                 Y => q14_copy19_c3);
   q14_c3 <= q14_copy19_c3; -- output copy to hold a pipeline register if needed

   with q14_c3  select 
      absq14D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q14_c3(2)  select 
   w13_c3<= betaw14_c3 - absq14D_c3 when '0',
         betaw14_c3 + absq14D_c3 when others;

   betaw13_c3 <= w13_c3(53 downto 0) & "00"; -- multiplication by the radix
   sel13_c3 <= betaw13_c3(55 downto 50) & D_c3(51 downto 49);
   SelFunctionTable13: selFunction_Freq100_uid4
      port map ( X => sel13_c3,
                 Y => q13_copy20_c3);
   q13_c3 <= q13_copy20_c3; -- output copy to hold a pipeline register if needed

   with q13_c3  select 
      absq13D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q13_c3(2)  select 
   w12_c3<= betaw13_c3 - absq13D_c3 when '0',
         betaw13_c3 + absq13D_c3 when others;

   betaw12_c3 <= w12_c3(53 downto 0) & "00"; -- multiplication by the radix
   sel12_c3 <= betaw12_c3(55 downto 50) & D_c3(51 downto 49);
   SelFunctionTable12: selFunction_Freq100_uid4
      port map ( X => sel12_c3,
                 Y => q12_copy21_c3);
   q12_c3 <= q12_copy21_c3; -- output copy to hold a pipeline register if needed

   with q12_c3  select 
      absq12D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q12_c3(2)  select 
   w11_c3<= betaw12_c3 - absq12D_c3 when '0',
         betaw12_c3 + absq12D_c3 when others;

   betaw11_c3 <= w11_c3(53 downto 0) & "00"; -- multiplication by the radix
   sel11_c3 <= betaw11_c3(55 downto 50) & D_c3(51 downto 49);
   SelFunctionTable11: selFunction_Freq100_uid4
      port map ( X => sel11_c3,
                 Y => q11_copy22_c3);
   q11_c3 <= q11_copy22_c3; -- output copy to hold a pipeline register if needed

   with q11_c3  select 
      absq11D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q11_c4(2)  select 
   w10_c4<= betaw11_c4 - absq11D_c4 when '0',
         betaw11_c4 + absq11D_c4 when others;

   betaw10_c4 <= w10_c4(53 downto 0) & "00"; -- multiplication by the radix
   sel10_c4 <= betaw10_c4(55 downto 50) & D_c4(51 downto 49);
   SelFunctionTable10: selFunction_Freq100_uid4
      port map ( X => sel10_c4,
                 Y => q10_copy23_c4);
   q10_c4 <= q10_copy23_c4; -- output copy to hold a pipeline register if needed

   with q10_c4  select 
      absq10D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q10_c4(2)  select 
   w9_c4<= betaw10_c4 - absq10D_c4 when '0',
         betaw10_c4 + absq10D_c4 when others;

   betaw9_c4 <= w9_c4(53 downto 0) & "00"; -- multiplication by the radix
   sel9_c4 <= betaw9_c4(55 downto 50) & D_c4(51 downto 49);
   SelFunctionTable9: selFunction_Freq100_uid4
      port map ( X => sel9_c4,
                 Y => q9_copy24_c4);
   q9_c4 <= q9_copy24_c4; -- output copy to hold a pipeline register if needed

   with q9_c4  select 
      absq9D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q9_c4(2)  select 
   w8_c4<= betaw9_c4 - absq9D_c4 when '0',
         betaw9_c4 + absq9D_c4 when others;

   betaw8_c4 <= w8_c4(53 downto 0) & "00"; -- multiplication by the radix
   sel8_c4 <= betaw8_c4(55 downto 50) & D_c4(51 downto 49);
   SelFunctionTable8: selFunction_Freq100_uid4
      port map ( X => sel8_c4,
                 Y => q8_copy25_c4);
   q8_c4 <= q8_copy25_c4; -- output copy to hold a pipeline register if needed

   with q8_c4  select 
      absq8D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q8_c4(2)  select 
   w7_c4<= betaw8_c4 - absq8D_c4 when '0',
         betaw8_c4 + absq8D_c4 when others;

   betaw7_c4 <= w7_c4(53 downto 0) & "00"; -- multiplication by the radix
   sel7_c4 <= betaw7_c4(55 downto 50) & D_c4(51 downto 49);
   SelFunctionTable7: selFunction_Freq100_uid4
      port map ( X => sel7_c4,
                 Y => q7_copy26_c4);
   q7_c4 <= q7_copy26_c4; -- output copy to hold a pipeline register if needed

   with q7_c4  select 
      absq7D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q7_c4(2)  select 
   w6_c4<= betaw7_c4 - absq7D_c4 when '0',
         betaw7_c4 + absq7D_c4 when others;

   betaw6_c4 <= w6_c4(53 downto 0) & "00"; -- multiplication by the radix
   sel6_c4 <= betaw6_c4(55 downto 50) & D_c4(51 downto 49);
   SelFunctionTable6: selFunction_Freq100_uid4
      port map ( X => sel6_c4,
                 Y => q6_copy27_c4);
   q6_c5 <= q6_copy27_c5; -- output copy to hold a pipeline register if needed

   with q6_c5  select 
      absq6D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q6_c5(2)  select 
   w5_c5<= betaw6_c5 - absq6D_c5 when '0',
         betaw6_c5 + absq6D_c5 when others;

   betaw5_c5 <= w5_c5(53 downto 0) & "00"; -- multiplication by the radix
   sel5_c5 <= betaw5_c5(55 downto 50) & D_c5(51 downto 49);
   SelFunctionTable5: selFunction_Freq100_uid4
      port map ( X => sel5_c5,
                 Y => q5_copy28_c5);
   q5_c5 <= q5_copy28_c5; -- output copy to hold a pipeline register if needed

   with q5_c5  select 
      absq5D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q5_c5(2)  select 
   w4_c5<= betaw5_c5 - absq5D_c5 when '0',
         betaw5_c5 + absq5D_c5 when others;

   betaw4_c5 <= w4_c5(53 downto 0) & "00"; -- multiplication by the radix
   sel4_c5 <= betaw4_c5(55 downto 50) & D_c5(51 downto 49);
   SelFunctionTable4: selFunction_Freq100_uid4
      port map ( X => sel4_c5,
                 Y => q4_copy29_c5);
   q4_c5 <= q4_copy29_c5; -- output copy to hold a pipeline register if needed

   with q4_c5  select 
      absq4D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q4_c5(2)  select 
   w3_c5<= betaw4_c5 - absq4D_c5 when '0',
         betaw4_c5 + absq4D_c5 when others;

   betaw3_c5 <= w3_c5(53 downto 0) & "00"; -- multiplication by the radix
   sel3_c5 <= betaw3_c5(55 downto 50) & D_c5(51 downto 49);
   SelFunctionTable3: selFunction_Freq100_uid4
      port map ( X => sel3_c5,
                 Y => q3_copy30_c5);
   q3_c5 <= q3_copy30_c5; -- output copy to hold a pipeline register if needed

   with q3_c5  select 
      absq3D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q3_c5(2)  select 
   w2_c5<= betaw3_c5 - absq3D_c5 when '0',
         betaw3_c5 + absq3D_c5 when others;

   betaw2_c5 <= w2_c5(53 downto 0) & "00"; -- multiplication by the radix
   sel2_c5 <= betaw2_c5(55 downto 50) & D_c5(51 downto 49);
   SelFunctionTable2: selFunction_Freq100_uid4
      port map ( X => sel2_c5,
                 Y => q2_copy31_c5);
   q2_c5 <= q2_copy31_c5; -- output copy to hold a pipeline register if needed

   with q2_c5  select 
      absq2D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q2_c6(2)  select 
   w1_c6<= betaw2_c6 - absq2D_c6 when '0',
         betaw2_c6 + absq2D_c6 when others;

   betaw1_c6 <= w1_c6(53 downto 0) & "00"; -- multiplication by the radix
   sel1_c6 <= betaw1_c6(55 downto 50) & D_c6(51 downto 49);
   SelFunctionTable1: selFunction_Freq100_uid4
      port map ( X => sel1_c6,
                 Y => q1_copy32_c6);
   q1_c6 <= q1_copy32_c6; -- output copy to hold a pipeline register if needed

   with q1_c6  select 
      absq1D_c6 <= 
         "000" & D_c6						 when "001" | "111", -- mult by 1
         "00" & D_c6 & "0"			   when "010" | "110", -- mult by 2
         (55 downto 0 => '0')	 when others;        -- mult by 0

   with q1_c6(2)  select 
   w0_c6<= betaw1_c6 - absq1D_c6 when '0',
         betaw1_c6 + absq1D_c6 when others;

   wfinal_c6 <= w0_c6(53 downto 0);
   qM0_c6 <= wfinal_c6(53); -- rounding bit is the sign of the remainder
   qP28_c0 <=      q28_c0(1 downto 0);
   qM28_c0 <=      q28_c0(2) & "0";
   qP27_c0 <=      q27_c0(1 downto 0);
   qM27_c0 <=      q27_c0(2) & "0";
   qP26_c0 <=      q26_c0(1 downto 0);
   qM26_c0 <=      q26_c0(2) & "0";
   qP25_c0 <=      q25_c0(1 downto 0);
   qM25_c0 <=      q25_c0(2) & "0";
   qP24_c0 <=      q24_c0(1 downto 0);
   qM24_c0 <=      q24_c0(2) & "0";
   qP23_c1 <=      q23_c1(1 downto 0);
   qM23_c1 <=      q23_c1(2) & "0";
   qP22_c1 <=      q22_c1(1 downto 0);
   qM22_c1 <=      q22_c1(2) & "0";
   qP21_c1 <=      q21_c1(1 downto 0);
   qM21_c1 <=      q21_c1(2) & "0";
   qP20_c1 <=      q20_c1(1 downto 0);
   qM20_c1 <=      q20_c1(2) & "0";
   qP19_c2 <=      q19_c2(1 downto 0);
   qM19_c2 <=      q19_c2(2) & "0";
   qP18_c2 <=      q18_c2(1 downto 0);
   qM18_c2 <=      q18_c2(2) & "0";
   qP17_c2 <=      q17_c2(1 downto 0);
   qM17_c2 <=      q17_c2(2) & "0";
   qP16_c2 <=      q16_c2(1 downto 0);
   qM16_c2 <=      q16_c2(2) & "0";
   qP15_c3 <=      q15_c3(1 downto 0);
   qM15_c3 <=      q15_c3(2) & "0";
   qP14_c3 <=      q14_c3(1 downto 0);
   qM14_c3 <=      q14_c3(2) & "0";
   qP13_c3 <=      q13_c3(1 downto 0);
   qM13_c3 <=      q13_c3(2) & "0";
   qP12_c3 <=      q12_c3(1 downto 0);
   qM12_c3 <=      q12_c3(2) & "0";
   qP11_c3 <=      q11_c3(1 downto 0);
   qM11_c3 <=      q11_c3(2) & "0";
   qP10_c4 <=      q10_c4(1 downto 0);
   qM10_c4 <=      q10_c4(2) & "0";
   qP9_c4 <=      q9_c4(1 downto 0);
   qM9_c4 <=      q9_c4(2) & "0";
   qP8_c4 <=      q8_c4(1 downto 0);
   qM8_c4 <=      q8_c4(2) & "0";
   qP7_c4 <=      q7_c4(1 downto 0);
   qM7_c4 <=      q7_c4(2) & "0";
   qP6_c5 <=      q6_c5(1 downto 0);
   qM6_c5 <=      q6_c5(2) & "0";
   qP5_c5 <=      q5_c5(1 downto 0);
   qM5_c5 <=      q5_c5(2) & "0";
   qP4_c5 <=      q4_c5(1 downto 0);
   qM4_c5 <=      q4_c5(2) & "0";
   qP3_c5 <=      q3_c5(1 downto 0);
   qM3_c5 <=      q3_c5(2) & "0";
   qP2_c5 <=      q2_c5(1 downto 0);
   qM2_c5 <=      q2_c5(2) & "0";
   qP1_c6 <=      q1_c6(1 downto 0);
   qM1_c6 <=      q1_c6(2) & "0";
   qP_c6 <= qP28_c6 & qP27_c6 & qP26_c6 & qP25_c6 & qP24_c6 & qP23_c6 & qP22_c6 & qP21_c6 & qP20_c6 & qP19_c6 & qP18_c6 & qP17_c6 & qP16_c6 & qP15_c6 & qP14_c6 & qP13_c6 & qP12_c6 & qP11_c6 & qP10_c6 & qP9_c6 & qP8_c6 & qP7_c6 & qP6_c6 & qP5_c6 & qP4_c6 & qP3_c6 & qP2_c6 & qP1_c6;
   qM_c6 <= qM28_c6(0) & qM27_c6 & qM26_c6 & qM25_c6 & qM24_c6 & qM23_c6 & qM22_c6 & qM21_c6 & qM20_c6 & qM19_c6 & qM18_c6 & qM17_c6 & qM16_c6 & qM15_c6 & qM14_c6 & qM13_c6 & qM12_c6 & qM11_c6 & qM10_c6 & qM9_c6 & qM8_c6 & qM7_c6 & qM6_c6 & qM5_c6 & qM4_c6 & qM3_c6 & qM2_c6 & qM1_c6 & qM0_c6;
   quotient_c6 <= qP_c6 - qM_c6;
   -- We need a mR in (0, -wf-2) format: 1+wF fraction bits, 1 round bit, and 1 guard bit for the normalisation,
   -- quotient is the truncation of the exact quotient to at least 2^(-wF-2) bits
   -- now discarding its possible known MSB zeroes, and dropping the possible extra LSB bit (due to radix 4) 
   mR_c6 <= quotient_c6(54 downto 0); 
   -- normalisation
   fRnorm_c6 <=    mR_c6(53 downto 1)  when mR_c6(54)= '1'
           else mR_c6(52 downto 0);  -- now fRnorm is a (-1, -wF-1) fraction
   round_c6 <= fRnorm_c6(0); 
   expR1_c6 <= expR0_c6 + ("000" & (9 downto 1 => '1') & mR_c6(54)); -- add back bias
   -- final rounding
   expfrac_c6 <= expR1_c6 & fRnorm_c6(52 downto 1) ;
   expfracR_c6 <= expfrac_c6 + ((64 downto 1 => '0') & round_c6);
   exnR_c6 <=      "00"  when expfracR_c6(64) = '1'   -- underflow
           else "10"  when  expfracR_c6(64 downto 63) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_c6  select 
      exnRfinal_c6 <= 
         exnR_c6   when "01", -- normal
         exnR0_c6  when others;
   R <= exnRfinal_c6 & sR_c6 & expfracR_c6(62 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          selFunction_Freq500_uid4
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity selFunction_Freq500_uid4 is
    port (X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of selFunction_Freq500_uid4 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000000000",
      "000" when "000000001",
      "000" when "000000010",
      "000" when "000000011",
      "000" when "000000100",
      "000" when "000000101",
      "000" when "000000110",
      "000" when "000000111",
      "000" when "000001000",
      "000" when "000001001",
      "000" when "000001010",
      "000" when "000001011",
      "000" when "000001100",
      "000" when "000001101",
      "000" when "000001110",
      "000" when "000001111",
      "001" when "000010000",
      "000" when "000010001",
      "000" when "000010010",
      "000" when "000010011",
      "000" when "000010100",
      "000" when "000010101",
      "000" when "000010110",
      "000" when "000010111",
      "001" when "000011000",
      "001" when "000011001",
      "001" when "000011010",
      "001" when "000011011",
      "000" when "000011100",
      "000" when "000011101",
      "000" when "000011110",
      "000" when "000011111",
      "001" when "000100000",
      "001" when "000100001",
      "001" when "000100010",
      "001" when "000100011",
      "001" when "000100100",
      "001" when "000100101",
      "001" when "000100110",
      "000" when "000100111",
      "001" when "000101000",
      "001" when "000101001",
      "001" when "000101010",
      "001" when "000101011",
      "001" when "000101100",
      "001" when "000101101",
      "001" when "000101110",
      "001" when "000101111",
      "010" when "000110000",
      "001" when "000110001",
      "001" when "000110010",
      "001" when "000110011",
      "001" when "000110100",
      "001" when "000110101",
      "001" when "000110110",
      "001" when "000110111",
      "010" when "000111000",
      "010" when "000111001",
      "001" when "000111010",
      "001" when "000111011",
      "001" when "000111100",
      "001" when "000111101",
      "001" when "000111110",
      "001" when "000111111",
      "010" when "001000000",
      "010" when "001000001",
      "010" when "001000010",
      "001" when "001000011",
      "001" when "001000100",
      "001" when "001000101",
      "001" when "001000110",
      "001" when "001000111",
      "010" when "001001000",
      "010" when "001001001",
      "010" when "001001010",
      "010" when "001001011",
      "001" when "001001100",
      "001" when "001001101",
      "001" when "001001110",
      "001" when "001001111",
      "010" when "001010000",
      "010" when "001010001",
      "010" when "001010010",
      "010" when "001010011",
      "010" when "001010100",
      "010" when "001010101",
      "001" when "001010110",
      "001" when "001010111",
      "010" when "001011000",
      "010" when "001011001",
      "010" when "001011010",
      "010" when "001011011",
      "010" when "001011100",
      "010" when "001011101",
      "010" when "001011110",
      "001" when "001011111",
      "010" when "001100000",
      "010" when "001100001",
      "010" when "001100010",
      "010" when "001100011",
      "010" when "001100100",
      "010" when "001100101",
      "010" when "001100110",
      "010" when "001100111",
      "010" when "001101000",
      "010" when "001101001",
      "010" when "001101010",
      "010" when "001101011",
      "010" when "001101100",
      "010" when "001101101",
      "010" when "001101110",
      "010" when "001101111",
      "010" when "001110000",
      "010" when "001110001",
      "010" when "001110010",
      "010" when "001110011",
      "010" when "001110100",
      "010" when "001110101",
      "010" when "001110110",
      "010" when "001110111",
      "010" when "001111000",
      "010" when "001111001",
      "010" when "001111010",
      "010" when "001111011",
      "010" when "001111100",
      "010" when "001111101",
      "010" when "001111110",
      "010" when "001111111",
      "010" when "010000000",
      "010" when "010000001",
      "010" when "010000010",
      "010" when "010000011",
      "010" when "010000100",
      "010" when "010000101",
      "010" when "010000110",
      "010" when "010000111",
      "010" when "010001000",
      "010" when "010001001",
      "010" when "010001010",
      "010" when "010001011",
      "010" when "010001100",
      "010" when "010001101",
      "010" when "010001110",
      "010" when "010001111",
      "010" when "010010000",
      "010" when "010010001",
      "010" when "010010010",
      "010" when "010010011",
      "010" when "010010100",
      "010" when "010010101",
      "010" when "010010110",
      "010" when "010010111",
      "010" when "010011000",
      "010" when "010011001",
      "010" when "010011010",
      "010" when "010011011",
      "010" when "010011100",
      "010" when "010011101",
      "010" when "010011110",
      "010" when "010011111",
      "010" when "010100000",
      "010" when "010100001",
      "010" when "010100010",
      "010" when "010100011",
      "010" when "010100100",
      "010" when "010100101",
      "010" when "010100110",
      "010" when "010100111",
      "010" when "010101000",
      "010" when "010101001",
      "010" when "010101010",
      "010" when "010101011",
      "010" when "010101100",
      "010" when "010101101",
      "010" when "010101110",
      "010" when "010101111",
      "010" when "010110000",
      "010" when "010110001",
      "010" when "010110010",
      "010" when "010110011",
      "010" when "010110100",
      "010" when "010110101",
      "010" when "010110110",
      "010" when "010110111",
      "010" when "010111000",
      "010" when "010111001",
      "010" when "010111010",
      "010" when "010111011",
      "010" when "010111100",
      "010" when "010111101",
      "010" when "010111110",
      "010" when "010111111",
      "010" when "011000000",
      "010" when "011000001",
      "010" when "011000010",
      "010" when "011000011",
      "010" when "011000100",
      "010" when "011000101",
      "010" when "011000110",
      "010" when "011000111",
      "010" when "011001000",
      "010" when "011001001",
      "010" when "011001010",
      "010" when "011001011",
      "010" when "011001100",
      "010" when "011001101",
      "010" when "011001110",
      "010" when "011001111",
      "010" when "011010000",
      "010" when "011010001",
      "010" when "011010010",
      "010" when "011010011",
      "010" when "011010100",
      "010" when "011010101",
      "010" when "011010110",
      "010" when "011010111",
      "010" when "011011000",
      "010" when "011011001",
      "010" when "011011010",
      "010" when "011011011",
      "010" when "011011100",
      "010" when "011011101",
      "010" when "011011110",
      "010" when "011011111",
      "010" when "011100000",
      "010" when "011100001",
      "010" when "011100010",
      "010" when "011100011",
      "010" when "011100100",
      "010" when "011100101",
      "010" when "011100110",
      "010" when "011100111",
      "010" when "011101000",
      "010" when "011101001",
      "010" when "011101010",
      "010" when "011101011",
      "010" when "011101100",
      "010" when "011101101",
      "010" when "011101110",
      "010" when "011101111",
      "010" when "011110000",
      "010" when "011110001",
      "010" when "011110010",
      "010" when "011110011",
      "010" when "011110100",
      "010" when "011110101",
      "010" when "011110110",
      "010" when "011110111",
      "010" when "011111000",
      "010" when "011111001",
      "010" when "011111010",
      "010" when "011111011",
      "010" when "011111100",
      "010" when "011111101",
      "010" when "011111110",
      "010" when "011111111",
      "110" when "100000000",
      "110" when "100000001",
      "110" when "100000010",
      "110" when "100000011",
      "110" when "100000100",
      "110" when "100000101",
      "110" when "100000110",
      "110" when "100000111",
      "110" when "100001000",
      "110" when "100001001",
      "110" when "100001010",
      "110" when "100001011",
      "110" when "100001100",
      "110" when "100001101",
      "110" when "100001110",
      "110" when "100001111",
      "110" when "100010000",
      "110" when "100010001",
      "110" when "100010010",
      "110" when "100010011",
      "110" when "100010100",
      "110" when "100010101",
      "110" when "100010110",
      "110" when "100010111",
      "110" when "100011000",
      "110" when "100011001",
      "110" when "100011010",
      "110" when "100011011",
      "110" when "100011100",
      "110" when "100011101",
      "110" when "100011110",
      "110" when "100011111",
      "110" when "100100000",
      "110" when "100100001",
      "110" when "100100010",
      "110" when "100100011",
      "110" when "100100100",
      "110" when "100100101",
      "110" when "100100110",
      "110" when "100100111",
      "110" when "100101000",
      "110" when "100101001",
      "110" when "100101010",
      "110" when "100101011",
      "110" when "100101100",
      "110" when "100101101",
      "110" when "100101110",
      "110" when "100101111",
      "110" when "100110000",
      "110" when "100110001",
      "110" when "100110010",
      "110" when "100110011",
      "110" when "100110100",
      "110" when "100110101",
      "110" when "100110110",
      "110" when "100110111",
      "110" when "100111000",
      "110" when "100111001",
      "110" when "100111010",
      "110" when "100111011",
      "110" when "100111100",
      "110" when "100111101",
      "110" when "100111110",
      "110" when "100111111",
      "110" when "101000000",
      "110" when "101000001",
      "110" when "101000010",
      "110" when "101000011",
      "110" when "101000100",
      "110" when "101000101",
      "110" when "101000110",
      "110" when "101000111",
      "110" when "101001000",
      "110" when "101001001",
      "110" when "101001010",
      "110" when "101001011",
      "110" when "101001100",
      "110" when "101001101",
      "110" when "101001110",
      "110" when "101001111",
      "110" when "101010000",
      "110" when "101010001",
      "110" when "101010010",
      "110" when "101010011",
      "110" when "101010100",
      "110" when "101010101",
      "110" when "101010110",
      "110" when "101010111",
      "110" when "101011000",
      "110" when "101011001",
      "110" when "101011010",
      "110" when "101011011",
      "110" when "101011100",
      "110" when "101011101",
      "110" when "101011110",
      "110" when "101011111",
      "110" when "101100000",
      "110" when "101100001",
      "110" when "101100010",
      "110" when "101100011",
      "110" when "101100100",
      "110" when "101100101",
      "110" when "101100110",
      "110" when "101100111",
      "110" when "101101000",
      "110" when "101101001",
      "110" when "101101010",
      "110" when "101101011",
      "110" when "101101100",
      "110" when "101101101",
      "110" when "101101110",
      "110" when "101101111",
      "110" when "101110000",
      "110" when "101110001",
      "110" when "101110010",
      "110" when "101110011",
      "110" when "101110100",
      "110" when "101110101",
      "110" when "101110110",
      "110" when "101110111",
      "110" when "101111000",
      "110" when "101111001",
      "110" when "101111010",
      "110" when "101111011",
      "110" when "101111100",
      "110" when "101111101",
      "110" when "101111110",
      "110" when "101111111",
      "110" when "110000000",
      "110" when "110000001",
      "110" when "110000010",
      "110" when "110000011",
      "110" when "110000100",
      "110" when "110000101",
      "110" when "110000110",
      "110" when "110000111",
      "110" when "110001000",
      "110" when "110001001",
      "110" when "110001010",
      "110" when "110001011",
      "110" when "110001100",
      "110" when "110001101",
      "110" when "110001110",
      "110" when "110001111",
      "110" when "110010000",
      "110" when "110010001",
      "110" when "110010010",
      "110" when "110010011",
      "110" when "110010100",
      "110" when "110010101",
      "110" when "110010110",
      "110" when "110010111",
      "110" when "110011000",
      "110" when "110011001",
      "110" when "110011010",
      "110" when "110011011",
      "110" when "110011100",
      "110" when "110011101",
      "110" when "110011110",
      "110" when "110011111",
      "110" when "110100000",
      "110" when "110100001",
      "110" when "110100010",
      "110" when "110100011",
      "110" when "110100100",
      "110" when "110100101",
      "110" when "110100110",
      "110" when "110100111",
      "110" when "110101000",
      "110" when "110101001",
      "110" when "110101010",
      "110" when "110101011",
      "110" when "110101100",
      "110" when "110101101",
      "110" when "110101110",
      "111" when "110101111",
      "110" when "110110000",
      "110" when "110110001",
      "110" when "110110010",
      "110" when "110110011",
      "110" when "110110100",
      "111" when "110110101",
      "111" when "110110110",
      "111" when "110110111",
      "110" when "110111000",
      "110" when "110111001",
      "110" when "110111010",
      "110" when "110111011",
      "111" when "110111100",
      "111" when "110111101",
      "111" when "110111110",
      "111" when "110111111",
      "110" when "111000000",
      "110" when "111000001",
      "111" when "111000010",
      "111" when "111000011",
      "111" when "111000100",
      "111" when "111000101",
      "111" when "111000110",
      "111" when "111000111",
      "110" when "111001000",
      "111" when "111001001",
      "111" when "111001010",
      "111" when "111001011",
      "111" when "111001100",
      "111" when "111001101",
      "111" when "111001110",
      "111" when "111001111",
      "111" when "111010000",
      "111" when "111010001",
      "111" when "111010010",
      "111" when "111010011",
      "111" when "111010100",
      "111" when "111010101",
      "111" when "111010110",
      "111" when "111010111",
      "111" when "111011000",
      "111" when "111011001",
      "111" when "111011010",
      "111" when "111011011",
      "111" when "111011100",
      "111" when "111011101",
      "111" when "111011110",
      "111" when "111011111",
      "111" when "111100000",
      "111" when "111100001",
      "111" when "111100010",
      "111" when "111100011",
      "111" when "111100100",
      "111" when "111100101",
      "111" when "111100110",
      "111" when "111100111",
      "111" when "111101000",
      "111" when "111101001",
      "111" when "111101010",
      "111" when "111101011",
      "000" when "111101100",
      "000" when "111101101",
      "000" when "111101110",
      "000" when "111101111",
      "000" when "111110000",
      "000" when "111110001",
      "000" when "111110010",
      "000" when "111110011",
      "000" when "111110100",
      "000" when "111110101",
      "000" when "111110110",
      "000" when "111110111",
      "000" when "111111000",
      "000" when "111111001",
      "000" when "111111010",
      "000" when "111111011",
      "000" when "111111100",
      "000" when "111111101",
      "000" when "111111110",
      "000" when "111111111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            FloatingPointDivider
--                         (FPDiv_8_23_Freq500_uid2)
-- VHDL generated for Kintex7 @ 500MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 15 cycles
-- Clock period (ns): 2
-- Target frequency (MHz): 500
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointDivider_32_3_812000 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9, ce_10, ce_11, ce_12, ce_13, ce_14, ce_15 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointDivider_32_3_812000 is
   component selFunction_Freq500_uid4 is
      port ( X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal fX_c0 :  std_logic_vector(23 downto 0);
signal fY_c0 :  std_logic_vector(23 downto 0);
signal expR0_c0, expR0_c1, expR0_c2, expR0_c3, expR0_c4, expR0_c5, expR0_c6, expR0_c7, expR0_c8, expR0_c9, expR0_c10, expR0_c11, expR0_c12, expR0_c13, expR0_c14, expR0_c15 :  std_logic_vector(9 downto 0);
signal sR_c0, sR_c1, sR_c2, sR_c3, sR_c4, sR_c5, sR_c6, sR_c7, sR_c8, sR_c9, sR_c10, sR_c11, sR_c12, sR_c13, sR_c14, sR_c15 :  std_logic;
signal exnXY_c0 :  std_logic_vector(3 downto 0);
signal exnR0_c0, exnR0_c1, exnR0_c2, exnR0_c3, exnR0_c4, exnR0_c5, exnR0_c6, exnR0_c7, exnR0_c8, exnR0_c9, exnR0_c10, exnR0_c11, exnR0_c12, exnR0_c13, exnR0_c14, exnR0_c15 :  std_logic_vector(1 downto 0);
signal D_c0, D_c1, D_c2, D_c3, D_c4, D_c5, D_c6, D_c7, D_c8, D_c9, D_c10, D_c11, D_c12, D_c13 :  std_logic_vector(23 downto 0);
signal psX_c0 :  std_logic_vector(24 downto 0);
signal betaw14_c0, betaw14_c1 :  std_logic_vector(26 downto 0);
signal sel14_c0 :  std_logic_vector(8 downto 0);
signal q14_c0, q14_c1 :  std_logic_vector(2 downto 0);
signal q14_copy5_c0 :  std_logic_vector(2 downto 0);
signal absq14D_c0, absq14D_c1 :  std_logic_vector(26 downto 0);
signal w13_c1 :  std_logic_vector(26 downto 0);
signal betaw13_c1, betaw13_c2 :  std_logic_vector(26 downto 0);
signal sel13_c1 :  std_logic_vector(8 downto 0);
signal q13_c1, q13_c2 :  std_logic_vector(2 downto 0);
signal q13_copy6_c1 :  std_logic_vector(2 downto 0);
signal absq13D_c1, absq13D_c2 :  std_logic_vector(26 downto 0);
signal w12_c2 :  std_logic_vector(26 downto 0);
signal betaw12_c2, betaw12_c3 :  std_logic_vector(26 downto 0);
signal sel12_c2 :  std_logic_vector(8 downto 0);
signal q12_c2, q12_c3 :  std_logic_vector(2 downto 0);
signal q12_copy7_c2 :  std_logic_vector(2 downto 0);
signal absq12D_c2, absq12D_c3 :  std_logic_vector(26 downto 0);
signal w11_c3 :  std_logic_vector(26 downto 0);
signal betaw11_c3, betaw11_c4 :  std_logic_vector(26 downto 0);
signal sel11_c3 :  std_logic_vector(8 downto 0);
signal q11_c3, q11_c4 :  std_logic_vector(2 downto 0);
signal q11_copy8_c3 :  std_logic_vector(2 downto 0);
signal absq11D_c3, absq11D_c4 :  std_logic_vector(26 downto 0);
signal w10_c4 :  std_logic_vector(26 downto 0);
signal betaw10_c4, betaw10_c5 :  std_logic_vector(26 downto 0);
signal sel10_c4 :  std_logic_vector(8 downto 0);
signal q10_c4, q10_c5 :  std_logic_vector(2 downto 0);
signal q10_copy9_c4 :  std_logic_vector(2 downto 0);
signal absq10D_c4, absq10D_c5 :  std_logic_vector(26 downto 0);
signal w9_c5 :  std_logic_vector(26 downto 0);
signal betaw9_c5, betaw9_c6 :  std_logic_vector(26 downto 0);
signal sel9_c5 :  std_logic_vector(8 downto 0);
signal q9_c5, q9_c6 :  std_logic_vector(2 downto 0);
signal q9_copy10_c5 :  std_logic_vector(2 downto 0);
signal absq9D_c5, absq9D_c6 :  std_logic_vector(26 downto 0);
signal w8_c6 :  std_logic_vector(26 downto 0);
signal betaw8_c6, betaw8_c7 :  std_logic_vector(26 downto 0);
signal sel8_c6 :  std_logic_vector(8 downto 0);
signal q8_c6, q8_c7 :  std_logic_vector(2 downto 0);
signal q8_copy11_c6 :  std_logic_vector(2 downto 0);
signal absq8D_c6, absq8D_c7 :  std_logic_vector(26 downto 0);
signal w7_c7 :  std_logic_vector(26 downto 0);
signal betaw7_c7, betaw7_c8 :  std_logic_vector(26 downto 0);
signal sel7_c7 :  std_logic_vector(8 downto 0);
signal q7_c7, q7_c8 :  std_logic_vector(2 downto 0);
signal q7_copy12_c7 :  std_logic_vector(2 downto 0);
signal absq7D_c7, absq7D_c8 :  std_logic_vector(26 downto 0);
signal w6_c8 :  std_logic_vector(26 downto 0);
signal betaw6_c8, betaw6_c9 :  std_logic_vector(26 downto 0);
signal sel6_c8 :  std_logic_vector(8 downto 0);
signal q6_c8, q6_c9 :  std_logic_vector(2 downto 0);
signal q6_copy13_c8 :  std_logic_vector(2 downto 0);
signal absq6D_c8, absq6D_c9 :  std_logic_vector(26 downto 0);
signal w5_c9 :  std_logic_vector(26 downto 0);
signal betaw5_c9, betaw5_c10 :  std_logic_vector(26 downto 0);
signal sel5_c9 :  std_logic_vector(8 downto 0);
signal q5_c9, q5_c10 :  std_logic_vector(2 downto 0);
signal q5_copy14_c9 :  std_logic_vector(2 downto 0);
signal absq5D_c9, absq5D_c10 :  std_logic_vector(26 downto 0);
signal w4_c10 :  std_logic_vector(26 downto 0);
signal betaw4_c10, betaw4_c11 :  std_logic_vector(26 downto 0);
signal sel4_c10 :  std_logic_vector(8 downto 0);
signal q4_c10, q4_c11 :  std_logic_vector(2 downto 0);
signal q4_copy15_c10 :  std_logic_vector(2 downto 0);
signal absq4D_c10, absq4D_c11 :  std_logic_vector(26 downto 0);
signal w3_c11 :  std_logic_vector(26 downto 0);
signal betaw3_c11, betaw3_c12 :  std_logic_vector(26 downto 0);
signal sel3_c11 :  std_logic_vector(8 downto 0);
signal q3_c11, q3_c12 :  std_logic_vector(2 downto 0);
signal q3_copy16_c11 :  std_logic_vector(2 downto 0);
signal absq3D_c11, absq3D_c12 :  std_logic_vector(26 downto 0);
signal w2_c12 :  std_logic_vector(26 downto 0);
signal betaw2_c12, betaw2_c13 :  std_logic_vector(26 downto 0);
signal sel2_c12 :  std_logic_vector(8 downto 0);
signal q2_c12, q2_c13 :  std_logic_vector(2 downto 0);
signal q2_copy17_c12 :  std_logic_vector(2 downto 0);
signal absq2D_c12, absq2D_c13 :  std_logic_vector(26 downto 0);
signal w1_c13 :  std_logic_vector(26 downto 0);
signal betaw1_c13, betaw1_c14 :  std_logic_vector(26 downto 0);
signal sel1_c13 :  std_logic_vector(8 downto 0);
signal q1_c13, q1_c14 :  std_logic_vector(2 downto 0);
signal q1_copy18_c13 :  std_logic_vector(2 downto 0);
signal absq1D_c13, absq1D_c14 :  std_logic_vector(26 downto 0);
signal w0_c14 :  std_logic_vector(26 downto 0);
signal wfinal_c14 :  std_logic_vector(24 downto 0);
signal qM0_c14 :  std_logic;
signal qP14_c0, qP14_c1, qP14_c2, qP14_c3, qP14_c4, qP14_c5, qP14_c6, qP14_c7, qP14_c8, qP14_c9, qP14_c10, qP14_c11, qP14_c12, qP14_c13 :  std_logic_vector(1 downto 0);
signal qM14_c0, qM14_c1, qM14_c2, qM14_c3, qM14_c4, qM14_c5, qM14_c6, qM14_c7, qM14_c8, qM14_c9, qM14_c10, qM14_c11, qM14_c12, qM14_c13, qM14_c14 :  std_logic_vector(1 downto 0);
signal qP13_c1, qP13_c2, qP13_c3, qP13_c4, qP13_c5, qP13_c6, qP13_c7, qP13_c8, qP13_c9, qP13_c10, qP13_c11, qP13_c12, qP13_c13 :  std_logic_vector(1 downto 0);
signal qM13_c1, qM13_c2, qM13_c3, qM13_c4, qM13_c5, qM13_c6, qM13_c7, qM13_c8, qM13_c9, qM13_c10, qM13_c11, qM13_c12, qM13_c13, qM13_c14 :  std_logic_vector(1 downto 0);
signal qP12_c2, qP12_c3, qP12_c4, qP12_c5, qP12_c6, qP12_c7, qP12_c8, qP12_c9, qP12_c10, qP12_c11, qP12_c12, qP12_c13 :  std_logic_vector(1 downto 0);
signal qM12_c2, qM12_c3, qM12_c4, qM12_c5, qM12_c6, qM12_c7, qM12_c8, qM12_c9, qM12_c10, qM12_c11, qM12_c12, qM12_c13, qM12_c14 :  std_logic_vector(1 downto 0);
signal qP11_c3, qP11_c4, qP11_c5, qP11_c6, qP11_c7, qP11_c8, qP11_c9, qP11_c10, qP11_c11, qP11_c12, qP11_c13 :  std_logic_vector(1 downto 0);
signal qM11_c3, qM11_c4, qM11_c5, qM11_c6, qM11_c7, qM11_c8, qM11_c9, qM11_c10, qM11_c11, qM11_c12, qM11_c13, qM11_c14 :  std_logic_vector(1 downto 0);
signal qP10_c4, qP10_c5, qP10_c6, qP10_c7, qP10_c8, qP10_c9, qP10_c10, qP10_c11, qP10_c12, qP10_c13 :  std_logic_vector(1 downto 0);
signal qM10_c4, qM10_c5, qM10_c6, qM10_c7, qM10_c8, qM10_c9, qM10_c10, qM10_c11, qM10_c12, qM10_c13, qM10_c14 :  std_logic_vector(1 downto 0);
signal qP9_c5, qP9_c6, qP9_c7, qP9_c8, qP9_c9, qP9_c10, qP9_c11, qP9_c12, qP9_c13 :  std_logic_vector(1 downto 0);
signal qM9_c5, qM9_c6, qM9_c7, qM9_c8, qM9_c9, qM9_c10, qM9_c11, qM9_c12, qM9_c13, qM9_c14 :  std_logic_vector(1 downto 0);
signal qP8_c6, qP8_c7, qP8_c8, qP8_c9, qP8_c10, qP8_c11, qP8_c12, qP8_c13 :  std_logic_vector(1 downto 0);
signal qM8_c6, qM8_c7, qM8_c8, qM8_c9, qM8_c10, qM8_c11, qM8_c12, qM8_c13, qM8_c14 :  std_logic_vector(1 downto 0);
signal qP7_c7, qP7_c8, qP7_c9, qP7_c10, qP7_c11, qP7_c12, qP7_c13 :  std_logic_vector(1 downto 0);
signal qM7_c7, qM7_c8, qM7_c9, qM7_c10, qM7_c11, qM7_c12, qM7_c13, qM7_c14 :  std_logic_vector(1 downto 0);
signal qP6_c8, qP6_c9, qP6_c10, qP6_c11, qP6_c12, qP6_c13 :  std_logic_vector(1 downto 0);
signal qM6_c8, qM6_c9, qM6_c10, qM6_c11, qM6_c12, qM6_c13, qM6_c14 :  std_logic_vector(1 downto 0);
signal qP5_c9, qP5_c10, qP5_c11, qP5_c12, qP5_c13 :  std_logic_vector(1 downto 0);
signal qM5_c9, qM5_c10, qM5_c11, qM5_c12, qM5_c13, qM5_c14 :  std_logic_vector(1 downto 0);
signal qP4_c10, qP4_c11, qP4_c12, qP4_c13 :  std_logic_vector(1 downto 0);
signal qM4_c10, qM4_c11, qM4_c12, qM4_c13, qM4_c14 :  std_logic_vector(1 downto 0);
signal qP3_c11, qP3_c12, qP3_c13 :  std_logic_vector(1 downto 0);
signal qM3_c11, qM3_c12, qM3_c13, qM3_c14 :  std_logic_vector(1 downto 0);
signal qP2_c12, qP2_c13 :  std_logic_vector(1 downto 0);
signal qM2_c12, qM2_c13, qM2_c14 :  std_logic_vector(1 downto 0);
signal qP1_c13 :  std_logic_vector(1 downto 0);
signal qM1_c13, qM1_c14 :  std_logic_vector(1 downto 0);
signal qP_c13, qP_c14, qP_c15 :  std_logic_vector(27 downto 0);
signal qM_c14, qM_c15 :  std_logic_vector(27 downto 0);
signal quotient_c15 :  std_logic_vector(27 downto 0);
signal mR_c15 :  std_logic_vector(25 downto 0);
signal fRnorm_c15 :  std_logic_vector(23 downto 0);
signal round_c15 :  std_logic;
signal expR1_c15 :  std_logic_vector(9 downto 0);
signal expfrac_c15 :  std_logic_vector(32 downto 0);
signal expfracR_c15 :  std_logic_vector(32 downto 0);
signal exnR_c15 :  std_logic_vector(1 downto 0);
signal exnRfinal_c15 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               expR0_c1 <= expR0_c0;
               sR_c1 <= sR_c0;
               exnR0_c1 <= exnR0_c0;
               D_c1 <= D_c0;
               betaw14_c1 <= betaw14_c0;
               q14_c1 <= q14_c0;
               absq14D_c1 <= absq14D_c0;
               qP14_c1 <= qP14_c0;
               qM14_c1 <= qM14_c0;
            end if;
            if ce_2 = '1' then
               expR0_c2 <= expR0_c1;
               sR_c2 <= sR_c1;
               exnR0_c2 <= exnR0_c1;
               D_c2 <= D_c1;
               betaw13_c2 <= betaw13_c1;
               q13_c2 <= q13_c1;
               absq13D_c2 <= absq13D_c1;
               qP14_c2 <= qP14_c1;
               qM14_c2 <= qM14_c1;
               qP13_c2 <= qP13_c1;
               qM13_c2 <= qM13_c1;
            end if;
            if ce_3 = '1' then
               expR0_c3 <= expR0_c2;
               sR_c3 <= sR_c2;
               exnR0_c3 <= exnR0_c2;
               D_c3 <= D_c2;
               betaw12_c3 <= betaw12_c2;
               q12_c3 <= q12_c2;
               absq12D_c3 <= absq12D_c2;
               qP14_c3 <= qP14_c2;
               qM14_c3 <= qM14_c2;
               qP13_c3 <= qP13_c2;
               qM13_c3 <= qM13_c2;
               qP12_c3 <= qP12_c2;
               qM12_c3 <= qM12_c2;
            end if;
            if ce_4 = '1' then
               expR0_c4 <= expR0_c3;
               sR_c4 <= sR_c3;
               exnR0_c4 <= exnR0_c3;
               D_c4 <= D_c3;
               betaw11_c4 <= betaw11_c3;
               q11_c4 <= q11_c3;
               absq11D_c4 <= absq11D_c3;
               qP14_c4 <= qP14_c3;
               qM14_c4 <= qM14_c3;
               qP13_c4 <= qP13_c3;
               qM13_c4 <= qM13_c3;
               qP12_c4 <= qP12_c3;
               qM12_c4 <= qM12_c3;
               qP11_c4 <= qP11_c3;
               qM11_c4 <= qM11_c3;
            end if;
            if ce_5 = '1' then
               expR0_c5 <= expR0_c4;
               sR_c5 <= sR_c4;
               exnR0_c5 <= exnR0_c4;
               D_c5 <= D_c4;
               betaw10_c5 <= betaw10_c4;
               q10_c5 <= q10_c4;
               absq10D_c5 <= absq10D_c4;
               qP14_c5 <= qP14_c4;
               qM14_c5 <= qM14_c4;
               qP13_c5 <= qP13_c4;
               qM13_c5 <= qM13_c4;
               qP12_c5 <= qP12_c4;
               qM12_c5 <= qM12_c4;
               qP11_c5 <= qP11_c4;
               qM11_c5 <= qM11_c4;
               qP10_c5 <= qP10_c4;
               qM10_c5 <= qM10_c4;
            end if;
            if ce_6 = '1' then
               expR0_c6 <= expR0_c5;
               sR_c6 <= sR_c5;
               exnR0_c6 <= exnR0_c5;
               D_c6 <= D_c5;
               betaw9_c6 <= betaw9_c5;
               q9_c6 <= q9_c5;
               absq9D_c6 <= absq9D_c5;
               qP14_c6 <= qP14_c5;
               qM14_c6 <= qM14_c5;
               qP13_c6 <= qP13_c5;
               qM13_c6 <= qM13_c5;
               qP12_c6 <= qP12_c5;
               qM12_c6 <= qM12_c5;
               qP11_c6 <= qP11_c5;
               qM11_c6 <= qM11_c5;
               qP10_c6 <= qP10_c5;
               qM10_c6 <= qM10_c5;
               qP9_c6 <= qP9_c5;
               qM9_c6 <= qM9_c5;
            end if;
            if ce_7 = '1' then
               expR0_c7 <= expR0_c6;
               sR_c7 <= sR_c6;
               exnR0_c7 <= exnR0_c6;
               D_c7 <= D_c6;
               betaw8_c7 <= betaw8_c6;
               q8_c7 <= q8_c6;
               absq8D_c7 <= absq8D_c6;
               qP14_c7 <= qP14_c6;
               qM14_c7 <= qM14_c6;
               qP13_c7 <= qP13_c6;
               qM13_c7 <= qM13_c6;
               qP12_c7 <= qP12_c6;
               qM12_c7 <= qM12_c6;
               qP11_c7 <= qP11_c6;
               qM11_c7 <= qM11_c6;
               qP10_c7 <= qP10_c6;
               qM10_c7 <= qM10_c6;
               qP9_c7 <= qP9_c6;
               qM9_c7 <= qM9_c6;
               qP8_c7 <= qP8_c6;
               qM8_c7 <= qM8_c6;
            end if;
            if ce_8 = '1' then
               expR0_c8 <= expR0_c7;
               sR_c8 <= sR_c7;
               exnR0_c8 <= exnR0_c7;
               D_c8 <= D_c7;
               betaw7_c8 <= betaw7_c7;
               q7_c8 <= q7_c7;
               absq7D_c8 <= absq7D_c7;
               qP14_c8 <= qP14_c7;
               qM14_c8 <= qM14_c7;
               qP13_c8 <= qP13_c7;
               qM13_c8 <= qM13_c7;
               qP12_c8 <= qP12_c7;
               qM12_c8 <= qM12_c7;
               qP11_c8 <= qP11_c7;
               qM11_c8 <= qM11_c7;
               qP10_c8 <= qP10_c7;
               qM10_c8 <= qM10_c7;
               qP9_c8 <= qP9_c7;
               qM9_c8 <= qM9_c7;
               qP8_c8 <= qP8_c7;
               qM8_c8 <= qM8_c7;
               qP7_c8 <= qP7_c7;
               qM7_c8 <= qM7_c7;
            end if;
            if ce_9 = '1' then
               expR0_c9 <= expR0_c8;
               sR_c9 <= sR_c8;
               exnR0_c9 <= exnR0_c8;
               D_c9 <= D_c8;
               betaw6_c9 <= betaw6_c8;
               q6_c9 <= q6_c8;
               absq6D_c9 <= absq6D_c8;
               qP14_c9 <= qP14_c8;
               qM14_c9 <= qM14_c8;
               qP13_c9 <= qP13_c8;
               qM13_c9 <= qM13_c8;
               qP12_c9 <= qP12_c8;
               qM12_c9 <= qM12_c8;
               qP11_c9 <= qP11_c8;
               qM11_c9 <= qM11_c8;
               qP10_c9 <= qP10_c8;
               qM10_c9 <= qM10_c8;
               qP9_c9 <= qP9_c8;
               qM9_c9 <= qM9_c8;
               qP8_c9 <= qP8_c8;
               qM8_c9 <= qM8_c8;
               qP7_c9 <= qP7_c8;
               qM7_c9 <= qM7_c8;
               qP6_c9 <= qP6_c8;
               qM6_c9 <= qM6_c8;
            end if;
            if ce_10 = '1' then
               expR0_c10 <= expR0_c9;
               sR_c10 <= sR_c9;
               exnR0_c10 <= exnR0_c9;
               D_c10 <= D_c9;
               betaw5_c10 <= betaw5_c9;
               q5_c10 <= q5_c9;
               absq5D_c10 <= absq5D_c9;
               qP14_c10 <= qP14_c9;
               qM14_c10 <= qM14_c9;
               qP13_c10 <= qP13_c9;
               qM13_c10 <= qM13_c9;
               qP12_c10 <= qP12_c9;
               qM12_c10 <= qM12_c9;
               qP11_c10 <= qP11_c9;
               qM11_c10 <= qM11_c9;
               qP10_c10 <= qP10_c9;
               qM10_c10 <= qM10_c9;
               qP9_c10 <= qP9_c9;
               qM9_c10 <= qM9_c9;
               qP8_c10 <= qP8_c9;
               qM8_c10 <= qM8_c9;
               qP7_c10 <= qP7_c9;
               qM7_c10 <= qM7_c9;
               qP6_c10 <= qP6_c9;
               qM6_c10 <= qM6_c9;
               qP5_c10 <= qP5_c9;
               qM5_c10 <= qM5_c9;
            end if;
            if ce_11 = '1' then
               expR0_c11 <= expR0_c10;
               sR_c11 <= sR_c10;
               exnR0_c11 <= exnR0_c10;
               D_c11 <= D_c10;
               betaw4_c11 <= betaw4_c10;
               q4_c11 <= q4_c10;
               absq4D_c11 <= absq4D_c10;
               qP14_c11 <= qP14_c10;
               qM14_c11 <= qM14_c10;
               qP13_c11 <= qP13_c10;
               qM13_c11 <= qM13_c10;
               qP12_c11 <= qP12_c10;
               qM12_c11 <= qM12_c10;
               qP11_c11 <= qP11_c10;
               qM11_c11 <= qM11_c10;
               qP10_c11 <= qP10_c10;
               qM10_c11 <= qM10_c10;
               qP9_c11 <= qP9_c10;
               qM9_c11 <= qM9_c10;
               qP8_c11 <= qP8_c10;
               qM8_c11 <= qM8_c10;
               qP7_c11 <= qP7_c10;
               qM7_c11 <= qM7_c10;
               qP6_c11 <= qP6_c10;
               qM6_c11 <= qM6_c10;
               qP5_c11 <= qP5_c10;
               qM5_c11 <= qM5_c10;
               qP4_c11 <= qP4_c10;
               qM4_c11 <= qM4_c10;
            end if;
            if ce_12 = '1' then
               expR0_c12 <= expR0_c11;
               sR_c12 <= sR_c11;
               exnR0_c12 <= exnR0_c11;
               D_c12 <= D_c11;
               betaw3_c12 <= betaw3_c11;
               q3_c12 <= q3_c11;
               absq3D_c12 <= absq3D_c11;
               qP14_c12 <= qP14_c11;
               qM14_c12 <= qM14_c11;
               qP13_c12 <= qP13_c11;
               qM13_c12 <= qM13_c11;
               qP12_c12 <= qP12_c11;
               qM12_c12 <= qM12_c11;
               qP11_c12 <= qP11_c11;
               qM11_c12 <= qM11_c11;
               qP10_c12 <= qP10_c11;
               qM10_c12 <= qM10_c11;
               qP9_c12 <= qP9_c11;
               qM9_c12 <= qM9_c11;
               qP8_c12 <= qP8_c11;
               qM8_c12 <= qM8_c11;
               qP7_c12 <= qP7_c11;
               qM7_c12 <= qM7_c11;
               qP6_c12 <= qP6_c11;
               qM6_c12 <= qM6_c11;
               qP5_c12 <= qP5_c11;
               qM5_c12 <= qM5_c11;
               qP4_c12 <= qP4_c11;
               qM4_c12 <= qM4_c11;
               qP3_c12 <= qP3_c11;
               qM3_c12 <= qM3_c11;
            end if;
            if ce_13 = '1' then
               expR0_c13 <= expR0_c12;
               sR_c13 <= sR_c12;
               exnR0_c13 <= exnR0_c12;
               D_c13 <= D_c12;
               betaw2_c13 <= betaw2_c12;
               q2_c13 <= q2_c12;
               absq2D_c13 <= absq2D_c12;
               qP14_c13 <= qP14_c12;
               qM14_c13 <= qM14_c12;
               qP13_c13 <= qP13_c12;
               qM13_c13 <= qM13_c12;
               qP12_c13 <= qP12_c12;
               qM12_c13 <= qM12_c12;
               qP11_c13 <= qP11_c12;
               qM11_c13 <= qM11_c12;
               qP10_c13 <= qP10_c12;
               qM10_c13 <= qM10_c12;
               qP9_c13 <= qP9_c12;
               qM9_c13 <= qM9_c12;
               qP8_c13 <= qP8_c12;
               qM8_c13 <= qM8_c12;
               qP7_c13 <= qP7_c12;
               qM7_c13 <= qM7_c12;
               qP6_c13 <= qP6_c12;
               qM6_c13 <= qM6_c12;
               qP5_c13 <= qP5_c12;
               qM5_c13 <= qM5_c12;
               qP4_c13 <= qP4_c12;
               qM4_c13 <= qM4_c12;
               qP3_c13 <= qP3_c12;
               qM3_c13 <= qM3_c12;
               qP2_c13 <= qP2_c12;
               qM2_c13 <= qM2_c12;
            end if;
            if ce_14 = '1' then
               expR0_c14 <= expR0_c13;
               sR_c14 <= sR_c13;
               exnR0_c14 <= exnR0_c13;
               betaw1_c14 <= betaw1_c13;
               q1_c14 <= q1_c13;
               absq1D_c14 <= absq1D_c13;
               qM14_c14 <= qM14_c13;
               qM13_c14 <= qM13_c13;
               qM12_c14 <= qM12_c13;
               qM11_c14 <= qM11_c13;
               qM10_c14 <= qM10_c13;
               qM9_c14 <= qM9_c13;
               qM8_c14 <= qM8_c13;
               qM7_c14 <= qM7_c13;
               qM6_c14 <= qM6_c13;
               qM5_c14 <= qM5_c13;
               qM4_c14 <= qM4_c13;
               qM3_c14 <= qM3_c13;
               qM2_c14 <= qM2_c13;
               qM1_c14 <= qM1_c13;
               qP_c14 <= qP_c13;
            end if;
            if ce_15 = '1' then
               expR0_c15 <= expR0_c14;
               sR_c15 <= sR_c14;
               exnR0_c15 <= exnR0_c14;
               qP_c15 <= qP_c14;
               qM_c15 <= qM_c14;
            end if;
         end if;
      end process;
   fX_c0 <= "1" & X(22 downto 0);
   fY_c0 <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have fewer bits to pipeline
   expR0_c0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR_c0 <= X(31) xor Y(31);
   -- early exception handling 
   exnXY_c0 <= X(33 downto 32) & Y(33 downto 32);
   with exnXY_c0  select 
      exnR0_c0 <= 
         "01"	 when "0101",										-- normal
         "00"	 when "0001" | "0010" | "0110", -- zero
         "10"	 when "0100" | "1000" | "1001", -- overflow
         "11"	 when others;										-- NaN
   D_c0 <= fY_c0 ;
   psX_c0 <= "0" & fX_c0 ;
   betaw14_c0 <=  "00" & psX_c0;
   sel14_c0 <= betaw14_c0(26 downto 21) & D_c0(22 downto 20);
   SelFunctionTable14: selFunction_Freq500_uid4
      port map ( X => sel14_c0,
                 Y => q14_copy5_c0);
   q14_c0 <= q14_copy5_c0; -- output copy to hold a pipeline register if needed

   with q14_c0  select 
      absq14D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q14_c1(2)  select 
   w13_c1<= betaw14_c1 - absq14D_c1 when '0',
         betaw14_c1 + absq14D_c1 when others;

   betaw13_c1 <= w13_c1(24 downto 0) & "00"; -- multiplication by the radix
   sel13_c1 <= betaw13_c1(26 downto 21) & D_c1(22 downto 20);
   SelFunctionTable13: selFunction_Freq500_uid4
      port map ( X => sel13_c1,
                 Y => q13_copy6_c1);
   q13_c1 <= q13_copy6_c1; -- output copy to hold a pipeline register if needed

   with q13_c1  select 
      absq13D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q13_c2(2)  select 
   w12_c2<= betaw13_c2 - absq13D_c2 when '0',
         betaw13_c2 + absq13D_c2 when others;

   betaw12_c2 <= w12_c2(24 downto 0) & "00"; -- multiplication by the radix
   sel12_c2 <= betaw12_c2(26 downto 21) & D_c2(22 downto 20);
   SelFunctionTable12: selFunction_Freq500_uid4
      port map ( X => sel12_c2,
                 Y => q12_copy7_c2);
   q12_c2 <= q12_copy7_c2; -- output copy to hold a pipeline register if needed

   with q12_c2  select 
      absq12D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q12_c3(2)  select 
   w11_c3<= betaw12_c3 - absq12D_c3 when '0',
         betaw12_c3 + absq12D_c3 when others;

   betaw11_c3 <= w11_c3(24 downto 0) & "00"; -- multiplication by the radix
   sel11_c3 <= betaw11_c3(26 downto 21) & D_c3(22 downto 20);
   SelFunctionTable11: selFunction_Freq500_uid4
      port map ( X => sel11_c3,
                 Y => q11_copy8_c3);
   q11_c3 <= q11_copy8_c3; -- output copy to hold a pipeline register if needed

   with q11_c3  select 
      absq11D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q11_c4(2)  select 
   w10_c4<= betaw11_c4 - absq11D_c4 when '0',
         betaw11_c4 + absq11D_c4 when others;

   betaw10_c4 <= w10_c4(24 downto 0) & "00"; -- multiplication by the radix
   sel10_c4 <= betaw10_c4(26 downto 21) & D_c4(22 downto 20);
   SelFunctionTable10: selFunction_Freq500_uid4
      port map ( X => sel10_c4,
                 Y => q10_copy9_c4);
   q10_c4 <= q10_copy9_c4; -- output copy to hold a pipeline register if needed

   with q10_c4  select 
      absq10D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q10_c5(2)  select 
   w9_c5<= betaw10_c5 - absq10D_c5 when '0',
         betaw10_c5 + absq10D_c5 when others;

   betaw9_c5 <= w9_c5(24 downto 0) & "00"; -- multiplication by the radix
   sel9_c5 <= betaw9_c5(26 downto 21) & D_c5(22 downto 20);
   SelFunctionTable9: selFunction_Freq500_uid4
      port map ( X => sel9_c5,
                 Y => q9_copy10_c5);
   q9_c5 <= q9_copy10_c5; -- output copy to hold a pipeline register if needed

   with q9_c5  select 
      absq9D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q9_c6(2)  select 
   w8_c6<= betaw9_c6 - absq9D_c6 when '0',
         betaw9_c6 + absq9D_c6 when others;

   betaw8_c6 <= w8_c6(24 downto 0) & "00"; -- multiplication by the radix
   sel8_c6 <= betaw8_c6(26 downto 21) & D_c6(22 downto 20);
   SelFunctionTable8: selFunction_Freq500_uid4
      port map ( X => sel8_c6,
                 Y => q8_copy11_c6);
   q8_c6 <= q8_copy11_c6; -- output copy to hold a pipeline register if needed

   with q8_c6  select 
      absq8D_c6 <= 
         "000" & D_c6						 when "001" | "111", -- mult by 1
         "00" & D_c6 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q8_c7(2)  select 
   w7_c7<= betaw8_c7 - absq8D_c7 when '0',
         betaw8_c7 + absq8D_c7 when others;

   betaw7_c7 <= w7_c7(24 downto 0) & "00"; -- multiplication by the radix
   sel7_c7 <= betaw7_c7(26 downto 21) & D_c7(22 downto 20);
   SelFunctionTable7: selFunction_Freq500_uid4
      port map ( X => sel7_c7,
                 Y => q7_copy12_c7);
   q7_c7 <= q7_copy12_c7; -- output copy to hold a pipeline register if needed

   with q7_c7  select 
      absq7D_c7 <= 
         "000" & D_c7						 when "001" | "111", -- mult by 1
         "00" & D_c7 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q7_c8(2)  select 
   w6_c8<= betaw7_c8 - absq7D_c8 when '0',
         betaw7_c8 + absq7D_c8 when others;

   betaw6_c8 <= w6_c8(24 downto 0) & "00"; -- multiplication by the radix
   sel6_c8 <= betaw6_c8(26 downto 21) & D_c8(22 downto 20);
   SelFunctionTable6: selFunction_Freq500_uid4
      port map ( X => sel6_c8,
                 Y => q6_copy13_c8);
   q6_c8 <= q6_copy13_c8; -- output copy to hold a pipeline register if needed

   with q6_c8  select 
      absq6D_c8 <= 
         "000" & D_c8						 when "001" | "111", -- mult by 1
         "00" & D_c8 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q6_c9(2)  select 
   w5_c9<= betaw6_c9 - absq6D_c9 when '0',
         betaw6_c9 + absq6D_c9 when others;

   betaw5_c9 <= w5_c9(24 downto 0) & "00"; -- multiplication by the radix
   sel5_c9 <= betaw5_c9(26 downto 21) & D_c9(22 downto 20);
   SelFunctionTable5: selFunction_Freq500_uid4
      port map ( X => sel5_c9,
                 Y => q5_copy14_c9);
   q5_c9 <= q5_copy14_c9; -- output copy to hold a pipeline register if needed

   with q5_c9  select 
      absq5D_c9 <= 
         "000" & D_c9						 when "001" | "111", -- mult by 1
         "00" & D_c9 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q5_c10(2)  select 
   w4_c10<= betaw5_c10 - absq5D_c10 when '0',
         betaw5_c10 + absq5D_c10 when others;

   betaw4_c10 <= w4_c10(24 downto 0) & "00"; -- multiplication by the radix
   sel4_c10 <= betaw4_c10(26 downto 21) & D_c10(22 downto 20);
   SelFunctionTable4: selFunction_Freq500_uid4
      port map ( X => sel4_c10,
                 Y => q4_copy15_c10);
   q4_c10 <= q4_copy15_c10; -- output copy to hold a pipeline register if needed

   with q4_c10  select 
      absq4D_c10 <= 
         "000" & D_c10						 when "001" | "111", -- mult by 1
         "00" & D_c10 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q4_c11(2)  select 
   w3_c11<= betaw4_c11 - absq4D_c11 when '0',
         betaw4_c11 + absq4D_c11 when others;

   betaw3_c11 <= w3_c11(24 downto 0) & "00"; -- multiplication by the radix
   sel3_c11 <= betaw3_c11(26 downto 21) & D_c11(22 downto 20);
   SelFunctionTable3: selFunction_Freq500_uid4
      port map ( X => sel3_c11,
                 Y => q3_copy16_c11);
   q3_c11 <= q3_copy16_c11; -- output copy to hold a pipeline register if needed

   with q3_c11  select 
      absq3D_c11 <= 
         "000" & D_c11						 when "001" | "111", -- mult by 1
         "00" & D_c11 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q3_c12(2)  select 
   w2_c12<= betaw3_c12 - absq3D_c12 when '0',
         betaw3_c12 + absq3D_c12 when others;

   betaw2_c12 <= w2_c12(24 downto 0) & "00"; -- multiplication by the radix
   sel2_c12 <= betaw2_c12(26 downto 21) & D_c12(22 downto 20);
   SelFunctionTable2: selFunction_Freq500_uid4
      port map ( X => sel2_c12,
                 Y => q2_copy17_c12);
   q2_c12 <= q2_copy17_c12; -- output copy to hold a pipeline register if needed

   with q2_c12  select 
      absq2D_c12 <= 
         "000" & D_c12						 when "001" | "111", -- mult by 1
         "00" & D_c12 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q2_c13(2)  select 
   w1_c13<= betaw2_c13 - absq2D_c13 when '0',
         betaw2_c13 + absq2D_c13 when others;

   betaw1_c13 <= w1_c13(24 downto 0) & "00"; -- multiplication by the radix
   sel1_c13 <= betaw1_c13(26 downto 21) & D_c13(22 downto 20);
   SelFunctionTable1: selFunction_Freq500_uid4
      port map ( X => sel1_c13,
                 Y => q1_copy18_c13);
   q1_c13 <= q1_copy18_c13; -- output copy to hold a pipeline register if needed

   with q1_c13  select 
      absq1D_c13 <= 
         "000" & D_c13						 when "001" | "111", -- mult by 1
         "00" & D_c13 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q1_c14(2)  select 
   w0_c14<= betaw1_c14 - absq1D_c14 when '0',
         betaw1_c14 + absq1D_c14 when others;

   wfinal_c14 <= w0_c14(24 downto 0);
   qM0_c14 <= wfinal_c14(24); -- rounding bit is the sign of the remainder
   qP14_c0 <=      q14_c0(1 downto 0);
   qM14_c0 <=      q14_c0(2) & "0";
   qP13_c1 <=      q13_c1(1 downto 0);
   qM13_c1 <=      q13_c1(2) & "0";
   qP12_c2 <=      q12_c2(1 downto 0);
   qM12_c2 <=      q12_c2(2) & "0";
   qP11_c3 <=      q11_c3(1 downto 0);
   qM11_c3 <=      q11_c3(2) & "0";
   qP10_c4 <=      q10_c4(1 downto 0);
   qM10_c4 <=      q10_c4(2) & "0";
   qP9_c5 <=      q9_c5(1 downto 0);
   qM9_c5 <=      q9_c5(2) & "0";
   qP8_c6 <=      q8_c6(1 downto 0);
   qM8_c6 <=      q8_c6(2) & "0";
   qP7_c7 <=      q7_c7(1 downto 0);
   qM7_c7 <=      q7_c7(2) & "0";
   qP6_c8 <=      q6_c8(1 downto 0);
   qM6_c8 <=      q6_c8(2) & "0";
   qP5_c9 <=      q5_c9(1 downto 0);
   qM5_c9 <=      q5_c9(2) & "0";
   qP4_c10 <=      q4_c10(1 downto 0);
   qM4_c10 <=      q4_c10(2) & "0";
   qP3_c11 <=      q3_c11(1 downto 0);
   qM3_c11 <=      q3_c11(2) & "0";
   qP2_c12 <=      q2_c12(1 downto 0);
   qM2_c12 <=      q2_c12(2) & "0";
   qP1_c13 <=      q1_c13(1 downto 0);
   qM1_c13 <=      q1_c13(2) & "0";
   qP_c13 <= qP14_c13 & qP13_c13 & qP12_c13 & qP11_c13 & qP10_c13 & qP9_c13 & qP8_c13 & qP7_c13 & qP6_c13 & qP5_c13 & qP4_c13 & qP3_c13 & qP2_c13 & qP1_c13;
   qM_c14 <= qM14_c14(0) & qM13_c14 & qM12_c14 & qM11_c14 & qM10_c14 & qM9_c14 & qM8_c14 & qM7_c14 & qM6_c14 & qM5_c14 & qM4_c14 & qM3_c14 & qM2_c14 & qM1_c14 & qM0_c14;
   quotient_c15 <= qP_c15 - qM_c15;
   -- We need a mR in (0, -wf-2) format: 1+wF fraction bits, 1 round bit, and 1 guard bit for the normalisation,
   -- quotient is the truncation of the exact quotient to at least 2^(-wF-2) bits
   -- now discarding its possible known MSB zeroes, and dropping the possible extra LSB bit (due to radix 4) 
   mR_c15 <= quotient_c15(26 downto 1); 
   -- normalisation
   fRnorm_c15 <=    mR_c15(24 downto 1)  when mR_c15(25)= '1'
           else mR_c15(23 downto 0);  -- now fRnorm is a (-1, -wF-1) fraction
   round_c15 <= fRnorm_c15(0); 
   expR1_c15 <= expR0_c15 + ("000" & (6 downto 1 => '1') & mR_c15(25)); -- add back bias
   -- final rounding
   expfrac_c15 <= expR1_c15 & fRnorm_c15(23 downto 1) ;
   expfracR_c15 <= expfrac_c15 + ((32 downto 1 => '0') & round_c15);
   exnR_c15 <=      "00"  when expfracR_c15(32) = '1'   -- underflow
           else "10"  when  expfracR_c15(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_c15  select 
      exnRfinal_c15 <= 
         exnR_c15   when "01", -- normal
         exnR0_c15  when others;
   R <= exnRfinal_c15 & sR_c15 & expfracR_c15(30 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          selFunction_Freq300_uid4
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity selFunction_Freq300_uid4 is
    port (X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of selFunction_Freq300_uid4 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000000000",
      "000" when "000000001",
      "000" when "000000010",
      "000" when "000000011",
      "000" when "000000100",
      "000" when "000000101",
      "000" when "000000110",
      "000" when "000000111",
      "000" when "000001000",
      "000" when "000001001",
      "000" when "000001010",
      "000" when "000001011",
      "000" when "000001100",
      "000" when "000001101",
      "000" when "000001110",
      "000" when "000001111",
      "001" when "000010000",
      "000" when "000010001",
      "000" when "000010010",
      "000" when "000010011",
      "000" when "000010100",
      "000" when "000010101",
      "000" when "000010110",
      "000" when "000010111",
      "001" when "000011000",
      "001" when "000011001",
      "001" when "000011010",
      "001" when "000011011",
      "000" when "000011100",
      "000" when "000011101",
      "000" when "000011110",
      "000" when "000011111",
      "001" when "000100000",
      "001" when "000100001",
      "001" when "000100010",
      "001" when "000100011",
      "001" when "000100100",
      "001" when "000100101",
      "001" when "000100110",
      "000" when "000100111",
      "001" when "000101000",
      "001" when "000101001",
      "001" when "000101010",
      "001" when "000101011",
      "001" when "000101100",
      "001" when "000101101",
      "001" when "000101110",
      "001" when "000101111",
      "010" when "000110000",
      "001" when "000110001",
      "001" when "000110010",
      "001" when "000110011",
      "001" when "000110100",
      "001" when "000110101",
      "001" when "000110110",
      "001" when "000110111",
      "010" when "000111000",
      "010" when "000111001",
      "001" when "000111010",
      "001" when "000111011",
      "001" when "000111100",
      "001" when "000111101",
      "001" when "000111110",
      "001" when "000111111",
      "010" when "001000000",
      "010" when "001000001",
      "010" when "001000010",
      "001" when "001000011",
      "001" when "001000100",
      "001" when "001000101",
      "001" when "001000110",
      "001" when "001000111",
      "010" when "001001000",
      "010" when "001001001",
      "010" when "001001010",
      "010" when "001001011",
      "001" when "001001100",
      "001" when "001001101",
      "001" when "001001110",
      "001" when "001001111",
      "010" when "001010000",
      "010" when "001010001",
      "010" when "001010010",
      "010" when "001010011",
      "010" when "001010100",
      "010" when "001010101",
      "001" when "001010110",
      "001" when "001010111",
      "010" when "001011000",
      "010" when "001011001",
      "010" when "001011010",
      "010" when "001011011",
      "010" when "001011100",
      "010" when "001011101",
      "010" when "001011110",
      "001" when "001011111",
      "010" when "001100000",
      "010" when "001100001",
      "010" when "001100010",
      "010" when "001100011",
      "010" when "001100100",
      "010" when "001100101",
      "010" when "001100110",
      "010" when "001100111",
      "010" when "001101000",
      "010" when "001101001",
      "010" when "001101010",
      "010" when "001101011",
      "010" when "001101100",
      "010" when "001101101",
      "010" when "001101110",
      "010" when "001101111",
      "010" when "001110000",
      "010" when "001110001",
      "010" when "001110010",
      "010" when "001110011",
      "010" when "001110100",
      "010" when "001110101",
      "010" when "001110110",
      "010" when "001110111",
      "010" when "001111000",
      "010" when "001111001",
      "010" when "001111010",
      "010" when "001111011",
      "010" when "001111100",
      "010" when "001111101",
      "010" when "001111110",
      "010" when "001111111",
      "010" when "010000000",
      "010" when "010000001",
      "010" when "010000010",
      "010" when "010000011",
      "010" when "010000100",
      "010" when "010000101",
      "010" when "010000110",
      "010" when "010000111",
      "010" when "010001000",
      "010" when "010001001",
      "010" when "010001010",
      "010" when "010001011",
      "010" when "010001100",
      "010" when "010001101",
      "010" when "010001110",
      "010" when "010001111",
      "010" when "010010000",
      "010" when "010010001",
      "010" when "010010010",
      "010" when "010010011",
      "010" when "010010100",
      "010" when "010010101",
      "010" when "010010110",
      "010" when "010010111",
      "010" when "010011000",
      "010" when "010011001",
      "010" when "010011010",
      "010" when "010011011",
      "010" when "010011100",
      "010" when "010011101",
      "010" when "010011110",
      "010" when "010011111",
      "010" when "010100000",
      "010" when "010100001",
      "010" when "010100010",
      "010" when "010100011",
      "010" when "010100100",
      "010" when "010100101",
      "010" when "010100110",
      "010" when "010100111",
      "010" when "010101000",
      "010" when "010101001",
      "010" when "010101010",
      "010" when "010101011",
      "010" when "010101100",
      "010" when "010101101",
      "010" when "010101110",
      "010" when "010101111",
      "010" when "010110000",
      "010" when "010110001",
      "010" when "010110010",
      "010" when "010110011",
      "010" when "010110100",
      "010" when "010110101",
      "010" when "010110110",
      "010" when "010110111",
      "010" when "010111000",
      "010" when "010111001",
      "010" when "010111010",
      "010" when "010111011",
      "010" when "010111100",
      "010" when "010111101",
      "010" when "010111110",
      "010" when "010111111",
      "010" when "011000000",
      "010" when "011000001",
      "010" when "011000010",
      "010" when "011000011",
      "010" when "011000100",
      "010" when "011000101",
      "010" when "011000110",
      "010" when "011000111",
      "010" when "011001000",
      "010" when "011001001",
      "010" when "011001010",
      "010" when "011001011",
      "010" when "011001100",
      "010" when "011001101",
      "010" when "011001110",
      "010" when "011001111",
      "010" when "011010000",
      "010" when "011010001",
      "010" when "011010010",
      "010" when "011010011",
      "010" when "011010100",
      "010" when "011010101",
      "010" when "011010110",
      "010" when "011010111",
      "010" when "011011000",
      "010" when "011011001",
      "010" when "011011010",
      "010" when "011011011",
      "010" when "011011100",
      "010" when "011011101",
      "010" when "011011110",
      "010" when "011011111",
      "010" when "011100000",
      "010" when "011100001",
      "010" when "011100010",
      "010" when "011100011",
      "010" when "011100100",
      "010" when "011100101",
      "010" when "011100110",
      "010" when "011100111",
      "010" when "011101000",
      "010" when "011101001",
      "010" when "011101010",
      "010" when "011101011",
      "010" when "011101100",
      "010" when "011101101",
      "010" when "011101110",
      "010" when "011101111",
      "010" when "011110000",
      "010" when "011110001",
      "010" when "011110010",
      "010" when "011110011",
      "010" when "011110100",
      "010" when "011110101",
      "010" when "011110110",
      "010" when "011110111",
      "010" when "011111000",
      "010" when "011111001",
      "010" when "011111010",
      "010" when "011111011",
      "010" when "011111100",
      "010" when "011111101",
      "010" when "011111110",
      "010" when "011111111",
      "110" when "100000000",
      "110" when "100000001",
      "110" when "100000010",
      "110" when "100000011",
      "110" when "100000100",
      "110" when "100000101",
      "110" when "100000110",
      "110" when "100000111",
      "110" when "100001000",
      "110" when "100001001",
      "110" when "100001010",
      "110" when "100001011",
      "110" when "100001100",
      "110" when "100001101",
      "110" when "100001110",
      "110" when "100001111",
      "110" when "100010000",
      "110" when "100010001",
      "110" when "100010010",
      "110" when "100010011",
      "110" when "100010100",
      "110" when "100010101",
      "110" when "100010110",
      "110" when "100010111",
      "110" when "100011000",
      "110" when "100011001",
      "110" when "100011010",
      "110" when "100011011",
      "110" when "100011100",
      "110" when "100011101",
      "110" when "100011110",
      "110" when "100011111",
      "110" when "100100000",
      "110" when "100100001",
      "110" when "100100010",
      "110" when "100100011",
      "110" when "100100100",
      "110" when "100100101",
      "110" when "100100110",
      "110" when "100100111",
      "110" when "100101000",
      "110" when "100101001",
      "110" when "100101010",
      "110" when "100101011",
      "110" when "100101100",
      "110" when "100101101",
      "110" when "100101110",
      "110" when "100101111",
      "110" when "100110000",
      "110" when "100110001",
      "110" when "100110010",
      "110" when "100110011",
      "110" when "100110100",
      "110" when "100110101",
      "110" when "100110110",
      "110" when "100110111",
      "110" when "100111000",
      "110" when "100111001",
      "110" when "100111010",
      "110" when "100111011",
      "110" when "100111100",
      "110" when "100111101",
      "110" when "100111110",
      "110" when "100111111",
      "110" when "101000000",
      "110" when "101000001",
      "110" when "101000010",
      "110" when "101000011",
      "110" when "101000100",
      "110" when "101000101",
      "110" when "101000110",
      "110" when "101000111",
      "110" when "101001000",
      "110" when "101001001",
      "110" when "101001010",
      "110" when "101001011",
      "110" when "101001100",
      "110" when "101001101",
      "110" when "101001110",
      "110" when "101001111",
      "110" when "101010000",
      "110" when "101010001",
      "110" when "101010010",
      "110" when "101010011",
      "110" when "101010100",
      "110" when "101010101",
      "110" when "101010110",
      "110" when "101010111",
      "110" when "101011000",
      "110" when "101011001",
      "110" when "101011010",
      "110" when "101011011",
      "110" when "101011100",
      "110" when "101011101",
      "110" when "101011110",
      "110" when "101011111",
      "110" when "101100000",
      "110" when "101100001",
      "110" when "101100010",
      "110" when "101100011",
      "110" when "101100100",
      "110" when "101100101",
      "110" when "101100110",
      "110" when "101100111",
      "110" when "101101000",
      "110" when "101101001",
      "110" when "101101010",
      "110" when "101101011",
      "110" when "101101100",
      "110" when "101101101",
      "110" when "101101110",
      "110" when "101101111",
      "110" when "101110000",
      "110" when "101110001",
      "110" when "101110010",
      "110" when "101110011",
      "110" when "101110100",
      "110" when "101110101",
      "110" when "101110110",
      "110" when "101110111",
      "110" when "101111000",
      "110" when "101111001",
      "110" when "101111010",
      "110" when "101111011",
      "110" when "101111100",
      "110" when "101111101",
      "110" when "101111110",
      "110" when "101111111",
      "110" when "110000000",
      "110" when "110000001",
      "110" when "110000010",
      "110" when "110000011",
      "110" when "110000100",
      "110" when "110000101",
      "110" when "110000110",
      "110" when "110000111",
      "110" when "110001000",
      "110" when "110001001",
      "110" when "110001010",
      "110" when "110001011",
      "110" when "110001100",
      "110" when "110001101",
      "110" when "110001110",
      "110" when "110001111",
      "110" when "110010000",
      "110" when "110010001",
      "110" when "110010010",
      "110" when "110010011",
      "110" when "110010100",
      "110" when "110010101",
      "110" when "110010110",
      "110" when "110010111",
      "110" when "110011000",
      "110" when "110011001",
      "110" when "110011010",
      "110" when "110011011",
      "110" when "110011100",
      "110" when "110011101",
      "110" when "110011110",
      "110" when "110011111",
      "110" when "110100000",
      "110" when "110100001",
      "110" when "110100010",
      "110" when "110100011",
      "110" when "110100100",
      "110" when "110100101",
      "110" when "110100110",
      "110" when "110100111",
      "110" when "110101000",
      "110" when "110101001",
      "110" when "110101010",
      "110" when "110101011",
      "110" when "110101100",
      "110" when "110101101",
      "110" when "110101110",
      "111" when "110101111",
      "110" when "110110000",
      "110" when "110110001",
      "110" when "110110010",
      "110" when "110110011",
      "110" when "110110100",
      "111" when "110110101",
      "111" when "110110110",
      "111" when "110110111",
      "110" when "110111000",
      "110" when "110111001",
      "110" when "110111010",
      "110" when "110111011",
      "111" when "110111100",
      "111" when "110111101",
      "111" when "110111110",
      "111" when "110111111",
      "110" when "111000000",
      "110" when "111000001",
      "111" when "111000010",
      "111" when "111000011",
      "111" when "111000100",
      "111" when "111000101",
      "111" when "111000110",
      "111" when "111000111",
      "110" when "111001000",
      "111" when "111001001",
      "111" when "111001010",
      "111" when "111001011",
      "111" when "111001100",
      "111" when "111001101",
      "111" when "111001110",
      "111" when "111001111",
      "111" when "111010000",
      "111" when "111010001",
      "111" when "111010010",
      "111" when "111010011",
      "111" when "111010100",
      "111" when "111010101",
      "111" when "111010110",
      "111" when "111010111",
      "111" when "111011000",
      "111" when "111011001",
      "111" when "111011010",
      "111" when "111011011",
      "111" when "111011100",
      "111" when "111011101",
      "111" when "111011110",
      "111" when "111011111",
      "111" when "111100000",
      "111" when "111100001",
      "111" when "111100010",
      "111" when "111100011",
      "111" when "111100100",
      "111" when "111100101",
      "111" when "111100110",
      "111" when "111100111",
      "111" when "111101000",
      "111" when "111101001",
      "111" when "111101010",
      "111" when "111101011",
      "000" when "111101100",
      "000" when "111101101",
      "000" when "111101110",
      "000" when "111101111",
      "000" when "111110000",
      "000" when "111110001",
      "000" when "111110010",
      "000" when "111110011",
      "000" when "111110100",
      "000" when "111110101",
      "000" when "111110110",
      "000" when "111110111",
      "000" when "111111000",
      "000" when "111111001",
      "000" when "111111010",
      "000" when "111111011",
      "000" when "111111100",
      "000" when "111111101",
      "000" when "111111110",
      "000" when "111111111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            FloatingPointDivider
--                         (FPDiv_8_23_Freq300_uid2)
-- VHDL generated for Kintex7 @ 300MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 9 cycles
-- Clock period (ns): 3.33333
-- Target frequency (MHz): 300
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointDivider_32_6_629333 is
    port (clk, ce_1, ce_2, ce_3, ce_4, ce_5, ce_6, ce_7, ce_8, ce_9 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointDivider_32_6_629333 is
   component selFunction_Freq300_uid4 is
      port ( X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal fX_c0 :  std_logic_vector(23 downto 0);
signal fY_c0 :  std_logic_vector(23 downto 0);
signal expR0_c0, expR0_c1, expR0_c2, expR0_c3, expR0_c4, expR0_c5, expR0_c6, expR0_c7, expR0_c8, expR0_c9 :  std_logic_vector(9 downto 0);
signal sR_c0, sR_c1, sR_c2, sR_c3, sR_c4, sR_c5, sR_c6, sR_c7, sR_c8, sR_c9 :  std_logic;
signal exnXY_c0 :  std_logic_vector(3 downto 0);
signal exnR0_c0, exnR0_c1, exnR0_c2, exnR0_c3, exnR0_c4, exnR0_c5, exnR0_c6, exnR0_c7, exnR0_c8, exnR0_c9 :  std_logic_vector(1 downto 0);
signal D_c0, D_c1, D_c2, D_c3, D_c4, D_c5, D_c6, D_c7 :  std_logic_vector(23 downto 0);
signal psX_c0 :  std_logic_vector(24 downto 0);
signal betaw14_c0 :  std_logic_vector(26 downto 0);
signal sel14_c0 :  std_logic_vector(8 downto 0);
signal q14_c0 :  std_logic_vector(2 downto 0);
signal q14_copy5_c0 :  std_logic_vector(2 downto 0);
signal absq14D_c0 :  std_logic_vector(26 downto 0);
signal w13_c0 :  std_logic_vector(26 downto 0);
signal betaw13_c0, betaw13_c1 :  std_logic_vector(26 downto 0);
signal sel13_c0 :  std_logic_vector(8 downto 0);
signal q13_c0, q13_c1 :  std_logic_vector(2 downto 0);
signal q13_copy6_c0 :  std_logic_vector(2 downto 0);
signal absq13D_c0, absq13D_c1 :  std_logic_vector(26 downto 0);
signal w12_c1 :  std_logic_vector(26 downto 0);
signal betaw12_c1 :  std_logic_vector(26 downto 0);
signal sel12_c1 :  std_logic_vector(8 downto 0);
signal q12_c1 :  std_logic_vector(2 downto 0);
signal q12_copy7_c1 :  std_logic_vector(2 downto 0);
signal absq12D_c1 :  std_logic_vector(26 downto 0);
signal w11_c1 :  std_logic_vector(26 downto 0);
signal betaw11_c1, betaw11_c2 :  std_logic_vector(26 downto 0);
signal sel11_c1 :  std_logic_vector(8 downto 0);
signal q11_c1, q11_c2 :  std_logic_vector(2 downto 0);
signal q11_copy8_c1 :  std_logic_vector(2 downto 0);
signal absq11D_c1, absq11D_c2 :  std_logic_vector(26 downto 0);
signal w10_c2 :  std_logic_vector(26 downto 0);
signal betaw10_c2 :  std_logic_vector(26 downto 0);
signal sel10_c2 :  std_logic_vector(8 downto 0);
signal q10_c2 :  std_logic_vector(2 downto 0);
signal q10_copy9_c2 :  std_logic_vector(2 downto 0);
signal absq10D_c2 :  std_logic_vector(26 downto 0);
signal w9_c2 :  std_logic_vector(26 downto 0);
signal betaw9_c2, betaw9_c3 :  std_logic_vector(26 downto 0);
signal sel9_c2 :  std_logic_vector(8 downto 0);
signal q9_c3 :  std_logic_vector(2 downto 0);
signal q9_copy10_c2, q9_copy10_c3 :  std_logic_vector(2 downto 0);
signal absq9D_c3 :  std_logic_vector(26 downto 0);
signal w8_c3 :  std_logic_vector(26 downto 0);
signal betaw8_c3, betaw8_c4 :  std_logic_vector(26 downto 0);
signal sel8_c3 :  std_logic_vector(8 downto 0);
signal q8_c3, q8_c4 :  std_logic_vector(2 downto 0);
signal q8_copy11_c3 :  std_logic_vector(2 downto 0);
signal absq8D_c3, absq8D_c4 :  std_logic_vector(26 downto 0);
signal w7_c4 :  std_logic_vector(26 downto 0);
signal betaw7_c4 :  std_logic_vector(26 downto 0);
signal sel7_c4 :  std_logic_vector(8 downto 0);
signal q7_c4 :  std_logic_vector(2 downto 0);
signal q7_copy12_c4 :  std_logic_vector(2 downto 0);
signal absq7D_c4 :  std_logic_vector(26 downto 0);
signal w6_c4 :  std_logic_vector(26 downto 0);
signal betaw6_c4, betaw6_c5 :  std_logic_vector(26 downto 0);
signal sel6_c4 :  std_logic_vector(8 downto 0);
signal q6_c4, q6_c5 :  std_logic_vector(2 downto 0);
signal q6_copy13_c4 :  std_logic_vector(2 downto 0);
signal absq6D_c4, absq6D_c5 :  std_logic_vector(26 downto 0);
signal w5_c5 :  std_logic_vector(26 downto 0);
signal betaw5_c5 :  std_logic_vector(26 downto 0);
signal sel5_c5 :  std_logic_vector(8 downto 0);
signal q5_c5 :  std_logic_vector(2 downto 0);
signal q5_copy14_c5 :  std_logic_vector(2 downto 0);
signal absq5D_c5 :  std_logic_vector(26 downto 0);
signal w4_c5 :  std_logic_vector(26 downto 0);
signal betaw4_c5, betaw4_c6 :  std_logic_vector(26 downto 0);
signal sel4_c5 :  std_logic_vector(8 downto 0);
signal q4_c6 :  std_logic_vector(2 downto 0);
signal q4_copy15_c5, q4_copy15_c6 :  std_logic_vector(2 downto 0);
signal absq4D_c6 :  std_logic_vector(26 downto 0);
signal w3_c6 :  std_logic_vector(26 downto 0);
signal betaw3_c6, betaw3_c7 :  std_logic_vector(26 downto 0);
signal sel3_c6 :  std_logic_vector(8 downto 0);
signal q3_c6, q3_c7 :  std_logic_vector(2 downto 0);
signal q3_copy16_c6 :  std_logic_vector(2 downto 0);
signal absq3D_c6, absq3D_c7 :  std_logic_vector(26 downto 0);
signal w2_c7 :  std_logic_vector(26 downto 0);
signal betaw2_c7 :  std_logic_vector(26 downto 0);
signal sel2_c7 :  std_logic_vector(8 downto 0);
signal q2_c7 :  std_logic_vector(2 downto 0);
signal q2_copy17_c7 :  std_logic_vector(2 downto 0);
signal absq2D_c7 :  std_logic_vector(26 downto 0);
signal w1_c7 :  std_logic_vector(26 downto 0);
signal betaw1_c7, betaw1_c8 :  std_logic_vector(26 downto 0);
signal sel1_c7 :  std_logic_vector(8 downto 0);
signal q1_c7, q1_c8 :  std_logic_vector(2 downto 0);
signal q1_copy18_c7 :  std_logic_vector(2 downto 0);
signal absq1D_c7, absq1D_c8 :  std_logic_vector(26 downto 0);
signal w0_c8 :  std_logic_vector(26 downto 0);
signal wfinal_c8 :  std_logic_vector(24 downto 0);
signal qM0_c8 :  std_logic;
signal qP14_c0, qP14_c1, qP14_c2, qP14_c3, qP14_c4, qP14_c5, qP14_c6, qP14_c7 :  std_logic_vector(1 downto 0);
signal qM14_c0, qM14_c1, qM14_c2, qM14_c3, qM14_c4, qM14_c5, qM14_c6, qM14_c7, qM14_c8 :  std_logic_vector(1 downto 0);
signal qP13_c0, qP13_c1, qP13_c2, qP13_c3, qP13_c4, qP13_c5, qP13_c6, qP13_c7 :  std_logic_vector(1 downto 0);
signal qM13_c0, qM13_c1, qM13_c2, qM13_c3, qM13_c4, qM13_c5, qM13_c6, qM13_c7, qM13_c8 :  std_logic_vector(1 downto 0);
signal qP12_c1, qP12_c2, qP12_c3, qP12_c4, qP12_c5, qP12_c6, qP12_c7 :  std_logic_vector(1 downto 0);
signal qM12_c1, qM12_c2, qM12_c3, qM12_c4, qM12_c5, qM12_c6, qM12_c7, qM12_c8 :  std_logic_vector(1 downto 0);
signal qP11_c1, qP11_c2, qP11_c3, qP11_c4, qP11_c5, qP11_c6, qP11_c7 :  std_logic_vector(1 downto 0);
signal qM11_c1, qM11_c2, qM11_c3, qM11_c4, qM11_c5, qM11_c6, qM11_c7, qM11_c8 :  std_logic_vector(1 downto 0);
signal qP10_c2, qP10_c3, qP10_c4, qP10_c5, qP10_c6, qP10_c7 :  std_logic_vector(1 downto 0);
signal qM10_c2, qM10_c3, qM10_c4, qM10_c5, qM10_c6, qM10_c7, qM10_c8 :  std_logic_vector(1 downto 0);
signal qP9_c3, qP9_c4, qP9_c5, qP9_c6, qP9_c7 :  std_logic_vector(1 downto 0);
signal qM9_c3, qM9_c4, qM9_c5, qM9_c6, qM9_c7, qM9_c8 :  std_logic_vector(1 downto 0);
signal qP8_c3, qP8_c4, qP8_c5, qP8_c6, qP8_c7 :  std_logic_vector(1 downto 0);
signal qM8_c3, qM8_c4, qM8_c5, qM8_c6, qM8_c7, qM8_c8 :  std_logic_vector(1 downto 0);
signal qP7_c4, qP7_c5, qP7_c6, qP7_c7 :  std_logic_vector(1 downto 0);
signal qM7_c4, qM7_c5, qM7_c6, qM7_c7, qM7_c8 :  std_logic_vector(1 downto 0);
signal qP6_c4, qP6_c5, qP6_c6, qP6_c7 :  std_logic_vector(1 downto 0);
signal qM6_c4, qM6_c5, qM6_c6, qM6_c7, qM6_c8 :  std_logic_vector(1 downto 0);
signal qP5_c5, qP5_c6, qP5_c7 :  std_logic_vector(1 downto 0);
signal qM5_c5, qM5_c6, qM5_c7, qM5_c8 :  std_logic_vector(1 downto 0);
signal qP4_c6, qP4_c7 :  std_logic_vector(1 downto 0);
signal qM4_c6, qM4_c7, qM4_c8 :  std_logic_vector(1 downto 0);
signal qP3_c6, qP3_c7 :  std_logic_vector(1 downto 0);
signal qM3_c6, qM3_c7, qM3_c8 :  std_logic_vector(1 downto 0);
signal qP2_c7 :  std_logic_vector(1 downto 0);
signal qM2_c7, qM2_c8 :  std_logic_vector(1 downto 0);
signal qP1_c7 :  std_logic_vector(1 downto 0);
signal qM1_c7, qM1_c8 :  std_logic_vector(1 downto 0);
signal qP_c7, qP_c8 :  std_logic_vector(27 downto 0);
signal qM_c8 :  std_logic_vector(27 downto 0);
signal quotient_c8 :  std_logic_vector(27 downto 0);
signal mR_c8, mR_c9 :  std_logic_vector(25 downto 0);
signal fRnorm_c8, fRnorm_c9 :  std_logic_vector(23 downto 0);
signal round_c8, round_c9 :  std_logic;
signal expR1_c9 :  std_logic_vector(9 downto 0);
signal expfrac_c9 :  std_logic_vector(32 downto 0);
signal expfracR_c9 :  std_logic_vector(32 downto 0);
signal exnR_c9 :  std_logic_vector(1 downto 0);
signal exnRfinal_c9 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               expR0_c1 <= expR0_c0;
               sR_c1 <= sR_c0;
               exnR0_c1 <= exnR0_c0;
               D_c1 <= D_c0;
               betaw13_c1 <= betaw13_c0;
               q13_c1 <= q13_c0;
               absq13D_c1 <= absq13D_c0;
               qP14_c1 <= qP14_c0;
               qM14_c1 <= qM14_c0;
               qP13_c1 <= qP13_c0;
               qM13_c1 <= qM13_c0;
            end if;
            if ce_2 = '1' then
               expR0_c2 <= expR0_c1;
               sR_c2 <= sR_c1;
               exnR0_c2 <= exnR0_c1;
               D_c2 <= D_c1;
               betaw11_c2 <= betaw11_c1;
               q11_c2 <= q11_c1;
               absq11D_c2 <= absq11D_c1;
               qP14_c2 <= qP14_c1;
               qM14_c2 <= qM14_c1;
               qP13_c2 <= qP13_c1;
               qM13_c2 <= qM13_c1;
               qP12_c2 <= qP12_c1;
               qM12_c2 <= qM12_c1;
               qP11_c2 <= qP11_c1;
               qM11_c2 <= qM11_c1;
            end if;
            if ce_3 = '1' then
               expR0_c3 <= expR0_c2;
               sR_c3 <= sR_c2;
               exnR0_c3 <= exnR0_c2;
               D_c3 <= D_c2;
               betaw9_c3 <= betaw9_c2;
               q9_copy10_c3 <= q9_copy10_c2;
               qP14_c3 <= qP14_c2;
               qM14_c3 <= qM14_c2;
               qP13_c3 <= qP13_c2;
               qM13_c3 <= qM13_c2;
               qP12_c3 <= qP12_c2;
               qM12_c3 <= qM12_c2;
               qP11_c3 <= qP11_c2;
               qM11_c3 <= qM11_c2;
               qP10_c3 <= qP10_c2;
               qM10_c3 <= qM10_c2;
            end if;
            if ce_4 = '1' then
               expR0_c4 <= expR0_c3;
               sR_c4 <= sR_c3;
               exnR0_c4 <= exnR0_c3;
               D_c4 <= D_c3;
               betaw8_c4 <= betaw8_c3;
               q8_c4 <= q8_c3;
               absq8D_c4 <= absq8D_c3;
               qP14_c4 <= qP14_c3;
               qM14_c4 <= qM14_c3;
               qP13_c4 <= qP13_c3;
               qM13_c4 <= qM13_c3;
               qP12_c4 <= qP12_c3;
               qM12_c4 <= qM12_c3;
               qP11_c4 <= qP11_c3;
               qM11_c4 <= qM11_c3;
               qP10_c4 <= qP10_c3;
               qM10_c4 <= qM10_c3;
               qP9_c4 <= qP9_c3;
               qM9_c4 <= qM9_c3;
               qP8_c4 <= qP8_c3;
               qM8_c4 <= qM8_c3;
            end if;
            if ce_5 = '1' then
               expR0_c5 <= expR0_c4;
               sR_c5 <= sR_c4;
               exnR0_c5 <= exnR0_c4;
               D_c5 <= D_c4;
               betaw6_c5 <= betaw6_c4;
               q6_c5 <= q6_c4;
               absq6D_c5 <= absq6D_c4;
               qP14_c5 <= qP14_c4;
               qM14_c5 <= qM14_c4;
               qP13_c5 <= qP13_c4;
               qM13_c5 <= qM13_c4;
               qP12_c5 <= qP12_c4;
               qM12_c5 <= qM12_c4;
               qP11_c5 <= qP11_c4;
               qM11_c5 <= qM11_c4;
               qP10_c5 <= qP10_c4;
               qM10_c5 <= qM10_c4;
               qP9_c5 <= qP9_c4;
               qM9_c5 <= qM9_c4;
               qP8_c5 <= qP8_c4;
               qM8_c5 <= qM8_c4;
               qP7_c5 <= qP7_c4;
               qM7_c5 <= qM7_c4;
               qP6_c5 <= qP6_c4;
               qM6_c5 <= qM6_c4;
            end if;
            if ce_6 = '1' then
               expR0_c6 <= expR0_c5;
               sR_c6 <= sR_c5;
               exnR0_c6 <= exnR0_c5;
               D_c6 <= D_c5;
               betaw4_c6 <= betaw4_c5;
               q4_copy15_c6 <= q4_copy15_c5;
               qP14_c6 <= qP14_c5;
               qM14_c6 <= qM14_c5;
               qP13_c6 <= qP13_c5;
               qM13_c6 <= qM13_c5;
               qP12_c6 <= qP12_c5;
               qM12_c6 <= qM12_c5;
               qP11_c6 <= qP11_c5;
               qM11_c6 <= qM11_c5;
               qP10_c6 <= qP10_c5;
               qM10_c6 <= qM10_c5;
               qP9_c6 <= qP9_c5;
               qM9_c6 <= qM9_c5;
               qP8_c6 <= qP8_c5;
               qM8_c6 <= qM8_c5;
               qP7_c6 <= qP7_c5;
               qM7_c6 <= qM7_c5;
               qP6_c6 <= qP6_c5;
               qM6_c6 <= qM6_c5;
               qP5_c6 <= qP5_c5;
               qM5_c6 <= qM5_c5;
            end if;
            if ce_7 = '1' then
               expR0_c7 <= expR0_c6;
               sR_c7 <= sR_c6;
               exnR0_c7 <= exnR0_c6;
               D_c7 <= D_c6;
               betaw3_c7 <= betaw3_c6;
               q3_c7 <= q3_c6;
               absq3D_c7 <= absq3D_c6;
               qP14_c7 <= qP14_c6;
               qM14_c7 <= qM14_c6;
               qP13_c7 <= qP13_c6;
               qM13_c7 <= qM13_c6;
               qP12_c7 <= qP12_c6;
               qM12_c7 <= qM12_c6;
               qP11_c7 <= qP11_c6;
               qM11_c7 <= qM11_c6;
               qP10_c7 <= qP10_c6;
               qM10_c7 <= qM10_c6;
               qP9_c7 <= qP9_c6;
               qM9_c7 <= qM9_c6;
               qP8_c7 <= qP8_c6;
               qM8_c7 <= qM8_c6;
               qP7_c7 <= qP7_c6;
               qM7_c7 <= qM7_c6;
               qP6_c7 <= qP6_c6;
               qM6_c7 <= qM6_c6;
               qP5_c7 <= qP5_c6;
               qM5_c7 <= qM5_c6;
               qP4_c7 <= qP4_c6;
               qM4_c7 <= qM4_c6;
               qP3_c7 <= qP3_c6;
               qM3_c7 <= qM3_c6;
            end if;
            if ce_8 = '1' then
               expR0_c8 <= expR0_c7;
               sR_c8 <= sR_c7;
               exnR0_c8 <= exnR0_c7;
               betaw1_c8 <= betaw1_c7;
               q1_c8 <= q1_c7;
               absq1D_c8 <= absq1D_c7;
               qM14_c8 <= qM14_c7;
               qM13_c8 <= qM13_c7;
               qM12_c8 <= qM12_c7;
               qM11_c8 <= qM11_c7;
               qM10_c8 <= qM10_c7;
               qM9_c8 <= qM9_c7;
               qM8_c8 <= qM8_c7;
               qM7_c8 <= qM7_c7;
               qM6_c8 <= qM6_c7;
               qM5_c8 <= qM5_c7;
               qM4_c8 <= qM4_c7;
               qM3_c8 <= qM3_c7;
               qM2_c8 <= qM2_c7;
               qM1_c8 <= qM1_c7;
               qP_c8 <= qP_c7;
            end if;
            if ce_9 = '1' then
               expR0_c9 <= expR0_c8;
               sR_c9 <= sR_c8;
               exnR0_c9 <= exnR0_c8;
               mR_c9 <= mR_c8;
               fRnorm_c9 <= fRnorm_c8;
               round_c9 <= round_c8;
            end if;
         end if;
      end process;
   fX_c0 <= "1" & X(22 downto 0);
   fY_c0 <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have fewer bits to pipeline
   expR0_c0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR_c0 <= X(31) xor Y(31);
   -- early exception handling 
   exnXY_c0 <= X(33 downto 32) & Y(33 downto 32);
   with exnXY_c0  select 
      exnR0_c0 <= 
         "01"	 when "0101",										-- normal
         "00"	 when "0001" | "0010" | "0110", -- zero
         "10"	 when "0100" | "1000" | "1001", -- overflow
         "11"	 when others;										-- NaN
   D_c0 <= fY_c0 ;
   psX_c0 <= "0" & fX_c0 ;
   betaw14_c0 <=  "00" & psX_c0;
   sel14_c0 <= betaw14_c0(26 downto 21) & D_c0(22 downto 20);
   SelFunctionTable14: selFunction_Freq300_uid4
      port map ( X => sel14_c0,
                 Y => q14_copy5_c0);
   q14_c0 <= q14_copy5_c0; -- output copy to hold a pipeline register if needed

   with q14_c0  select 
      absq14D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q14_c0(2)  select 
   w13_c0<= betaw14_c0 - absq14D_c0 when '0',
         betaw14_c0 + absq14D_c0 when others;

   betaw13_c0 <= w13_c0(24 downto 0) & "00"; -- multiplication by the radix
   sel13_c0 <= betaw13_c0(26 downto 21) & D_c0(22 downto 20);
   SelFunctionTable13: selFunction_Freq300_uid4
      port map ( X => sel13_c0,
                 Y => q13_copy6_c0);
   q13_c0 <= q13_copy6_c0; -- output copy to hold a pipeline register if needed

   with q13_c0  select 
      absq13D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q13_c1(2)  select 
   w12_c1<= betaw13_c1 - absq13D_c1 when '0',
         betaw13_c1 + absq13D_c1 when others;

   betaw12_c1 <= w12_c1(24 downto 0) & "00"; -- multiplication by the radix
   sel12_c1 <= betaw12_c1(26 downto 21) & D_c1(22 downto 20);
   SelFunctionTable12: selFunction_Freq300_uid4
      port map ( X => sel12_c1,
                 Y => q12_copy7_c1);
   q12_c1 <= q12_copy7_c1; -- output copy to hold a pipeline register if needed

   with q12_c1  select 
      absq12D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q12_c1(2)  select 
   w11_c1<= betaw12_c1 - absq12D_c1 when '0',
         betaw12_c1 + absq12D_c1 when others;

   betaw11_c1 <= w11_c1(24 downto 0) & "00"; -- multiplication by the radix
   sel11_c1 <= betaw11_c1(26 downto 21) & D_c1(22 downto 20);
   SelFunctionTable11: selFunction_Freq300_uid4
      port map ( X => sel11_c1,
                 Y => q11_copy8_c1);
   q11_c1 <= q11_copy8_c1; -- output copy to hold a pipeline register if needed

   with q11_c1  select 
      absq11D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q11_c2(2)  select 
   w10_c2<= betaw11_c2 - absq11D_c2 when '0',
         betaw11_c2 + absq11D_c2 when others;

   betaw10_c2 <= w10_c2(24 downto 0) & "00"; -- multiplication by the radix
   sel10_c2 <= betaw10_c2(26 downto 21) & D_c2(22 downto 20);
   SelFunctionTable10: selFunction_Freq300_uid4
      port map ( X => sel10_c2,
                 Y => q10_copy9_c2);
   q10_c2 <= q10_copy9_c2; -- output copy to hold a pipeline register if needed

   with q10_c2  select 
      absq10D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q10_c2(2)  select 
   w9_c2<= betaw10_c2 - absq10D_c2 when '0',
         betaw10_c2 + absq10D_c2 when others;

   betaw9_c2 <= w9_c2(24 downto 0) & "00"; -- multiplication by the radix
   sel9_c2 <= betaw9_c2(26 downto 21) & D_c2(22 downto 20);
   SelFunctionTable9: selFunction_Freq300_uid4
      port map ( X => sel9_c2,
                 Y => q9_copy10_c2);
   q9_c3 <= q9_copy10_c3; -- output copy to hold a pipeline register if needed

   with q9_c3  select 
      absq9D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q9_c3(2)  select 
   w8_c3<= betaw9_c3 - absq9D_c3 when '0',
         betaw9_c3 + absq9D_c3 when others;

   betaw8_c3 <= w8_c3(24 downto 0) & "00"; -- multiplication by the radix
   sel8_c3 <= betaw8_c3(26 downto 21) & D_c3(22 downto 20);
   SelFunctionTable8: selFunction_Freq300_uid4
      port map ( X => sel8_c3,
                 Y => q8_copy11_c3);
   q8_c3 <= q8_copy11_c3; -- output copy to hold a pipeline register if needed

   with q8_c3  select 
      absq8D_c3 <= 
         "000" & D_c3						 when "001" | "111", -- mult by 1
         "00" & D_c3 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q8_c4(2)  select 
   w7_c4<= betaw8_c4 - absq8D_c4 when '0',
         betaw8_c4 + absq8D_c4 when others;

   betaw7_c4 <= w7_c4(24 downto 0) & "00"; -- multiplication by the radix
   sel7_c4 <= betaw7_c4(26 downto 21) & D_c4(22 downto 20);
   SelFunctionTable7: selFunction_Freq300_uid4
      port map ( X => sel7_c4,
                 Y => q7_copy12_c4);
   q7_c4 <= q7_copy12_c4; -- output copy to hold a pipeline register if needed

   with q7_c4  select 
      absq7D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q7_c4(2)  select 
   w6_c4<= betaw7_c4 - absq7D_c4 when '0',
         betaw7_c4 + absq7D_c4 when others;

   betaw6_c4 <= w6_c4(24 downto 0) & "00"; -- multiplication by the radix
   sel6_c4 <= betaw6_c4(26 downto 21) & D_c4(22 downto 20);
   SelFunctionTable6: selFunction_Freq300_uid4
      port map ( X => sel6_c4,
                 Y => q6_copy13_c4);
   q6_c4 <= q6_copy13_c4; -- output copy to hold a pipeline register if needed

   with q6_c4  select 
      absq6D_c4 <= 
         "000" & D_c4						 when "001" | "111", -- mult by 1
         "00" & D_c4 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q6_c5(2)  select 
   w5_c5<= betaw6_c5 - absq6D_c5 when '0',
         betaw6_c5 + absq6D_c5 when others;

   betaw5_c5 <= w5_c5(24 downto 0) & "00"; -- multiplication by the radix
   sel5_c5 <= betaw5_c5(26 downto 21) & D_c5(22 downto 20);
   SelFunctionTable5: selFunction_Freq300_uid4
      port map ( X => sel5_c5,
                 Y => q5_copy14_c5);
   q5_c5 <= q5_copy14_c5; -- output copy to hold a pipeline register if needed

   with q5_c5  select 
      absq5D_c5 <= 
         "000" & D_c5						 when "001" | "111", -- mult by 1
         "00" & D_c5 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q5_c5(2)  select 
   w4_c5<= betaw5_c5 - absq5D_c5 when '0',
         betaw5_c5 + absq5D_c5 when others;

   betaw4_c5 <= w4_c5(24 downto 0) & "00"; -- multiplication by the radix
   sel4_c5 <= betaw4_c5(26 downto 21) & D_c5(22 downto 20);
   SelFunctionTable4: selFunction_Freq300_uid4
      port map ( X => sel4_c5,
                 Y => q4_copy15_c5);
   q4_c6 <= q4_copy15_c6; -- output copy to hold a pipeline register if needed

   with q4_c6  select 
      absq4D_c6 <= 
         "000" & D_c6						 when "001" | "111", -- mult by 1
         "00" & D_c6 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q4_c6(2)  select 
   w3_c6<= betaw4_c6 - absq4D_c6 when '0',
         betaw4_c6 + absq4D_c6 when others;

   betaw3_c6 <= w3_c6(24 downto 0) & "00"; -- multiplication by the radix
   sel3_c6 <= betaw3_c6(26 downto 21) & D_c6(22 downto 20);
   SelFunctionTable3: selFunction_Freq300_uid4
      port map ( X => sel3_c6,
                 Y => q3_copy16_c6);
   q3_c6 <= q3_copy16_c6; -- output copy to hold a pipeline register if needed

   with q3_c6  select 
      absq3D_c6 <= 
         "000" & D_c6						 when "001" | "111", -- mult by 1
         "00" & D_c6 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q3_c7(2)  select 
   w2_c7<= betaw3_c7 - absq3D_c7 when '0',
         betaw3_c7 + absq3D_c7 when others;

   betaw2_c7 <= w2_c7(24 downto 0) & "00"; -- multiplication by the radix
   sel2_c7 <= betaw2_c7(26 downto 21) & D_c7(22 downto 20);
   SelFunctionTable2: selFunction_Freq300_uid4
      port map ( X => sel2_c7,
                 Y => q2_copy17_c7);
   q2_c7 <= q2_copy17_c7; -- output copy to hold a pipeline register if needed

   with q2_c7  select 
      absq2D_c7 <= 
         "000" & D_c7						 when "001" | "111", -- mult by 1
         "00" & D_c7 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q2_c7(2)  select 
   w1_c7<= betaw2_c7 - absq2D_c7 when '0',
         betaw2_c7 + absq2D_c7 when others;

   betaw1_c7 <= w1_c7(24 downto 0) & "00"; -- multiplication by the radix
   sel1_c7 <= betaw1_c7(26 downto 21) & D_c7(22 downto 20);
   SelFunctionTable1: selFunction_Freq300_uid4
      port map ( X => sel1_c7,
                 Y => q1_copy18_c7);
   q1_c7 <= q1_copy18_c7; -- output copy to hold a pipeline register if needed

   with q1_c7  select 
      absq1D_c7 <= 
         "000" & D_c7						 when "001" | "111", -- mult by 1
         "00" & D_c7 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q1_c8(2)  select 
   w0_c8<= betaw1_c8 - absq1D_c8 when '0',
         betaw1_c8 + absq1D_c8 when others;

   wfinal_c8 <= w0_c8(24 downto 0);
   qM0_c8 <= wfinal_c8(24); -- rounding bit is the sign of the remainder
   qP14_c0 <=      q14_c0(1 downto 0);
   qM14_c0 <=      q14_c0(2) & "0";
   qP13_c0 <=      q13_c0(1 downto 0);
   qM13_c0 <=      q13_c0(2) & "0";
   qP12_c1 <=      q12_c1(1 downto 0);
   qM12_c1 <=      q12_c1(2) & "0";
   qP11_c1 <=      q11_c1(1 downto 0);
   qM11_c1 <=      q11_c1(2) & "0";
   qP10_c2 <=      q10_c2(1 downto 0);
   qM10_c2 <=      q10_c2(2) & "0";
   qP9_c3 <=      q9_c3(1 downto 0);
   qM9_c3 <=      q9_c3(2) & "0";
   qP8_c3 <=      q8_c3(1 downto 0);
   qM8_c3 <=      q8_c3(2) & "0";
   qP7_c4 <=      q7_c4(1 downto 0);
   qM7_c4 <=      q7_c4(2) & "0";
   qP6_c4 <=      q6_c4(1 downto 0);
   qM6_c4 <=      q6_c4(2) & "0";
   qP5_c5 <=      q5_c5(1 downto 0);
   qM5_c5 <=      q5_c5(2) & "0";
   qP4_c6 <=      q4_c6(1 downto 0);
   qM4_c6 <=      q4_c6(2) & "0";
   qP3_c6 <=      q3_c6(1 downto 0);
   qM3_c6 <=      q3_c6(2) & "0";
   qP2_c7 <=      q2_c7(1 downto 0);
   qM2_c7 <=      q2_c7(2) & "0";
   qP1_c7 <=      q1_c7(1 downto 0);
   qM1_c7 <=      q1_c7(2) & "0";
   qP_c7 <= qP14_c7 & qP13_c7 & qP12_c7 & qP11_c7 & qP10_c7 & qP9_c7 & qP8_c7 & qP7_c7 & qP6_c7 & qP5_c7 & qP4_c7 & qP3_c7 & qP2_c7 & qP1_c7;
   qM_c8 <= qM14_c8(0) & qM13_c8 & qM12_c8 & qM11_c8 & qM10_c8 & qM9_c8 & qM8_c8 & qM7_c8 & qM6_c8 & qM5_c8 & qM4_c8 & qM3_c8 & qM2_c8 & qM1_c8 & qM0_c8;
   quotient_c8 <= qP_c8 - qM_c8;
   -- We need a mR in (0, -wf-2) format: 1+wF fraction bits, 1 round bit, and 1 guard bit for the normalisation,
   -- quotient is the truncation of the exact quotient to at least 2^(-wF-2) bits
   -- now discarding its possible known MSB zeroes, and dropping the possible extra LSB bit (due to radix 4) 
   mR_c8 <= quotient_c8(26 downto 1); 
   -- normalisation
   fRnorm_c8 <=    mR_c8(24 downto 1)  when mR_c8(25)= '1'
           else mR_c8(23 downto 0);  -- now fRnorm is a (-1, -wF-1) fraction
   round_c8 <= fRnorm_c8(0); 
   expR1_c9 <= expR0_c9 + ("000" & (6 downto 1 => '1') & mR_c9(25)); -- add back bias
   -- final rounding
   expfrac_c9 <= expR1_c9 & fRnorm_c9(23 downto 1) ;
   expfracR_c9 <= expfrac_c9 + ((32 downto 1 => '0') & round_c9);
   exnR_c9 <=      "00"  when expfracR_c9(32) = '1'   -- underflow
           else "10"  when  expfracR_c9(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_c9  select 
      exnRfinal_c9 <= 
         exnR_c9   when "01", -- normal
         exnR0_c9  when others;
   R <= exnRfinal_c9 & sR_c9 & expfracR_c9(30 downto 0);
end architecture;




--------------------------------------------------------------------------------
--                          selFunction_Freq100_uid4
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X
-- Output signals: Y

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity selFunction_Freq100_uid4 is
    port (X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of selFunction_Freq100_uid4 is
signal Y0 :  std_logic_vector(2 downto 0);
attribute ram_extract: string;
attribute ram_style: string;
attribute ram_extract of Y0: signal is "yes";
attribute ram_style of Y0: signal is "distributed";
signal Y1 :  std_logic_vector(2 downto 0);
begin
   with X  select  Y0 <= 
      "000" when "000000000",
      "000" when "000000001",
      "000" when "000000010",
      "000" when "000000011",
      "000" when "000000100",
      "000" when "000000101",
      "000" when "000000110",
      "000" when "000000111",
      "000" when "000001000",
      "000" when "000001001",
      "000" when "000001010",
      "000" when "000001011",
      "000" when "000001100",
      "000" when "000001101",
      "000" when "000001110",
      "000" when "000001111",
      "001" when "000010000",
      "000" when "000010001",
      "000" when "000010010",
      "000" when "000010011",
      "000" when "000010100",
      "000" when "000010101",
      "000" when "000010110",
      "000" when "000010111",
      "001" when "000011000",
      "001" when "000011001",
      "001" when "000011010",
      "001" when "000011011",
      "000" when "000011100",
      "000" when "000011101",
      "000" when "000011110",
      "000" when "000011111",
      "001" when "000100000",
      "001" when "000100001",
      "001" when "000100010",
      "001" when "000100011",
      "001" when "000100100",
      "001" when "000100101",
      "001" when "000100110",
      "000" when "000100111",
      "001" when "000101000",
      "001" when "000101001",
      "001" when "000101010",
      "001" when "000101011",
      "001" when "000101100",
      "001" when "000101101",
      "001" when "000101110",
      "001" when "000101111",
      "010" when "000110000",
      "001" when "000110001",
      "001" when "000110010",
      "001" when "000110011",
      "001" when "000110100",
      "001" when "000110101",
      "001" when "000110110",
      "001" when "000110111",
      "010" when "000111000",
      "010" when "000111001",
      "001" when "000111010",
      "001" when "000111011",
      "001" when "000111100",
      "001" when "000111101",
      "001" when "000111110",
      "001" when "000111111",
      "010" when "001000000",
      "010" when "001000001",
      "010" when "001000010",
      "001" when "001000011",
      "001" when "001000100",
      "001" when "001000101",
      "001" when "001000110",
      "001" when "001000111",
      "010" when "001001000",
      "010" when "001001001",
      "010" when "001001010",
      "010" when "001001011",
      "001" when "001001100",
      "001" when "001001101",
      "001" when "001001110",
      "001" when "001001111",
      "010" when "001010000",
      "010" when "001010001",
      "010" when "001010010",
      "010" when "001010011",
      "010" when "001010100",
      "010" when "001010101",
      "001" when "001010110",
      "001" when "001010111",
      "010" when "001011000",
      "010" when "001011001",
      "010" when "001011010",
      "010" when "001011011",
      "010" when "001011100",
      "010" when "001011101",
      "010" when "001011110",
      "001" when "001011111",
      "010" when "001100000",
      "010" when "001100001",
      "010" when "001100010",
      "010" when "001100011",
      "010" when "001100100",
      "010" when "001100101",
      "010" when "001100110",
      "010" when "001100111",
      "010" when "001101000",
      "010" when "001101001",
      "010" when "001101010",
      "010" when "001101011",
      "010" when "001101100",
      "010" when "001101101",
      "010" when "001101110",
      "010" when "001101111",
      "010" when "001110000",
      "010" when "001110001",
      "010" when "001110010",
      "010" when "001110011",
      "010" when "001110100",
      "010" when "001110101",
      "010" when "001110110",
      "010" when "001110111",
      "010" when "001111000",
      "010" when "001111001",
      "010" when "001111010",
      "010" when "001111011",
      "010" when "001111100",
      "010" when "001111101",
      "010" when "001111110",
      "010" when "001111111",
      "010" when "010000000",
      "010" when "010000001",
      "010" when "010000010",
      "010" when "010000011",
      "010" when "010000100",
      "010" when "010000101",
      "010" when "010000110",
      "010" when "010000111",
      "010" when "010001000",
      "010" when "010001001",
      "010" when "010001010",
      "010" when "010001011",
      "010" when "010001100",
      "010" when "010001101",
      "010" when "010001110",
      "010" when "010001111",
      "010" when "010010000",
      "010" when "010010001",
      "010" when "010010010",
      "010" when "010010011",
      "010" when "010010100",
      "010" when "010010101",
      "010" when "010010110",
      "010" when "010010111",
      "010" when "010011000",
      "010" when "010011001",
      "010" when "010011010",
      "010" when "010011011",
      "010" when "010011100",
      "010" when "010011101",
      "010" when "010011110",
      "010" when "010011111",
      "010" when "010100000",
      "010" when "010100001",
      "010" when "010100010",
      "010" when "010100011",
      "010" when "010100100",
      "010" when "010100101",
      "010" when "010100110",
      "010" when "010100111",
      "010" when "010101000",
      "010" when "010101001",
      "010" when "010101010",
      "010" when "010101011",
      "010" when "010101100",
      "010" when "010101101",
      "010" when "010101110",
      "010" when "010101111",
      "010" when "010110000",
      "010" when "010110001",
      "010" when "010110010",
      "010" when "010110011",
      "010" when "010110100",
      "010" when "010110101",
      "010" when "010110110",
      "010" when "010110111",
      "010" when "010111000",
      "010" when "010111001",
      "010" when "010111010",
      "010" when "010111011",
      "010" when "010111100",
      "010" when "010111101",
      "010" when "010111110",
      "010" when "010111111",
      "010" when "011000000",
      "010" when "011000001",
      "010" when "011000010",
      "010" when "011000011",
      "010" when "011000100",
      "010" when "011000101",
      "010" when "011000110",
      "010" when "011000111",
      "010" when "011001000",
      "010" when "011001001",
      "010" when "011001010",
      "010" when "011001011",
      "010" when "011001100",
      "010" when "011001101",
      "010" when "011001110",
      "010" when "011001111",
      "010" when "011010000",
      "010" when "011010001",
      "010" when "011010010",
      "010" when "011010011",
      "010" when "011010100",
      "010" when "011010101",
      "010" when "011010110",
      "010" when "011010111",
      "010" when "011011000",
      "010" when "011011001",
      "010" when "011011010",
      "010" when "011011011",
      "010" when "011011100",
      "010" when "011011101",
      "010" when "011011110",
      "010" when "011011111",
      "010" when "011100000",
      "010" when "011100001",
      "010" when "011100010",
      "010" when "011100011",
      "010" when "011100100",
      "010" when "011100101",
      "010" when "011100110",
      "010" when "011100111",
      "010" when "011101000",
      "010" when "011101001",
      "010" when "011101010",
      "010" when "011101011",
      "010" when "011101100",
      "010" when "011101101",
      "010" when "011101110",
      "010" when "011101111",
      "010" when "011110000",
      "010" when "011110001",
      "010" when "011110010",
      "010" when "011110011",
      "010" when "011110100",
      "010" when "011110101",
      "010" when "011110110",
      "010" when "011110111",
      "010" when "011111000",
      "010" when "011111001",
      "010" when "011111010",
      "010" when "011111011",
      "010" when "011111100",
      "010" when "011111101",
      "010" when "011111110",
      "010" when "011111111",
      "110" when "100000000",
      "110" when "100000001",
      "110" when "100000010",
      "110" when "100000011",
      "110" when "100000100",
      "110" when "100000101",
      "110" when "100000110",
      "110" when "100000111",
      "110" when "100001000",
      "110" when "100001001",
      "110" when "100001010",
      "110" when "100001011",
      "110" when "100001100",
      "110" when "100001101",
      "110" when "100001110",
      "110" when "100001111",
      "110" when "100010000",
      "110" when "100010001",
      "110" when "100010010",
      "110" when "100010011",
      "110" when "100010100",
      "110" when "100010101",
      "110" when "100010110",
      "110" when "100010111",
      "110" when "100011000",
      "110" when "100011001",
      "110" when "100011010",
      "110" when "100011011",
      "110" when "100011100",
      "110" when "100011101",
      "110" when "100011110",
      "110" when "100011111",
      "110" when "100100000",
      "110" when "100100001",
      "110" when "100100010",
      "110" when "100100011",
      "110" when "100100100",
      "110" when "100100101",
      "110" when "100100110",
      "110" when "100100111",
      "110" when "100101000",
      "110" when "100101001",
      "110" when "100101010",
      "110" when "100101011",
      "110" when "100101100",
      "110" when "100101101",
      "110" when "100101110",
      "110" when "100101111",
      "110" when "100110000",
      "110" when "100110001",
      "110" when "100110010",
      "110" when "100110011",
      "110" when "100110100",
      "110" when "100110101",
      "110" when "100110110",
      "110" when "100110111",
      "110" when "100111000",
      "110" when "100111001",
      "110" when "100111010",
      "110" when "100111011",
      "110" when "100111100",
      "110" when "100111101",
      "110" when "100111110",
      "110" when "100111111",
      "110" when "101000000",
      "110" when "101000001",
      "110" when "101000010",
      "110" when "101000011",
      "110" when "101000100",
      "110" when "101000101",
      "110" when "101000110",
      "110" when "101000111",
      "110" when "101001000",
      "110" when "101001001",
      "110" when "101001010",
      "110" when "101001011",
      "110" when "101001100",
      "110" when "101001101",
      "110" when "101001110",
      "110" when "101001111",
      "110" when "101010000",
      "110" when "101010001",
      "110" when "101010010",
      "110" when "101010011",
      "110" when "101010100",
      "110" when "101010101",
      "110" when "101010110",
      "110" when "101010111",
      "110" when "101011000",
      "110" when "101011001",
      "110" when "101011010",
      "110" when "101011011",
      "110" when "101011100",
      "110" when "101011101",
      "110" when "101011110",
      "110" when "101011111",
      "110" when "101100000",
      "110" when "101100001",
      "110" when "101100010",
      "110" when "101100011",
      "110" when "101100100",
      "110" when "101100101",
      "110" when "101100110",
      "110" when "101100111",
      "110" when "101101000",
      "110" when "101101001",
      "110" when "101101010",
      "110" when "101101011",
      "110" when "101101100",
      "110" when "101101101",
      "110" when "101101110",
      "110" when "101101111",
      "110" when "101110000",
      "110" when "101110001",
      "110" when "101110010",
      "110" when "101110011",
      "110" when "101110100",
      "110" when "101110101",
      "110" when "101110110",
      "110" when "101110111",
      "110" when "101111000",
      "110" when "101111001",
      "110" when "101111010",
      "110" when "101111011",
      "110" when "101111100",
      "110" when "101111101",
      "110" when "101111110",
      "110" when "101111111",
      "110" when "110000000",
      "110" when "110000001",
      "110" when "110000010",
      "110" when "110000011",
      "110" when "110000100",
      "110" when "110000101",
      "110" when "110000110",
      "110" when "110000111",
      "110" when "110001000",
      "110" when "110001001",
      "110" when "110001010",
      "110" when "110001011",
      "110" when "110001100",
      "110" when "110001101",
      "110" when "110001110",
      "110" when "110001111",
      "110" when "110010000",
      "110" when "110010001",
      "110" when "110010010",
      "110" when "110010011",
      "110" when "110010100",
      "110" when "110010101",
      "110" when "110010110",
      "110" when "110010111",
      "110" when "110011000",
      "110" when "110011001",
      "110" when "110011010",
      "110" when "110011011",
      "110" when "110011100",
      "110" when "110011101",
      "110" when "110011110",
      "110" when "110011111",
      "110" when "110100000",
      "110" when "110100001",
      "110" when "110100010",
      "110" when "110100011",
      "110" when "110100100",
      "110" when "110100101",
      "110" when "110100110",
      "110" when "110100111",
      "110" when "110101000",
      "110" when "110101001",
      "110" when "110101010",
      "110" when "110101011",
      "110" when "110101100",
      "110" when "110101101",
      "110" when "110101110",
      "111" when "110101111",
      "110" when "110110000",
      "110" when "110110001",
      "110" when "110110010",
      "110" when "110110011",
      "110" when "110110100",
      "111" when "110110101",
      "111" when "110110110",
      "111" when "110110111",
      "110" when "110111000",
      "110" when "110111001",
      "110" when "110111010",
      "110" when "110111011",
      "111" when "110111100",
      "111" when "110111101",
      "111" when "110111110",
      "111" when "110111111",
      "110" when "111000000",
      "110" when "111000001",
      "111" when "111000010",
      "111" when "111000011",
      "111" when "111000100",
      "111" when "111000101",
      "111" when "111000110",
      "111" when "111000111",
      "110" when "111001000",
      "111" when "111001001",
      "111" when "111001010",
      "111" when "111001011",
      "111" when "111001100",
      "111" when "111001101",
      "111" when "111001110",
      "111" when "111001111",
      "111" when "111010000",
      "111" when "111010001",
      "111" when "111010010",
      "111" when "111010011",
      "111" when "111010100",
      "111" when "111010101",
      "111" when "111010110",
      "111" when "111010111",
      "111" when "111011000",
      "111" when "111011001",
      "111" when "111011010",
      "111" when "111011011",
      "111" when "111011100",
      "111" when "111011101",
      "111" when "111011110",
      "111" when "111011111",
      "111" when "111100000",
      "111" when "111100001",
      "111" when "111100010",
      "111" when "111100011",
      "111" when "111100100",
      "111" when "111100101",
      "111" when "111100110",
      "111" when "111100111",
      "111" when "111101000",
      "111" when "111101001",
      "111" when "111101010",
      "111" when "111101011",
      "000" when "111101100",
      "000" when "111101101",
      "000" when "111101110",
      "000" when "111101111",
      "000" when "111110000",
      "000" when "111110001",
      "000" when "111110010",
      "000" when "111110011",
      "000" when "111110100",
      "000" when "111110101",
      "000" when "111110110",
      "000" when "111110111",
      "000" when "111111000",
      "000" when "111111001",
      "000" when "111111010",
      "000" when "111111011",
      "000" when "111111100",
      "000" when "111111101",
      "000" when "111111110",
      "000" when "111111111",
      "---" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                            FloatingPointDivider
--                         (FPDiv_8_23_Freq100_uid2)
-- VHDL generated for Kintex7 @ 100MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Maxime Christ, Florent de Dinechin (2015)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 10
-- Target frequency (MHz): 100
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FloatingPointDivider_32_14_152000 is
    port (clk, ce_1, ce_2 : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0)   );
end entity;

architecture arch of FloatingPointDivider_32_14_152000 is
   component selFunction_Freq100_uid4 is
      port ( X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(2 downto 0)   );
   end component;

signal fX_c0 :  std_logic_vector(23 downto 0);
signal fY_c0 :  std_logic_vector(23 downto 0);
signal expR0_c0, expR0_c1, expR0_c2 :  std_logic_vector(9 downto 0);
signal sR_c0, sR_c1, sR_c2 :  std_logic;
signal exnXY_c0 :  std_logic_vector(3 downto 0);
signal exnR0_c0, exnR0_c1, exnR0_c2 :  std_logic_vector(1 downto 0);
signal D_c0, D_c1, D_c2 :  std_logic_vector(23 downto 0);
signal psX_c0 :  std_logic_vector(24 downto 0);
signal betaw14_c0 :  std_logic_vector(26 downto 0);
signal sel14_c0 :  std_logic_vector(8 downto 0);
signal q14_c0 :  std_logic_vector(2 downto 0);
signal q14_copy5_c0 :  std_logic_vector(2 downto 0);
signal absq14D_c0 :  std_logic_vector(26 downto 0);
signal w13_c0 :  std_logic_vector(26 downto 0);
signal betaw13_c0 :  std_logic_vector(26 downto 0);
signal sel13_c0 :  std_logic_vector(8 downto 0);
signal q13_c0 :  std_logic_vector(2 downto 0);
signal q13_copy6_c0 :  std_logic_vector(2 downto 0);
signal absq13D_c0 :  std_logic_vector(26 downto 0);
signal w12_c0 :  std_logic_vector(26 downto 0);
signal betaw12_c0 :  std_logic_vector(26 downto 0);
signal sel12_c0 :  std_logic_vector(8 downto 0);
signal q12_c0 :  std_logic_vector(2 downto 0);
signal q12_copy7_c0 :  std_logic_vector(2 downto 0);
signal absq12D_c0 :  std_logic_vector(26 downto 0);
signal w11_c0 :  std_logic_vector(26 downto 0);
signal betaw11_c0 :  std_logic_vector(26 downto 0);
signal sel11_c0 :  std_logic_vector(8 downto 0);
signal q11_c0 :  std_logic_vector(2 downto 0);
signal q11_copy8_c0 :  std_logic_vector(2 downto 0);
signal absq11D_c0 :  std_logic_vector(26 downto 0);
signal w10_c0 :  std_logic_vector(26 downto 0);
signal betaw10_c0 :  std_logic_vector(26 downto 0);
signal sel10_c0 :  std_logic_vector(8 downto 0);
signal q10_c0 :  std_logic_vector(2 downto 0);
signal q10_copy9_c0 :  std_logic_vector(2 downto 0);
signal absq10D_c0 :  std_logic_vector(26 downto 0);
signal w9_c0 :  std_logic_vector(26 downto 0);
signal betaw9_c0, betaw9_c1 :  std_logic_vector(26 downto 0);
signal sel9_c0 :  std_logic_vector(8 downto 0);
signal q9_c0, q9_c1 :  std_logic_vector(2 downto 0);
signal q9_copy10_c0 :  std_logic_vector(2 downto 0);
signal absq9D_c0, absq9D_c1 :  std_logic_vector(26 downto 0);
signal w8_c1 :  std_logic_vector(26 downto 0);
signal betaw8_c1 :  std_logic_vector(26 downto 0);
signal sel8_c1 :  std_logic_vector(8 downto 0);
signal q8_c1 :  std_logic_vector(2 downto 0);
signal q8_copy11_c1 :  std_logic_vector(2 downto 0);
signal absq8D_c1 :  std_logic_vector(26 downto 0);
signal w7_c1 :  std_logic_vector(26 downto 0);
signal betaw7_c1 :  std_logic_vector(26 downto 0);
signal sel7_c1 :  std_logic_vector(8 downto 0);
signal q7_c1 :  std_logic_vector(2 downto 0);
signal q7_copy12_c1 :  std_logic_vector(2 downto 0);
signal absq7D_c1 :  std_logic_vector(26 downto 0);
signal w6_c1 :  std_logic_vector(26 downto 0);
signal betaw6_c1 :  std_logic_vector(26 downto 0);
signal sel6_c1 :  std_logic_vector(8 downto 0);
signal q6_c1 :  std_logic_vector(2 downto 0);
signal q6_copy13_c1 :  std_logic_vector(2 downto 0);
signal absq6D_c1 :  std_logic_vector(26 downto 0);
signal w5_c1 :  std_logic_vector(26 downto 0);
signal betaw5_c1 :  std_logic_vector(26 downto 0);
signal sel5_c1 :  std_logic_vector(8 downto 0);
signal q5_c1 :  std_logic_vector(2 downto 0);
signal q5_copy14_c1 :  std_logic_vector(2 downto 0);
signal absq5D_c1 :  std_logic_vector(26 downto 0);
signal w4_c1 :  std_logic_vector(26 downto 0);
signal betaw4_c1, betaw4_c2 :  std_logic_vector(26 downto 0);
signal sel4_c1 :  std_logic_vector(8 downto 0);
signal q4_c1, q4_c2 :  std_logic_vector(2 downto 0);
signal q4_copy15_c1 :  std_logic_vector(2 downto 0);
signal absq4D_c1, absq4D_c2 :  std_logic_vector(26 downto 0);
signal w3_c2 :  std_logic_vector(26 downto 0);
signal betaw3_c2 :  std_logic_vector(26 downto 0);
signal sel3_c2 :  std_logic_vector(8 downto 0);
signal q3_c2 :  std_logic_vector(2 downto 0);
signal q3_copy16_c2 :  std_logic_vector(2 downto 0);
signal absq3D_c2 :  std_logic_vector(26 downto 0);
signal w2_c2 :  std_logic_vector(26 downto 0);
signal betaw2_c2 :  std_logic_vector(26 downto 0);
signal sel2_c2 :  std_logic_vector(8 downto 0);
signal q2_c2 :  std_logic_vector(2 downto 0);
signal q2_copy17_c2 :  std_logic_vector(2 downto 0);
signal absq2D_c2 :  std_logic_vector(26 downto 0);
signal w1_c2 :  std_logic_vector(26 downto 0);
signal betaw1_c2 :  std_logic_vector(26 downto 0);
signal sel1_c2 :  std_logic_vector(8 downto 0);
signal q1_c2 :  std_logic_vector(2 downto 0);
signal q1_copy18_c2 :  std_logic_vector(2 downto 0);
signal absq1D_c2 :  std_logic_vector(26 downto 0);
signal w0_c2 :  std_logic_vector(26 downto 0);
signal wfinal_c2 :  std_logic_vector(24 downto 0);
signal qM0_c2 :  std_logic;
signal qP14_c0, qP14_c1, qP14_c2 :  std_logic_vector(1 downto 0);
signal qM14_c0, qM14_c1, qM14_c2 :  std_logic_vector(1 downto 0);
signal qP13_c0, qP13_c1, qP13_c2 :  std_logic_vector(1 downto 0);
signal qM13_c0, qM13_c1, qM13_c2 :  std_logic_vector(1 downto 0);
signal qP12_c0, qP12_c1, qP12_c2 :  std_logic_vector(1 downto 0);
signal qM12_c0, qM12_c1, qM12_c2 :  std_logic_vector(1 downto 0);
signal qP11_c0, qP11_c1, qP11_c2 :  std_logic_vector(1 downto 0);
signal qM11_c0, qM11_c1, qM11_c2 :  std_logic_vector(1 downto 0);
signal qP10_c0, qP10_c1, qP10_c2 :  std_logic_vector(1 downto 0);
signal qM10_c0, qM10_c1, qM10_c2 :  std_logic_vector(1 downto 0);
signal qP9_c0, qP9_c1, qP9_c2 :  std_logic_vector(1 downto 0);
signal qM9_c0, qM9_c1, qM9_c2 :  std_logic_vector(1 downto 0);
signal qP8_c1, qP8_c2 :  std_logic_vector(1 downto 0);
signal qM8_c1, qM8_c2 :  std_logic_vector(1 downto 0);
signal qP7_c1, qP7_c2 :  std_logic_vector(1 downto 0);
signal qM7_c1, qM7_c2 :  std_logic_vector(1 downto 0);
signal qP6_c1, qP6_c2 :  std_logic_vector(1 downto 0);
signal qM6_c1, qM6_c2 :  std_logic_vector(1 downto 0);
signal qP5_c1, qP5_c2 :  std_logic_vector(1 downto 0);
signal qM5_c1, qM5_c2 :  std_logic_vector(1 downto 0);
signal qP4_c1, qP4_c2 :  std_logic_vector(1 downto 0);
signal qM4_c1, qM4_c2 :  std_logic_vector(1 downto 0);
signal qP3_c2 :  std_logic_vector(1 downto 0);
signal qM3_c2 :  std_logic_vector(1 downto 0);
signal qP2_c2 :  std_logic_vector(1 downto 0);
signal qM2_c2 :  std_logic_vector(1 downto 0);
signal qP1_c2 :  std_logic_vector(1 downto 0);
signal qM1_c2 :  std_logic_vector(1 downto 0);
signal qP_c2 :  std_logic_vector(27 downto 0);
signal qM_c2 :  std_logic_vector(27 downto 0);
signal quotient_c2 :  std_logic_vector(27 downto 0);
signal mR_c2 :  std_logic_vector(25 downto 0);
signal fRnorm_c2 :  std_logic_vector(23 downto 0);
signal round_c2 :  std_logic;
signal expR1_c2 :  std_logic_vector(9 downto 0);
signal expfrac_c2 :  std_logic_vector(32 downto 0);
signal expfracR_c2 :  std_logic_vector(32 downto 0);
signal exnR_c2 :  std_logic_vector(1 downto 0);
signal exnRfinal_c2 :  std_logic_vector(1 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            if ce_1 = '1' then
               expR0_c1 <= expR0_c0;
               sR_c1 <= sR_c0;
               exnR0_c1 <= exnR0_c0;
               D_c1 <= D_c0;
               betaw9_c1 <= betaw9_c0;
               q9_c1 <= q9_c0;
               absq9D_c1 <= absq9D_c0;
               qP14_c1 <= qP14_c0;
               qM14_c1 <= qM14_c0;
               qP13_c1 <= qP13_c0;
               qM13_c1 <= qM13_c0;
               qP12_c1 <= qP12_c0;
               qM12_c1 <= qM12_c0;
               qP11_c1 <= qP11_c0;
               qM11_c1 <= qM11_c0;
               qP10_c1 <= qP10_c0;
               qM10_c1 <= qM10_c0;
               qP9_c1 <= qP9_c0;
               qM9_c1 <= qM9_c0;
            end if;
            if ce_2 = '1' then
               expR0_c2 <= expR0_c1;
               sR_c2 <= sR_c1;
               exnR0_c2 <= exnR0_c1;
               D_c2 <= D_c1;
               betaw4_c2 <= betaw4_c1;
               q4_c2 <= q4_c1;
               absq4D_c2 <= absq4D_c1;
               qP14_c2 <= qP14_c1;
               qM14_c2 <= qM14_c1;
               qP13_c2 <= qP13_c1;
               qM13_c2 <= qM13_c1;
               qP12_c2 <= qP12_c1;
               qM12_c2 <= qM12_c1;
               qP11_c2 <= qP11_c1;
               qM11_c2 <= qM11_c1;
               qP10_c2 <= qP10_c1;
               qM10_c2 <= qM10_c1;
               qP9_c2 <= qP9_c1;
               qM9_c2 <= qM9_c1;
               qP8_c2 <= qP8_c1;
               qM8_c2 <= qM8_c1;
               qP7_c2 <= qP7_c1;
               qM7_c2 <= qM7_c1;
               qP6_c2 <= qP6_c1;
               qM6_c2 <= qM6_c1;
               qP5_c2 <= qP5_c1;
               qM5_c2 <= qM5_c1;
               qP4_c2 <= qP4_c1;
               qM4_c2 <= qM4_c1;
            end if;
         end if;
      end process;
   fX_c0 <= "1" & X(22 downto 0);
   fY_c0 <= "1" & Y(22 downto 0);
   -- exponent difference, sign and exception combination computed early, to have fewer bits to pipeline
   expR0_c0 <= ("00" & X(30 downto 23)) - ("00" & Y(30 downto 23));
   sR_c0 <= X(31) xor Y(31);
   -- early exception handling 
   exnXY_c0 <= X(33 downto 32) & Y(33 downto 32);
   with exnXY_c0  select 
      exnR0_c0 <= 
         "01"	 when "0101",										-- normal
         "00"	 when "0001" | "0010" | "0110", -- zero
         "10"	 when "0100" | "1000" | "1001", -- overflow
         "11"	 when others;										-- NaN
   D_c0 <= fY_c0 ;
   psX_c0 <= "0" & fX_c0 ;
   betaw14_c0 <=  "00" & psX_c0;
   sel14_c0 <= betaw14_c0(26 downto 21) & D_c0(22 downto 20);
   SelFunctionTable14: selFunction_Freq100_uid4
      port map ( X => sel14_c0,
                 Y => q14_copy5_c0);
   q14_c0 <= q14_copy5_c0; -- output copy to hold a pipeline register if needed

   with q14_c0  select 
      absq14D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q14_c0(2)  select 
   w13_c0<= betaw14_c0 - absq14D_c0 when '0',
         betaw14_c0 + absq14D_c0 when others;

   betaw13_c0 <= w13_c0(24 downto 0) & "00"; -- multiplication by the radix
   sel13_c0 <= betaw13_c0(26 downto 21) & D_c0(22 downto 20);
   SelFunctionTable13: selFunction_Freq100_uid4
      port map ( X => sel13_c0,
                 Y => q13_copy6_c0);
   q13_c0 <= q13_copy6_c0; -- output copy to hold a pipeline register if needed

   with q13_c0  select 
      absq13D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q13_c0(2)  select 
   w12_c0<= betaw13_c0 - absq13D_c0 when '0',
         betaw13_c0 + absq13D_c0 when others;

   betaw12_c0 <= w12_c0(24 downto 0) & "00"; -- multiplication by the radix
   sel12_c0 <= betaw12_c0(26 downto 21) & D_c0(22 downto 20);
   SelFunctionTable12: selFunction_Freq100_uid4
      port map ( X => sel12_c0,
                 Y => q12_copy7_c0);
   q12_c0 <= q12_copy7_c0; -- output copy to hold a pipeline register if needed

   with q12_c0  select 
      absq12D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q12_c0(2)  select 
   w11_c0<= betaw12_c0 - absq12D_c0 when '0',
         betaw12_c0 + absq12D_c0 when others;

   betaw11_c0 <= w11_c0(24 downto 0) & "00"; -- multiplication by the radix
   sel11_c0 <= betaw11_c0(26 downto 21) & D_c0(22 downto 20);
   SelFunctionTable11: selFunction_Freq100_uid4
      port map ( X => sel11_c0,
                 Y => q11_copy8_c0);
   q11_c0 <= q11_copy8_c0; -- output copy to hold a pipeline register if needed

   with q11_c0  select 
      absq11D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q11_c0(2)  select 
   w10_c0<= betaw11_c0 - absq11D_c0 when '0',
         betaw11_c0 + absq11D_c0 when others;

   betaw10_c0 <= w10_c0(24 downto 0) & "00"; -- multiplication by the radix
   sel10_c0 <= betaw10_c0(26 downto 21) & D_c0(22 downto 20);
   SelFunctionTable10: selFunction_Freq100_uid4
      port map ( X => sel10_c0,
                 Y => q10_copy9_c0);
   q10_c0 <= q10_copy9_c0; -- output copy to hold a pipeline register if needed

   with q10_c0  select 
      absq10D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q10_c0(2)  select 
   w9_c0<= betaw10_c0 - absq10D_c0 when '0',
         betaw10_c0 + absq10D_c0 when others;

   betaw9_c0 <= w9_c0(24 downto 0) & "00"; -- multiplication by the radix
   sel9_c0 <= betaw9_c0(26 downto 21) & D_c0(22 downto 20);
   SelFunctionTable9: selFunction_Freq100_uid4
      port map ( X => sel9_c0,
                 Y => q9_copy10_c0);
   q9_c0 <= q9_copy10_c0; -- output copy to hold a pipeline register if needed

   with q9_c0  select 
      absq9D_c0 <= 
         "000" & D_c0						 when "001" | "111", -- mult by 1
         "00" & D_c0 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q9_c1(2)  select 
   w8_c1<= betaw9_c1 - absq9D_c1 when '0',
         betaw9_c1 + absq9D_c1 when others;

   betaw8_c1 <= w8_c1(24 downto 0) & "00"; -- multiplication by the radix
   sel8_c1 <= betaw8_c1(26 downto 21) & D_c1(22 downto 20);
   SelFunctionTable8: selFunction_Freq100_uid4
      port map ( X => sel8_c1,
                 Y => q8_copy11_c1);
   q8_c1 <= q8_copy11_c1; -- output copy to hold a pipeline register if needed

   with q8_c1  select 
      absq8D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q8_c1(2)  select 
   w7_c1<= betaw8_c1 - absq8D_c1 when '0',
         betaw8_c1 + absq8D_c1 when others;

   betaw7_c1 <= w7_c1(24 downto 0) & "00"; -- multiplication by the radix
   sel7_c1 <= betaw7_c1(26 downto 21) & D_c1(22 downto 20);
   SelFunctionTable7: selFunction_Freq100_uid4
      port map ( X => sel7_c1,
                 Y => q7_copy12_c1);
   q7_c1 <= q7_copy12_c1; -- output copy to hold a pipeline register if needed

   with q7_c1  select 
      absq7D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q7_c1(2)  select 
   w6_c1<= betaw7_c1 - absq7D_c1 when '0',
         betaw7_c1 + absq7D_c1 when others;

   betaw6_c1 <= w6_c1(24 downto 0) & "00"; -- multiplication by the radix
   sel6_c1 <= betaw6_c1(26 downto 21) & D_c1(22 downto 20);
   SelFunctionTable6: selFunction_Freq100_uid4
      port map ( X => sel6_c1,
                 Y => q6_copy13_c1);
   q6_c1 <= q6_copy13_c1; -- output copy to hold a pipeline register if needed

   with q6_c1  select 
      absq6D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q6_c1(2)  select 
   w5_c1<= betaw6_c1 - absq6D_c1 when '0',
         betaw6_c1 + absq6D_c1 when others;

   betaw5_c1 <= w5_c1(24 downto 0) & "00"; -- multiplication by the radix
   sel5_c1 <= betaw5_c1(26 downto 21) & D_c1(22 downto 20);
   SelFunctionTable5: selFunction_Freq100_uid4
      port map ( X => sel5_c1,
                 Y => q5_copy14_c1);
   q5_c1 <= q5_copy14_c1; -- output copy to hold a pipeline register if needed

   with q5_c1  select 
      absq5D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q5_c1(2)  select 
   w4_c1<= betaw5_c1 - absq5D_c1 when '0',
         betaw5_c1 + absq5D_c1 when others;

   betaw4_c1 <= w4_c1(24 downto 0) & "00"; -- multiplication by the radix
   sel4_c1 <= betaw4_c1(26 downto 21) & D_c1(22 downto 20);
   SelFunctionTable4: selFunction_Freq100_uid4
      port map ( X => sel4_c1,
                 Y => q4_copy15_c1);
   q4_c1 <= q4_copy15_c1; -- output copy to hold a pipeline register if needed

   with q4_c1  select 
      absq4D_c1 <= 
         "000" & D_c1						 when "001" | "111", -- mult by 1
         "00" & D_c1 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q4_c2(2)  select 
   w3_c2<= betaw4_c2 - absq4D_c2 when '0',
         betaw4_c2 + absq4D_c2 when others;

   betaw3_c2 <= w3_c2(24 downto 0) & "00"; -- multiplication by the radix
   sel3_c2 <= betaw3_c2(26 downto 21) & D_c2(22 downto 20);
   SelFunctionTable3: selFunction_Freq100_uid4
      port map ( X => sel3_c2,
                 Y => q3_copy16_c2);
   q3_c2 <= q3_copy16_c2; -- output copy to hold a pipeline register if needed

   with q3_c2  select 
      absq3D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q3_c2(2)  select 
   w2_c2<= betaw3_c2 - absq3D_c2 when '0',
         betaw3_c2 + absq3D_c2 when others;

   betaw2_c2 <= w2_c2(24 downto 0) & "00"; -- multiplication by the radix
   sel2_c2 <= betaw2_c2(26 downto 21) & D_c2(22 downto 20);
   SelFunctionTable2: selFunction_Freq100_uid4
      port map ( X => sel2_c2,
                 Y => q2_copy17_c2);
   q2_c2 <= q2_copy17_c2; -- output copy to hold a pipeline register if needed

   with q2_c2  select 
      absq2D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q2_c2(2)  select 
   w1_c2<= betaw2_c2 - absq2D_c2 when '0',
         betaw2_c2 + absq2D_c2 when others;

   betaw1_c2 <= w1_c2(24 downto 0) & "00"; -- multiplication by the radix
   sel1_c2 <= betaw1_c2(26 downto 21) & D_c2(22 downto 20);
   SelFunctionTable1: selFunction_Freq100_uid4
      port map ( X => sel1_c2,
                 Y => q1_copy18_c2);
   q1_c2 <= q1_copy18_c2; -- output copy to hold a pipeline register if needed

   with q1_c2  select 
      absq1D_c2 <= 
         "000" & D_c2						 when "001" | "111", -- mult by 1
         "00" & D_c2 & "0"			   when "010" | "110", -- mult by 2
         (26 downto 0 => '0')	 when others;        -- mult by 0

   with q1_c2(2)  select 
   w0_c2<= betaw1_c2 - absq1D_c2 when '0',
         betaw1_c2 + absq1D_c2 when others;

   wfinal_c2 <= w0_c2(24 downto 0);
   qM0_c2 <= wfinal_c2(24); -- rounding bit is the sign of the remainder
   qP14_c0 <=      q14_c0(1 downto 0);
   qM14_c0 <=      q14_c0(2) & "0";
   qP13_c0 <=      q13_c0(1 downto 0);
   qM13_c0 <=      q13_c0(2) & "0";
   qP12_c0 <=      q12_c0(1 downto 0);
   qM12_c0 <=      q12_c0(2) & "0";
   qP11_c0 <=      q11_c0(1 downto 0);
   qM11_c0 <=      q11_c0(2) & "0";
   qP10_c0 <=      q10_c0(1 downto 0);
   qM10_c0 <=      q10_c0(2) & "0";
   qP9_c0 <=      q9_c0(1 downto 0);
   qM9_c0 <=      q9_c0(2) & "0";
   qP8_c1 <=      q8_c1(1 downto 0);
   qM8_c1 <=      q8_c1(2) & "0";
   qP7_c1 <=      q7_c1(1 downto 0);
   qM7_c1 <=      q7_c1(2) & "0";
   qP6_c1 <=      q6_c1(1 downto 0);
   qM6_c1 <=      q6_c1(2) & "0";
   qP5_c1 <=      q5_c1(1 downto 0);
   qM5_c1 <=      q5_c1(2) & "0";
   qP4_c1 <=      q4_c1(1 downto 0);
   qM4_c1 <=      q4_c1(2) & "0";
   qP3_c2 <=      q3_c2(1 downto 0);
   qM3_c2 <=      q3_c2(2) & "0";
   qP2_c2 <=      q2_c2(1 downto 0);
   qM2_c2 <=      q2_c2(2) & "0";
   qP1_c2 <=      q1_c2(1 downto 0);
   qM1_c2 <=      q1_c2(2) & "0";
   qP_c2 <= qP14_c2 & qP13_c2 & qP12_c2 & qP11_c2 & qP10_c2 & qP9_c2 & qP8_c2 & qP7_c2 & qP6_c2 & qP5_c2 & qP4_c2 & qP3_c2 & qP2_c2 & qP1_c2;
   qM_c2 <= qM14_c2(0) & qM13_c2 & qM12_c2 & qM11_c2 & qM10_c2 & qM9_c2 & qM8_c2 & qM7_c2 & qM6_c2 & qM5_c2 & qM4_c2 & qM3_c2 & qM2_c2 & qM1_c2 & qM0_c2;
   quotient_c2 <= qP_c2 - qM_c2;
   -- We need a mR in (0, -wf-2) format: 1+wF fraction bits, 1 round bit, and 1 guard bit for the normalisation,
   -- quotient is the truncation of the exact quotient to at least 2^(-wF-2) bits
   -- now discarding its possible known MSB zeroes, and dropping the possible extra LSB bit (due to radix 4) 
   mR_c2 <= quotient_c2(26 downto 1); 
   -- normalisation
   fRnorm_c2 <=    mR_c2(24 downto 1)  when mR_c2(25)= '1'
           else mR_c2(23 downto 0);  -- now fRnorm is a (-1, -wF-1) fraction
   round_c2 <= fRnorm_c2(0); 
   expR1_c2 <= expR0_c2 + ("000" & (6 downto 1 => '1') & mR_c2(25)); -- add back bias
   -- final rounding
   expfrac_c2 <= expR1_c2 & fRnorm_c2(23 downto 1) ;
   expfracR_c2 <= expfrac_c2 + ((32 downto 1 => '0') & round_c2);
   exnR_c2 <=      "00"  when expfracR_c2(32) = '1'   -- underflow
           else "10"  when  expfracR_c2(32 downto 31) =  "01" -- overflow
           else "01";      -- 00, normal case
   with exnR0_c2  select 
      exnRfinal_c2 <= 
         exnR_c2   when "01", -- normal
         exnR0_c2  when others;
   R <= exnRfinal_c2 & sR_c2 & expfracR_c2(30 downto 0);
end architecture;




